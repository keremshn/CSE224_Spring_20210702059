magic
tech sky130A
magscale 1 2
timestamp 1746359154
<< viali >>
rect 34989 69445 35023 69479
rect 7113 69377 7147 69411
rect 21925 69377 21959 69411
rect 7665 69309 7699 69343
rect 22385 69309 22419 69343
rect 35725 69309 35759 69343
rect 11989 68765 12023 68799
rect 12173 68765 12207 68799
rect 12541 68765 12575 68799
rect 12817 68765 12851 68799
rect 13001 68765 13035 68799
rect 13461 68765 13495 68799
rect 31309 68765 31343 68799
rect 31493 68765 31527 68799
rect 31125 68629 31159 68663
rect 23029 68289 23063 68323
rect 23581 68289 23615 68323
rect 13093 67881 13127 67915
rect 12817 67813 12851 67847
rect 38025 67813 38059 67847
rect 12173 67745 12207 67779
rect 13277 67745 13311 67779
rect 1409 67677 1443 67711
rect 12541 67677 12575 67711
rect 12633 67677 12667 67711
rect 13461 67677 13495 67711
rect 13553 67677 13587 67711
rect 35265 67677 35299 67711
rect 36093 67677 36127 67711
rect 36185 67677 36219 67711
rect 37105 67677 37139 67711
rect 37473 67677 37507 67711
rect 37841 67677 37875 67711
rect 2237 67609 2271 67643
rect 35357 67609 35391 67643
rect 37657 67541 37691 67575
rect 37749 67541 37783 67575
rect 39681 67269 39715 67303
rect 9965 67201 9999 67235
rect 10241 67201 10275 67235
rect 10793 67201 10827 67235
rect 18061 67201 18095 67235
rect 18613 67201 18647 67235
rect 18981 67201 19015 67235
rect 38025 67201 38059 67235
rect 38301 67201 38335 67235
rect 40509 67201 40543 67235
rect 10517 67065 10551 67099
rect 18153 67065 18187 67099
rect 8125 66725 8159 66759
rect 7481 66589 7515 66623
rect 8217 66589 8251 66623
rect 26157 66589 26191 66623
rect 26341 66589 26375 66623
rect 26433 66589 26467 66623
rect 26525 66589 26559 66623
rect 26617 66589 26651 66623
rect 29653 66589 29687 66623
rect 30113 66589 30147 66623
rect 30389 66589 30423 66623
rect 26801 66453 26835 66487
rect 29653 66453 29687 66487
rect 4169 66113 4203 66147
rect 4353 66113 4387 66147
rect 4537 66113 4571 66147
rect 4997 66113 5031 66147
rect 35449 66113 35483 66147
rect 35817 66113 35851 66147
rect 36461 66113 36495 66147
rect 36737 66113 36771 66147
rect 35541 65909 35575 65943
rect 1961 65637 1995 65671
rect 2789 65569 2823 65603
rect 2479 65501 2513 65535
rect 2881 65501 2915 65535
rect 11897 65501 11931 65535
rect 2237 65433 2271 65467
rect 12265 65433 12299 65467
rect 3249 65365 3283 65399
rect 20821 64617 20855 64651
rect 7665 64549 7699 64583
rect 8309 64481 8343 64515
rect 20177 64481 20211 64515
rect 7849 64413 7883 64447
rect 8217 64413 8251 64447
rect 20085 64413 20119 64447
rect 20361 64413 20395 64447
rect 20453 64413 20487 64447
rect 20729 64413 20763 64447
rect 21097 64413 21131 64447
rect 21741 64413 21775 64447
rect 33701 64413 33735 64447
rect 33977 64413 34011 64447
rect 33609 64345 33643 64379
rect 20637 64277 20671 64311
rect 37749 63937 37783 63971
rect 37933 63937 37967 63971
rect 38117 63937 38151 63971
rect 37289 63869 37323 63903
rect 26985 63529 27019 63563
rect 27353 63529 27387 63563
rect 27537 63325 27571 63359
rect 27905 63325 27939 63359
rect 26709 63257 26743 63291
rect 17877 63189 17911 63223
rect 27721 63189 27755 63223
rect 18245 62985 18279 63019
rect 8125 62849 8159 62883
rect 8309 62849 8343 62883
rect 18307 62849 18341 62883
rect 17785 62781 17819 62815
rect 8493 62645 8527 62679
rect 17877 62645 17911 62679
rect 18429 62645 18463 62679
rect 20177 62373 20211 62407
rect 13277 62305 13311 62339
rect 34713 62305 34747 62339
rect 7389 62237 7423 62271
rect 7573 62237 7607 62271
rect 12173 62237 12207 62271
rect 12541 62237 12575 62271
rect 12909 62237 12943 62271
rect 13369 62237 13403 62271
rect 20453 62237 20487 62271
rect 34897 62237 34931 62271
rect 35265 62237 35299 62271
rect 35633 62237 35667 62271
rect 20361 62169 20395 62203
rect 20913 62169 20947 62203
rect 7481 62101 7515 62135
rect 17877 62101 17911 62135
rect 13277 61761 13311 61795
rect 13185 61693 13219 61727
rect 13737 61693 13771 61727
rect 17877 61557 17911 61591
rect 1501 61217 1535 61251
rect 1593 61149 1627 61183
rect 2421 61149 2455 61183
rect 4261 61149 4295 61183
rect 8953 61149 8987 61183
rect 9229 61149 9263 61183
rect 2329 61081 2363 61115
rect 4077 61081 4111 61115
rect 4169 61081 4203 61115
rect 4445 61081 4479 61115
rect 9137 61081 9171 61115
rect 9689 61081 9723 61115
rect 3893 61013 3927 61047
rect 4813 61013 4847 61047
rect 8125 60673 8159 60707
rect 8493 60673 8527 60707
rect 29009 60673 29043 60707
rect 29561 60673 29595 60707
rect 38669 60673 38703 60707
rect 38761 60673 38795 60707
rect 38945 60673 38979 60707
rect 8217 60605 8251 60639
rect 8677 60605 8711 60639
rect 38301 60537 38335 60571
rect 8861 60469 8895 60503
rect 19349 60469 19383 60503
rect 29101 60469 29135 60503
rect 39129 60469 39163 60503
rect 19625 60265 19659 60299
rect 34713 60265 34747 60299
rect 29653 60129 29687 60163
rect 19257 60061 19291 60095
rect 21741 60061 21775 60095
rect 22109 60061 22143 60095
rect 22201 60061 22235 60095
rect 30205 60061 30239 60095
rect 32689 60061 32723 60095
rect 33149 60061 33183 60095
rect 33425 60061 33459 60095
rect 33793 60061 33827 60095
rect 34161 60061 34195 60095
rect 34989 60061 35023 60095
rect 21281 59993 21315 60027
rect 32597 59993 32631 60027
rect 34713 59993 34747 60027
rect 19625 59925 19659 59959
rect 19809 59925 19843 59959
rect 34897 59925 34931 59959
rect 40325 59585 40359 59619
rect 39681 59517 39715 59551
rect 19349 59381 19383 59415
rect 7205 59109 7239 59143
rect 4721 59041 4755 59075
rect 30941 59041 30975 59075
rect 38117 59041 38151 59075
rect 4353 58973 4387 59007
rect 6745 58973 6779 59007
rect 22937 58973 22971 59007
rect 23213 58973 23247 59007
rect 29929 58973 29963 59007
rect 30481 58973 30515 59007
rect 38209 58973 38243 59007
rect 38393 58973 38427 59007
rect 4169 58905 4203 58939
rect 23121 58905 23155 58939
rect 23673 58905 23707 58939
rect 30021 58837 30055 58871
rect 2605 58565 2639 58599
rect 1409 58497 1443 58531
rect 13921 58497 13955 58531
rect 14381 58497 14415 58531
rect 14749 58497 14783 58531
rect 38669 58497 38703 58531
rect 39221 58497 39255 58531
rect 14013 58429 14047 58463
rect 26893 58089 26927 58123
rect 27537 58089 27571 58123
rect 19901 57953 19935 57987
rect 20085 57885 20119 57919
rect 20637 57885 20671 57919
rect 21005 57885 21039 57919
rect 24685 57885 24719 57919
rect 27813 57885 27847 57919
rect 27169 57817 27203 57851
rect 24501 57749 24535 57783
rect 27546 57749 27580 57783
rect 17141 57409 17175 57443
rect 39037 57409 39071 57443
rect 39589 57409 39623 57443
rect 39865 57409 39899 57443
rect 40233 57409 40267 57443
rect 16681 57341 16715 57375
rect 17233 57341 17267 57375
rect 39129 57273 39163 57307
rect 10149 56865 10183 56899
rect 26433 56865 26467 56899
rect 10057 56797 10091 56831
rect 10793 56797 10827 56831
rect 10885 56797 10919 56831
rect 11529 56797 11563 56831
rect 26341 56797 26375 56831
rect 26801 56797 26835 56831
rect 15945 55845 15979 55879
rect 9597 55777 9631 55811
rect 9505 55709 9539 55743
rect 9964 55709 9998 55743
rect 15853 55709 15887 55743
rect 16375 55709 16409 55743
rect 10149 55641 10183 55675
rect 16313 55573 16347 55607
rect 16497 55573 16531 55607
rect 4905 55233 4939 55267
rect 5273 55233 5307 55267
rect 5825 55029 5859 55063
rect 15485 54689 15519 54723
rect 6837 54621 6871 54655
rect 15761 54621 15795 54655
rect 33885 54621 33919 54655
rect 5549 54553 5583 54587
rect 6561 54553 6595 54587
rect 6929 54553 6963 54587
rect 4261 54485 4295 54519
rect 6745 54485 6779 54519
rect 7113 54485 7147 54519
rect 33977 54485 34011 54519
rect 15577 54213 15611 54247
rect 15393 54145 15427 54179
rect 28273 54145 28307 54179
rect 28641 54145 28675 54179
rect 29009 54145 29043 54179
rect 28365 53941 28399 53975
rect 4077 53533 4111 53567
rect 4353 53533 4387 53567
rect 15117 53533 15151 53567
rect 15393 53533 15427 53567
rect 38301 53533 38335 53567
rect 4537 53465 4571 53499
rect 15485 53465 15519 53499
rect 15853 53465 15887 53499
rect 39221 53465 39255 53499
rect 15301 53397 15335 53431
rect 37013 53125 37047 53159
rect 15301 53057 15335 53091
rect 15577 53057 15611 53091
rect 36829 53057 36863 53091
rect 15945 52989 15979 53023
rect 15301 52921 15335 52955
rect 36737 52853 36771 52887
rect 39313 52649 39347 52683
rect 39129 52581 39163 52615
rect 7389 52513 7423 52547
rect 35265 52513 35299 52547
rect 5549 52445 5583 52479
rect 6469 52445 6503 52479
rect 35081 52445 35115 52479
rect 35541 52445 35575 52479
rect 35817 52445 35851 52479
rect 36553 52445 36587 52479
rect 38853 52445 38887 52479
rect 34713 52377 34747 52411
rect 34897 52309 34931 52343
rect 34989 52309 35023 52343
rect 35817 52105 35851 52139
rect 21373 52037 21407 52071
rect 4721 51969 4755 52003
rect 4905 51969 4939 52003
rect 5457 51969 5491 52003
rect 21160 51969 21194 52003
rect 21281 51969 21315 52003
rect 21557 51969 21591 52003
rect 5365 51901 5399 51935
rect 20637 51901 20671 51935
rect 36277 51901 36311 51935
rect 21005 51765 21039 51799
rect 31769 51357 31803 51391
rect 32689 51357 32723 51391
rect 30849 51289 30883 51323
rect 10149 51017 10183 51051
rect 12475 51017 12509 51051
rect 12265 50949 12299 50983
rect 22109 50949 22143 50983
rect 10701 50881 10735 50915
rect 10885 50881 10919 50915
rect 12967 50881 13001 50915
rect 21833 50881 21867 50915
rect 22017 50881 22051 50915
rect 22201 50881 22235 50915
rect 22293 50881 22327 50915
rect 13277 50813 13311 50847
rect 13369 50813 13403 50847
rect 12633 50745 12667 50779
rect 12449 50677 12483 50711
rect 12817 50677 12851 50711
rect 22477 50677 22511 50711
rect 2973 50405 3007 50439
rect 2237 50337 2271 50371
rect 3249 50337 3283 50371
rect 2513 50269 2547 50303
rect 12541 50201 12575 50235
rect 12633 50133 12667 50167
rect 2605 49861 2639 49895
rect 39681 49861 39715 49895
rect 1409 49793 1443 49827
rect 13921 49793 13955 49827
rect 14197 49793 14231 49827
rect 23673 49793 23707 49827
rect 23949 49793 23983 49827
rect 24317 49793 24351 49827
rect 24685 49793 24719 49827
rect 35817 49793 35851 49827
rect 36369 49793 36403 49827
rect 36645 49793 36679 49827
rect 40509 49793 40543 49827
rect 14289 49725 14323 49759
rect 25053 49725 25087 49759
rect 36001 49657 36035 49691
rect 24409 49181 24443 49215
rect 24777 49113 24811 49147
rect 24593 49045 24627 49079
rect 24685 49045 24719 49079
rect 24869 49045 24903 49079
rect 17325 48841 17359 48875
rect 37381 48841 37415 48875
rect 10241 48705 10275 48739
rect 10425 48705 10459 48739
rect 16773 48705 16807 48739
rect 17049 48705 17083 48739
rect 17141 48705 17175 48739
rect 22385 48705 22419 48739
rect 22569 48705 22603 48739
rect 37289 48705 37323 48739
rect 37841 48705 37875 48739
rect 10793 48637 10827 48671
rect 10701 48569 10735 48603
rect 22477 48569 22511 48603
rect 16865 48501 16899 48535
rect 31033 47617 31067 47651
rect 31769 47549 31803 47583
rect 32505 45985 32539 46019
rect 32137 45917 32171 45951
rect 32597 45917 32631 45951
rect 23213 45509 23247 45543
rect 6469 45441 6503 45475
rect 6745 45441 6779 45475
rect 7481 45441 7515 45475
rect 8217 45441 8251 45475
rect 6653 45237 6687 45271
rect 24501 45237 24535 45271
rect 19809 44897 19843 44931
rect 32413 44897 32447 44931
rect 6377 44829 6411 44863
rect 6745 44829 6779 44863
rect 19625 44829 19659 44863
rect 32505 44829 32539 44863
rect 32873 44829 32907 44863
rect 32781 44761 32815 44795
rect 19441 44693 19475 44727
rect 10425 44421 10459 44455
rect 4721 44353 4755 44387
rect 4997 44353 5031 44387
rect 5181 44353 5215 44387
rect 18889 44353 18923 44387
rect 18981 44353 19015 44387
rect 19257 44353 19291 44387
rect 37473 44353 37507 44387
rect 38117 44353 38151 44387
rect 10241 44217 10275 44251
rect 5089 44149 5123 44183
rect 37565 44149 37599 44183
rect 9597 43265 9631 43299
rect 9689 43265 9723 43299
rect 11621 43265 11655 43299
rect 11713 43265 11747 43299
rect 12081 43265 12115 43299
rect 9781 43197 9815 43231
rect 9873 43197 9907 43231
rect 12265 43129 12299 43163
rect 9413 43061 9447 43095
rect 21557 42789 21591 42823
rect 20361 42653 20395 42687
rect 20637 42653 20671 42687
rect 20729 42653 20763 42687
rect 22477 42653 22511 42687
rect 23029 42653 23063 42687
rect 21097 42585 21131 42619
rect 22845 42585 22879 42619
rect 22661 42517 22695 42551
rect 22753 42517 22787 42551
rect 23581 42177 23615 42211
rect 23673 42177 23707 42211
rect 23949 42177 23983 42211
rect 24133 42177 24167 42211
rect 26985 42177 27019 42211
rect 32137 42177 32171 42211
rect 33701 42177 33735 42211
rect 27445 42109 27479 42143
rect 32873 42109 32907 42143
rect 33977 42109 34011 42143
rect 23029 41973 23063 42007
rect 33241 41633 33275 41667
rect 32689 41565 32723 41599
rect 33057 41565 33091 41599
rect 33793 41565 33827 41599
rect 2789 41089 2823 41123
rect 8033 41089 8067 41123
rect 8401 41089 8435 41123
rect 25881 41089 25915 41123
rect 28549 41089 28583 41123
rect 29285 41089 29319 41123
rect 29561 41089 29595 41123
rect 29929 41089 29963 41123
rect 30573 41089 30607 41123
rect 30941 41089 30975 41123
rect 3433 41021 3467 41055
rect 8493 41021 8527 41055
rect 30113 41021 30147 41055
rect 31033 41021 31067 41055
rect 7849 40953 7883 40987
rect 28641 40953 28675 40987
rect 25697 40885 25731 40919
rect 17141 40681 17175 40715
rect 22477 40681 22511 40715
rect 17233 40545 17267 40579
rect 31585 40545 31619 40579
rect 39221 40545 39255 40579
rect 2237 40477 2271 40511
rect 2881 40477 2915 40511
rect 3525 40477 3559 40511
rect 16957 40477 16991 40511
rect 22293 40477 22327 40511
rect 23121 40477 23155 40511
rect 23581 40477 23615 40511
rect 25145 40477 25179 40511
rect 32045 40477 32079 40511
rect 32137 40477 32171 40511
rect 3065 40409 3099 40443
rect 24593 40409 24627 40443
rect 16773 40341 16807 40375
rect 38669 40341 38703 40375
rect 1409 40069 1443 40103
rect 39313 40069 39347 40103
rect 40509 40001 40543 40035
rect 2237 39933 2271 39967
rect 12817 39593 12851 39627
rect 30481 39593 30515 39627
rect 28641 39525 28675 39559
rect 31309 39457 31343 39491
rect 13001 39389 13035 39423
rect 13093 39389 13127 39423
rect 13277 39389 13311 39423
rect 13369 39389 13403 39423
rect 23213 39389 23247 39423
rect 23305 39389 23339 39423
rect 23489 39389 23523 39423
rect 23673 39389 23707 39423
rect 25605 39389 25639 39423
rect 25973 39389 26007 39423
rect 26157 39389 26191 39423
rect 30021 39389 30055 39423
rect 30757 39389 30791 39423
rect 33149 39389 33183 39423
rect 23397 39321 23431 39355
rect 28825 39321 28859 39355
rect 23029 39253 23063 39287
rect 25697 39253 25731 39287
rect 32689 39253 32723 39287
rect 32337 39049 32371 39083
rect 32505 39049 32539 39083
rect 30389 38981 30423 39015
rect 32137 38981 32171 39015
rect 32781 38981 32815 39015
rect 20453 38913 20487 38947
rect 21281 38913 21315 38947
rect 29193 38913 29227 38947
rect 29285 38913 29319 38947
rect 29653 38913 29687 38947
rect 30757 38913 30791 38947
rect 30941 38913 30975 38947
rect 21557 38845 21591 38879
rect 23857 38845 23891 38879
rect 29561 38845 29595 38879
rect 20269 38777 20303 38811
rect 23397 38709 23431 38743
rect 30205 38709 30239 38743
rect 32321 38709 32355 38743
rect 19533 38505 19567 38539
rect 25145 38505 25179 38539
rect 24777 38369 24811 38403
rect 19809 38301 19843 38335
rect 24409 38301 24443 38335
rect 24593 38301 24627 38335
rect 24685 38301 24719 38335
rect 24961 38301 24995 38335
rect 19349 38165 19383 38199
rect 37381 37961 37415 37995
rect 37565 37961 37599 37995
rect 14565 37893 14599 37927
rect 25237 37893 25271 37927
rect 37657 37893 37691 37927
rect 12817 37825 12851 37859
rect 25697 37825 25731 37859
rect 25789 37825 25823 37859
rect 27077 37825 27111 37859
rect 27353 37825 27387 37859
rect 37749 37825 37783 37859
rect 27077 37689 27111 37723
rect 37933 37689 37967 37723
rect 25973 37621 26007 37655
rect 18429 37417 18463 37451
rect 39405 37349 39439 37383
rect 18521 37213 18555 37247
rect 35173 37213 35207 37247
rect 38853 37213 38887 37247
rect 39037 37213 39071 37247
rect 39221 37213 39255 37247
rect 17601 37077 17635 37111
rect 18061 37077 18095 37111
rect 35633 37077 35667 37111
rect 24961 36805 24995 36839
rect 38209 36805 38243 36839
rect 23949 36737 23983 36771
rect 24409 36737 24443 36771
rect 37933 36737 37967 36771
rect 38025 36737 38059 36771
rect 9873 36329 9907 36363
rect 35449 36261 35483 36295
rect 9689 36125 9723 36159
rect 9873 36125 9907 36159
rect 34897 36125 34931 36159
rect 35081 36125 35115 36159
rect 35265 36125 35299 36159
rect 3893 35785 3927 35819
rect 29837 35717 29871 35751
rect 4077 35649 4111 35683
rect 4169 35649 4203 35683
rect 4445 35649 4479 35683
rect 30205 35649 30239 35683
rect 30297 35649 30331 35683
rect 30113 35581 30147 35615
rect 29377 35513 29411 35547
rect 4353 35445 4387 35479
rect 3893 35241 3927 35275
rect 4077 35241 4111 35275
rect 10425 35241 10459 35275
rect 3525 35173 3559 35207
rect 12449 35105 12483 35139
rect 16681 35105 16715 35139
rect 27169 35105 27203 35139
rect 3249 35037 3283 35071
rect 3341 35037 3375 35071
rect 3525 35037 3559 35071
rect 9781 35037 9815 35071
rect 9873 35037 9907 35071
rect 10057 35037 10091 35071
rect 10241 35037 10275 35071
rect 12992 35037 13026 35071
rect 13185 35037 13219 35071
rect 13553 35037 13587 35071
rect 13737 35037 13771 35071
rect 13829 35037 13863 35071
rect 16497 35037 16531 35071
rect 17049 35037 17083 35071
rect 26617 35037 26651 35071
rect 26985 35037 27019 35071
rect 4261 34969 4295 35003
rect 10149 34969 10183 35003
rect 26709 34969 26743 35003
rect 4077 34901 4111 34935
rect 7573 34697 7607 34731
rect 38117 34697 38151 34731
rect 7205 34629 7239 34663
rect 7297 34629 7331 34663
rect 7021 34561 7055 34595
rect 7389 34561 7423 34595
rect 15577 34561 15611 34595
rect 15761 34561 15795 34595
rect 15945 34561 15979 34595
rect 21833 34561 21867 34595
rect 38301 34561 38335 34595
rect 38393 34561 38427 34595
rect 38669 34561 38703 34595
rect 23029 34493 23063 34527
rect 38577 34493 38611 34527
rect 2421 34085 2455 34119
rect 2237 33949 2271 33983
rect 2513 33949 2547 33983
rect 17049 33949 17083 33983
rect 32597 33949 32631 33983
rect 33333 33881 33367 33915
rect 2053 33813 2087 33847
rect 17233 33813 17267 33847
rect 18429 33609 18463 33643
rect 18597 33609 18631 33643
rect 6377 33541 6411 33575
rect 17785 33541 17819 33575
rect 18797 33541 18831 33575
rect 24869 33541 24903 33575
rect 6561 33473 6595 33507
rect 13737 33473 13771 33507
rect 14197 33473 14231 33507
rect 14657 33473 14691 33507
rect 15117 33473 15151 33507
rect 17693 33473 17727 33507
rect 17877 33473 17911 33507
rect 23213 33473 23247 33507
rect 23489 33473 23523 33507
rect 25421 33473 25455 33507
rect 26157 33473 26191 33507
rect 14289 33405 14323 33439
rect 6653 33269 6687 33303
rect 18613 33269 18647 33303
rect 16589 32997 16623 33031
rect 37289 32997 37323 33031
rect 39221 32997 39255 33031
rect 38669 32929 38703 32963
rect 33241 32861 33275 32895
rect 33517 32861 33551 32895
rect 37473 32861 37507 32895
rect 38117 32861 38151 32895
rect 38761 32861 38795 32895
rect 16773 32793 16807 32827
rect 6929 32521 6963 32555
rect 17049 32453 17083 32487
rect 29285 32453 29319 32487
rect 6377 32385 6411 32419
rect 6653 32385 6687 32419
rect 6745 32385 6779 32419
rect 16865 32385 16899 32419
rect 19901 32385 19935 32419
rect 19993 32385 20027 32419
rect 28641 32385 28675 32419
rect 28825 32385 28859 32419
rect 28917 32385 28951 32419
rect 29010 32385 29044 32419
rect 6469 32317 6503 32351
rect 20177 32317 20211 32351
rect 17233 32249 17267 32283
rect 16957 31909 16991 31943
rect 18521 31909 18555 31943
rect 18613 31909 18647 31943
rect 9689 31841 9723 31875
rect 1409 31773 1443 31807
rect 1685 31773 1719 31807
rect 9045 31773 9079 31807
rect 17417 31773 17451 31807
rect 30941 31773 30975 31807
rect 31125 31773 31159 31807
rect 31309 31773 31343 31807
rect 18981 31705 19015 31739
rect 16849 31365 16883 31399
rect 17049 31365 17083 31399
rect 40509 31297 40543 31331
rect 39681 31229 39715 31263
rect 16681 31093 16715 31127
rect 16865 31093 16899 31127
rect 36829 30821 36863 30855
rect 2053 30685 2087 30719
rect 2145 30685 2179 30719
rect 2329 30685 2363 30719
rect 2421 30685 2455 30719
rect 36399 30685 36433 30719
rect 36921 30685 36955 30719
rect 1869 30549 1903 30583
rect 36277 30549 36311 30583
rect 36461 30549 36495 30583
rect 31217 30209 31251 30243
rect 30389 30141 30423 30175
rect 30481 30141 30515 30175
rect 31309 30141 31343 30175
rect 35633 29801 35667 29835
rect 36461 29801 36495 29835
rect 20913 29665 20947 29699
rect 32597 29665 32631 29699
rect 21649 29597 21683 29631
rect 21741 29597 21775 29631
rect 22017 29597 22051 29631
rect 22109 29597 22143 29631
rect 31309 29597 31343 29631
rect 36001 29597 36035 29631
rect 36093 29597 36127 29631
rect 36277 29597 36311 29631
rect 36829 29597 36863 29631
rect 21925 29529 21959 29563
rect 31861 29529 31895 29563
rect 20453 29461 20487 29495
rect 22293 29461 22327 29495
rect 32137 29461 32171 29495
rect 38945 29257 38979 29291
rect 9045 29121 9079 29155
rect 9413 29121 9447 29155
rect 9689 29121 9723 29155
rect 11989 29121 12023 29155
rect 12357 29121 12391 29155
rect 38485 29121 38519 29155
rect 38761 29121 38795 29155
rect 10701 29053 10735 29087
rect 11345 29053 11379 29087
rect 12449 29053 12483 29087
rect 38577 29053 38611 29087
rect 11805 28985 11839 29019
rect 9137 28917 9171 28951
rect 10885 28713 10919 28747
rect 17417 28577 17451 28611
rect 17785 28577 17819 28611
rect 24501 28577 24535 28611
rect 10793 28509 10827 28543
rect 10977 28509 11011 28543
rect 16313 28509 16347 28543
rect 16405 28509 16439 28543
rect 16589 28509 16623 28543
rect 17325 28509 17359 28543
rect 24777 28509 24811 28543
rect 17141 28441 17175 28475
rect 16773 28373 16807 28407
rect 24869 28169 24903 28203
rect 24409 28033 24443 28067
rect 24685 28033 24719 28067
rect 31033 28033 31067 28067
rect 31401 28033 31435 28067
rect 31769 27965 31803 27999
rect 24501 27897 24535 27931
rect 31033 27897 31067 27931
rect 34805 27625 34839 27659
rect 34713 27421 34747 27455
rect 35081 27421 35115 27455
rect 35449 27421 35483 27455
rect 17969 26945 18003 26979
rect 18429 26945 18463 26979
rect 18521 26945 18555 26979
rect 18705 26877 18739 26911
rect 32597 26537 32631 26571
rect 31217 26469 31251 26503
rect 32137 26401 32171 26435
rect 32229 26401 32263 26435
rect 4077 26333 4111 26367
rect 4261 26333 4295 26367
rect 4629 26333 4663 26367
rect 31585 26333 31619 26367
rect 31770 26333 31804 26367
rect 30849 26197 30883 26231
rect 17601 25993 17635 26027
rect 18061 25925 18095 25959
rect 25237 25925 25271 25959
rect 6653 25857 6687 25891
rect 7389 25857 7423 25891
rect 7665 25857 7699 25891
rect 8125 25857 8159 25891
rect 24685 25857 24719 25891
rect 24869 25857 24903 25891
rect 6929 25789 6963 25823
rect 17693 25721 17727 25755
rect 10701 25381 10735 25415
rect 10517 25313 10551 25347
rect 38117 25313 38151 25347
rect 38577 25313 38611 25347
rect 10793 25245 10827 25279
rect 38393 25245 38427 25279
rect 37565 25177 37599 25211
rect 10333 25109 10367 25143
rect 7665 24769 7699 24803
rect 10517 24769 10551 24803
rect 10977 24769 11011 24803
rect 18337 24769 18371 24803
rect 19993 24769 20027 24803
rect 11253 24701 11287 24735
rect 10425 24633 10459 24667
rect 7205 24565 7239 24599
rect 33701 24361 33735 24395
rect 18981 24225 19015 24259
rect 7205 24157 7239 24191
rect 17785 24157 17819 24191
rect 18153 24157 18187 24191
rect 18705 24157 18739 24191
rect 33425 24157 33459 24191
rect 33517 24157 33551 24191
rect 8033 24089 8067 24123
rect 26065 24089 26099 24123
rect 26433 24089 26467 24123
rect 33701 24089 33735 24123
rect 26249 24021 26283 24055
rect 26341 24021 26375 24055
rect 26525 24021 26559 24055
rect 6929 23749 6963 23783
rect 34897 23749 34931 23783
rect 6653 23681 6687 23715
rect 6837 23681 6871 23715
rect 7073 23681 7107 23715
rect 7665 23681 7699 23715
rect 33885 23681 33919 23715
rect 34253 23681 34287 23715
rect 7757 23613 7791 23647
rect 33977 23613 34011 23647
rect 34161 23613 34195 23647
rect 7205 23545 7239 23579
rect 8217 23477 8251 23511
rect 6745 23205 6779 23239
rect 8401 23137 8435 23171
rect 6929 23069 6963 23103
rect 7297 23069 7331 23103
rect 7389 23069 7423 23103
rect 8309 23069 8343 23103
rect 20637 23069 20671 23103
rect 21189 23001 21223 23035
rect 7941 22933 7975 22967
rect 11713 22729 11747 22763
rect 11805 22729 11839 22763
rect 1685 22661 1719 22695
rect 11897 22661 11931 22695
rect 12265 22661 12299 22695
rect 14933 22661 14967 22695
rect 15025 22661 15059 22695
rect 1409 22593 1443 22627
rect 14657 22593 14691 22627
rect 17325 22593 17359 22627
rect 17601 22593 17635 22627
rect 18797 22593 18831 22627
rect 40509 22593 40543 22627
rect 11529 22525 11563 22559
rect 14519 22525 14553 22559
rect 19349 22525 19383 22559
rect 39681 22525 39715 22559
rect 16681 22457 16715 22491
rect 14381 22389 14415 22423
rect 15301 22049 15335 22083
rect 14841 21981 14875 22015
rect 15025 21981 15059 22015
rect 14565 21913 14599 21947
rect 7113 20961 7147 20995
rect 22109 20961 22143 20995
rect 22293 20961 22327 20995
rect 23029 20961 23063 20995
rect 3157 20893 3191 20927
rect 3249 20893 3283 20927
rect 3433 20893 3467 20927
rect 3525 20893 3559 20927
rect 7481 20893 7515 20927
rect 7849 20893 7883 20927
rect 22017 20893 22051 20927
rect 22385 20893 22419 20927
rect 8033 20825 8067 20859
rect 2973 20757 3007 20791
rect 1685 20553 1719 20587
rect 24869 20553 24903 20587
rect 1961 20485 1995 20519
rect 33149 20485 33183 20519
rect 1777 20417 1811 20451
rect 24133 20417 24167 20451
rect 24317 20417 24351 20451
rect 24777 20417 24811 20451
rect 25329 20417 25363 20451
rect 33333 20417 33367 20451
rect 33425 20417 33459 20451
rect 24685 20349 24719 20383
rect 25789 20349 25823 20383
rect 24593 20281 24627 20315
rect 33149 20213 33183 20247
rect 38117 19941 38151 19975
rect 4169 19873 4203 19907
rect 7573 19873 7607 19907
rect 37473 19873 37507 19907
rect 4077 19805 4111 19839
rect 4353 19805 4387 19839
rect 15761 19805 15795 19839
rect 33241 19805 33275 19839
rect 33793 19805 33827 19839
rect 37565 19805 37599 19839
rect 37933 19805 37967 19839
rect 16957 19737 16991 19771
rect 7113 19669 7147 19703
rect 13553 19397 13587 19431
rect 7113 19329 7147 19363
rect 7481 19329 7515 19363
rect 7849 19329 7883 19363
rect 12909 19329 12943 19363
rect 7757 19261 7791 19295
rect 17601 18853 17635 18887
rect 25789 18785 25823 18819
rect 26709 18785 26743 18819
rect 17877 18717 17911 18751
rect 18705 18717 18739 18751
rect 19257 18717 19291 18751
rect 26249 18717 26283 18751
rect 26433 18717 26467 18751
rect 26801 18717 26835 18751
rect 19441 18581 19475 18615
rect 29561 18377 29595 18411
rect 29469 18241 29503 18275
rect 30021 18241 30055 18275
rect 30297 18173 30331 18207
rect 38669 17833 38703 17867
rect 39129 17697 39163 17731
rect 38853 17629 38887 17663
rect 38945 17629 38979 17663
rect 39037 17629 39071 17663
rect 6561 16609 6595 16643
rect 7113 16609 7147 16643
rect 24501 16609 24535 16643
rect 25053 16609 25087 16643
rect 7021 16541 7055 16575
rect 24961 16541 24995 16575
rect 2421 16201 2455 16235
rect 1961 16065 1995 16099
rect 2480 16065 2514 16099
rect 2053 15997 2087 16031
rect 2605 15861 2639 15895
rect 13001 15657 13035 15691
rect 13461 15657 13495 15691
rect 13185 15453 13219 15487
rect 34713 15453 34747 15487
rect 13277 15385 13311 15419
rect 35541 15385 35575 15419
rect 14565 15045 14599 15079
rect 31033 15045 31067 15079
rect 37841 15045 37875 15079
rect 38393 15045 38427 15079
rect 15301 14977 15335 15011
rect 15577 14977 15611 15011
rect 31401 14977 31435 15011
rect 33701 14977 33735 15011
rect 34253 14977 34287 15011
rect 34529 14977 34563 15011
rect 35357 14977 35391 15011
rect 38301 14977 38335 15011
rect 15117 14909 15151 14943
rect 15485 14909 15519 14943
rect 34345 14909 34379 14943
rect 34989 14909 35023 14943
rect 35265 14909 35299 14943
rect 31769 14841 31803 14875
rect 38577 14773 38611 14807
rect 38669 14569 38703 14603
rect 31493 14501 31527 14535
rect 31953 14501 31987 14535
rect 39405 14433 39439 14467
rect 39497 14433 39531 14467
rect 31125 14365 31159 14399
rect 31309 14365 31343 14399
rect 31677 14365 31711 14399
rect 32229 14365 32263 14399
rect 32689 14365 32723 14399
rect 39221 14365 39255 14399
rect 39313 14365 39347 14399
rect 31033 14297 31067 14331
rect 39037 14229 39071 14263
rect 39037 14025 39071 14059
rect 1409 13889 1443 13923
rect 38025 13889 38059 13923
rect 38393 13889 38427 13923
rect 38761 13889 38795 13923
rect 40325 13889 40359 13923
rect 3157 13821 3191 13855
rect 39681 13821 39715 13855
rect 39589 13481 39623 13515
rect 39037 13277 39071 13311
rect 39410 13277 39444 13311
rect 39221 13209 39255 13243
rect 39313 13209 39347 13243
rect 23305 12937 23339 12971
rect 39037 12937 39071 12971
rect 23213 12801 23247 12835
rect 23397 12801 23431 12835
rect 16497 12189 16531 12223
rect 16681 12189 16715 12223
rect 16865 12189 16899 12223
rect 17325 12121 17359 12155
rect 2421 11101 2455 11135
rect 14933 11101 14967 11135
rect 15117 11101 15151 11135
rect 15301 11101 15335 11135
rect 32413 11101 32447 11135
rect 32597 11101 32631 11135
rect 33609 11101 33643 11135
rect 37473 11101 37507 11135
rect 3433 11033 3467 11067
rect 15761 11033 15795 11067
rect 36461 11033 36495 11067
rect 2697 10625 2731 10659
rect 3065 10625 3099 10659
rect 3157 10557 3191 10591
rect 2513 10489 2547 10523
rect 14197 9605 14231 9639
rect 16681 9605 16715 9639
rect 16865 9605 16899 9639
rect 13645 9537 13679 9571
rect 13829 9537 13863 9571
rect 14013 9537 14047 9571
rect 14289 9537 14323 9571
rect 17141 9537 17175 9571
rect 16865 9333 16899 9367
rect 35173 9129 35207 9163
rect 34805 9061 34839 9095
rect 1869 8993 1903 9027
rect 2329 8993 2363 9027
rect 34713 8993 34747 9027
rect 2237 8925 2271 8959
rect 2605 8925 2639 8959
rect 2789 8925 2823 8959
rect 27077 8925 27111 8959
rect 27537 8925 27571 8959
rect 34989 8925 35023 8959
rect 27169 8041 27203 8075
rect 37749 7973 37783 8007
rect 37473 7905 37507 7939
rect 15669 7837 15703 7871
rect 15853 7837 15887 7871
rect 16037 7837 16071 7871
rect 27721 7837 27755 7871
rect 28089 7837 28123 7871
rect 16497 7769 16531 7803
rect 37933 7701 37967 7735
rect 19809 7361 19843 7395
rect 20269 7361 20303 7395
rect 20729 7361 20763 7395
rect 21005 7361 21039 7395
rect 19901 7293 19935 7327
rect 34897 6749 34931 6783
rect 35541 6749 35575 6783
rect 35633 6749 35667 6783
rect 34713 6681 34747 6715
rect 5733 6409 5767 6443
rect 17417 6341 17451 6375
rect 5917 6273 5951 6307
rect 6193 6273 6227 6307
rect 16681 6273 16715 6307
rect 16773 6273 16807 6307
rect 16957 6273 16991 6307
rect 31217 6273 31251 6307
rect 31585 6273 31619 6307
rect 31861 6273 31895 6307
rect 5181 6205 5215 6239
rect 6101 6137 6135 6171
rect 8401 5253 8435 5287
rect 8217 5185 8251 5219
rect 8493 5185 8527 5219
rect 8590 5185 8624 5219
rect 8769 5049 8803 5083
rect 7205 4777 7239 4811
rect 38577 4709 38611 4743
rect 2237 4641 2271 4675
rect 3801 4641 3835 4675
rect 6745 4641 6779 4675
rect 14105 4641 14139 4675
rect 19993 4641 20027 4675
rect 37381 4641 37415 4675
rect 1409 4573 1443 4607
rect 4353 4573 4387 4607
rect 6653 4573 6687 4607
rect 6929 4573 6963 4607
rect 7021 4573 7055 4607
rect 14289 4573 14323 4607
rect 14933 4573 14967 4607
rect 15301 4573 15335 4607
rect 19441 4573 19475 4607
rect 19533 4573 19567 4607
rect 37473 4573 37507 4607
rect 37749 4573 37783 4607
rect 37933 4573 37967 4607
rect 38025 4573 38059 4607
rect 38393 4573 38427 4607
rect 4169 4505 4203 4539
rect 4261 4505 4295 4539
rect 4537 4505 4571 4539
rect 19257 4505 19291 4539
rect 19625 4505 19659 4539
rect 40509 4165 40543 4199
rect 6469 4097 6503 4131
rect 7573 4097 7607 4131
rect 34161 4097 34195 4131
rect 7481 4029 7515 4063
rect 39681 4029 39715 4063
rect 34161 3689 34195 3723
rect 10977 3621 11011 3655
rect 10333 3553 10367 3587
rect 7205 3485 7239 3519
rect 8217 3485 8251 3519
rect 10425 3485 10459 3519
rect 11161 3485 11195 3519
rect 12817 3485 12851 3519
rect 13369 3485 13403 3519
rect 13645 3485 13679 3519
rect 13921 3485 13955 3519
rect 8217 3349 8251 3383
rect 34161 3145 34195 3179
rect 28549 3077 28583 3111
rect 29653 3077 29687 3111
rect 28181 3009 28215 3043
rect 28641 3009 28675 3043
rect 28733 3009 28767 3043
rect 28917 3009 28951 3043
rect 29929 2873 29963 2907
rect 30113 2805 30147 2839
rect 39037 2533 39071 2567
rect 2513 2465 2547 2499
rect 2973 2397 3007 2431
rect 8125 2397 8159 2431
rect 13461 2397 13495 2431
rect 18153 2397 18187 2431
rect 18705 2397 18739 2431
rect 23673 2397 23707 2431
rect 29009 2397 29043 2431
rect 34161 2397 34195 2431
rect 39405 2397 39439 2431
rect 7757 2329 7791 2363
rect 23305 2329 23339 2363
rect 28641 2329 28675 2363
rect 13277 2261 13311 2295
rect 18521 2261 18555 2295
rect 23857 2261 23891 2295
rect 29193 2261 29227 2295
rect 34345 2261 34379 2295
rect 39589 2261 39623 2295
<< metal1 >>
rect 1104 69658 40848 69680
rect 1104 69606 2610 69658
rect 2662 69606 2674 69658
rect 2726 69606 2738 69658
rect 2790 69606 2802 69658
rect 2854 69606 2866 69658
rect 2918 69606 7610 69658
rect 7662 69606 7674 69658
rect 7726 69606 7738 69658
rect 7790 69606 7802 69658
rect 7854 69606 7866 69658
rect 7918 69606 12610 69658
rect 12662 69606 12674 69658
rect 12726 69606 12738 69658
rect 12790 69606 12802 69658
rect 12854 69606 12866 69658
rect 12918 69606 17610 69658
rect 17662 69606 17674 69658
rect 17726 69606 17738 69658
rect 17790 69606 17802 69658
rect 17854 69606 17866 69658
rect 17918 69606 22610 69658
rect 22662 69606 22674 69658
rect 22726 69606 22738 69658
rect 22790 69606 22802 69658
rect 22854 69606 22866 69658
rect 22918 69606 27610 69658
rect 27662 69606 27674 69658
rect 27726 69606 27738 69658
rect 27790 69606 27802 69658
rect 27854 69606 27866 69658
rect 27918 69606 32610 69658
rect 32662 69606 32674 69658
rect 32726 69606 32738 69658
rect 32790 69606 32802 69658
rect 32854 69606 32866 69658
rect 32918 69606 37610 69658
rect 37662 69606 37674 69658
rect 37726 69606 37738 69658
rect 37790 69606 37802 69658
rect 37854 69606 37866 69658
rect 37918 69606 40848 69658
rect 1104 69584 40848 69606
rect 34974 69436 34980 69488
rect 35032 69436 35038 69488
rect 7098 69368 7104 69420
rect 7156 69368 7162 69420
rect 20898 69368 20904 69420
rect 20956 69408 20962 69420
rect 21913 69411 21971 69417
rect 21913 69408 21925 69411
rect 20956 69380 21925 69408
rect 20956 69368 20962 69380
rect 21913 69377 21925 69380
rect 21959 69377 21971 69411
rect 21913 69371 21971 69377
rect 7653 69343 7711 69349
rect 7653 69309 7665 69343
rect 7699 69340 7711 69343
rect 9582 69340 9588 69352
rect 7699 69312 9588 69340
rect 7699 69309 7711 69312
rect 7653 69303 7711 69309
rect 9582 69300 9588 69312
rect 9640 69300 9646 69352
rect 22370 69300 22376 69352
rect 22428 69300 22434 69352
rect 35434 69300 35440 69352
rect 35492 69340 35498 69352
rect 35713 69343 35771 69349
rect 35713 69340 35725 69343
rect 35492 69312 35725 69340
rect 35492 69300 35498 69312
rect 35713 69309 35725 69312
rect 35759 69309 35771 69343
rect 35713 69303 35771 69309
rect 1104 69114 40848 69136
rect 1104 69062 1950 69114
rect 2002 69062 2014 69114
rect 2066 69062 2078 69114
rect 2130 69062 2142 69114
rect 2194 69062 2206 69114
rect 2258 69062 6950 69114
rect 7002 69062 7014 69114
rect 7066 69062 7078 69114
rect 7130 69062 7142 69114
rect 7194 69062 7206 69114
rect 7258 69062 11950 69114
rect 12002 69062 12014 69114
rect 12066 69062 12078 69114
rect 12130 69062 12142 69114
rect 12194 69062 12206 69114
rect 12258 69062 16950 69114
rect 17002 69062 17014 69114
rect 17066 69062 17078 69114
rect 17130 69062 17142 69114
rect 17194 69062 17206 69114
rect 17258 69062 21950 69114
rect 22002 69062 22014 69114
rect 22066 69062 22078 69114
rect 22130 69062 22142 69114
rect 22194 69062 22206 69114
rect 22258 69062 26950 69114
rect 27002 69062 27014 69114
rect 27066 69062 27078 69114
rect 27130 69062 27142 69114
rect 27194 69062 27206 69114
rect 27258 69062 31950 69114
rect 32002 69062 32014 69114
rect 32066 69062 32078 69114
rect 32130 69062 32142 69114
rect 32194 69062 32206 69114
rect 32258 69062 36950 69114
rect 37002 69062 37014 69114
rect 37066 69062 37078 69114
rect 37130 69062 37142 69114
rect 37194 69062 37206 69114
rect 37258 69062 40848 69114
rect 1104 69040 40848 69062
rect 11422 68756 11428 68808
rect 11480 68796 11486 68808
rect 11977 68799 12035 68805
rect 11977 68796 11989 68799
rect 11480 68768 11989 68796
rect 11480 68756 11486 68768
rect 11977 68765 11989 68768
rect 12023 68765 12035 68799
rect 11977 68759 12035 68765
rect 12161 68799 12219 68805
rect 12161 68765 12173 68799
rect 12207 68765 12219 68799
rect 12161 68759 12219 68765
rect 12529 68799 12587 68805
rect 12529 68765 12541 68799
rect 12575 68765 12587 68799
rect 12529 68759 12587 68765
rect 12805 68799 12863 68805
rect 12805 68765 12817 68799
rect 12851 68765 12863 68799
rect 12805 68759 12863 68765
rect 12989 68799 13047 68805
rect 12989 68765 13001 68799
rect 13035 68796 13047 68799
rect 13170 68796 13176 68808
rect 13035 68768 13176 68796
rect 13035 68765 13047 68768
rect 12989 68759 13047 68765
rect 11514 68688 11520 68740
rect 11572 68728 11578 68740
rect 12176 68728 12204 68759
rect 11572 68700 12204 68728
rect 11572 68688 11578 68700
rect 12544 68660 12572 68759
rect 12820 68728 12848 68759
rect 13170 68756 13176 68768
rect 13228 68756 13234 68808
rect 13449 68799 13507 68805
rect 13449 68765 13461 68799
rect 13495 68796 13507 68799
rect 15562 68796 15568 68808
rect 13495 68768 15568 68796
rect 13495 68765 13507 68768
rect 13449 68759 13507 68765
rect 15562 68756 15568 68768
rect 15620 68756 15626 68808
rect 28718 68756 28724 68808
rect 28776 68796 28782 68808
rect 31297 68799 31355 68805
rect 31297 68796 31309 68799
rect 28776 68768 31309 68796
rect 28776 68756 28782 68768
rect 31297 68765 31309 68768
rect 31343 68765 31355 68799
rect 31297 68759 31355 68765
rect 31478 68756 31484 68808
rect 31536 68756 31542 68808
rect 13262 68728 13268 68740
rect 12820 68700 13268 68728
rect 13262 68688 13268 68700
rect 13320 68688 13326 68740
rect 20162 68660 20168 68672
rect 12544 68632 20168 68660
rect 20162 68620 20168 68632
rect 20220 68620 20226 68672
rect 31110 68620 31116 68672
rect 31168 68620 31174 68672
rect 1104 68570 40848 68592
rect 1104 68518 2610 68570
rect 2662 68518 2674 68570
rect 2726 68518 2738 68570
rect 2790 68518 2802 68570
rect 2854 68518 2866 68570
rect 2918 68518 7610 68570
rect 7662 68518 7674 68570
rect 7726 68518 7738 68570
rect 7790 68518 7802 68570
rect 7854 68518 7866 68570
rect 7918 68518 12610 68570
rect 12662 68518 12674 68570
rect 12726 68518 12738 68570
rect 12790 68518 12802 68570
rect 12854 68518 12866 68570
rect 12918 68518 17610 68570
rect 17662 68518 17674 68570
rect 17726 68518 17738 68570
rect 17790 68518 17802 68570
rect 17854 68518 17866 68570
rect 17918 68518 22610 68570
rect 22662 68518 22674 68570
rect 22726 68518 22738 68570
rect 22790 68518 22802 68570
rect 22854 68518 22866 68570
rect 22918 68518 27610 68570
rect 27662 68518 27674 68570
rect 27726 68518 27738 68570
rect 27790 68518 27802 68570
rect 27854 68518 27866 68570
rect 27918 68518 32610 68570
rect 32662 68518 32674 68570
rect 32726 68518 32738 68570
rect 32790 68518 32802 68570
rect 32854 68518 32866 68570
rect 32918 68518 37610 68570
rect 37662 68518 37674 68570
rect 37726 68518 37738 68570
rect 37790 68518 37802 68570
rect 37854 68518 37866 68570
rect 37918 68518 40848 68570
rect 1104 68496 40848 68518
rect 23842 68348 23848 68400
rect 23900 68388 23906 68400
rect 23900 68360 23966 68388
rect 23900 68348 23906 68360
rect 19794 68280 19800 68332
rect 19852 68320 19858 68332
rect 23017 68323 23075 68329
rect 23017 68320 23029 68323
rect 19852 68292 23029 68320
rect 19852 68280 19858 68292
rect 23017 68289 23029 68292
rect 23063 68289 23075 68323
rect 23017 68283 23075 68289
rect 23106 68280 23112 68332
rect 23164 68320 23170 68332
rect 23569 68323 23627 68329
rect 23569 68320 23581 68323
rect 23164 68292 23581 68320
rect 23164 68280 23170 68292
rect 23569 68289 23581 68292
rect 23615 68289 23627 68323
rect 23569 68283 23627 68289
rect 1104 68026 40848 68048
rect 1104 67974 1950 68026
rect 2002 67974 2014 68026
rect 2066 67974 2078 68026
rect 2130 67974 2142 68026
rect 2194 67974 2206 68026
rect 2258 67974 6950 68026
rect 7002 67974 7014 68026
rect 7066 67974 7078 68026
rect 7130 67974 7142 68026
rect 7194 67974 7206 68026
rect 7258 67974 11950 68026
rect 12002 67974 12014 68026
rect 12066 67974 12078 68026
rect 12130 67974 12142 68026
rect 12194 67974 12206 68026
rect 12258 67974 16950 68026
rect 17002 67974 17014 68026
rect 17066 67974 17078 68026
rect 17130 67974 17142 68026
rect 17194 67974 17206 68026
rect 17258 67974 21950 68026
rect 22002 67974 22014 68026
rect 22066 67974 22078 68026
rect 22130 67974 22142 68026
rect 22194 67974 22206 68026
rect 22258 67974 26950 68026
rect 27002 67974 27014 68026
rect 27066 67974 27078 68026
rect 27130 67974 27142 68026
rect 27194 67974 27206 68026
rect 27258 67974 31950 68026
rect 32002 67974 32014 68026
rect 32066 67974 32078 68026
rect 32130 67974 32142 68026
rect 32194 67974 32206 68026
rect 32258 67974 36950 68026
rect 37002 67974 37014 68026
rect 37066 67974 37078 68026
rect 37130 67974 37142 68026
rect 37194 67974 37206 68026
rect 37258 67974 40848 68026
rect 1104 67952 40848 67974
rect 8938 67872 8944 67924
rect 8996 67912 9002 67924
rect 13081 67915 13139 67921
rect 13081 67912 13093 67915
rect 8996 67884 13093 67912
rect 8996 67872 9002 67884
rect 13081 67881 13093 67884
rect 13127 67881 13139 67915
rect 13081 67875 13139 67881
rect 35342 67872 35348 67924
rect 35400 67912 35406 67924
rect 35400 67884 38240 67912
rect 35400 67872 35406 67884
rect 12805 67847 12863 67853
rect 12805 67813 12817 67847
rect 12851 67844 12863 67847
rect 13630 67844 13636 67856
rect 12851 67816 13636 67844
rect 12851 67813 12863 67816
rect 12805 67807 12863 67813
rect 13630 67804 13636 67816
rect 13688 67804 13694 67856
rect 36188 67816 37964 67844
rect 12161 67779 12219 67785
rect 12161 67745 12173 67779
rect 12207 67776 12219 67779
rect 13265 67779 13323 67785
rect 12207 67748 12664 67776
rect 12207 67745 12219 67748
rect 12161 67739 12219 67745
rect 1394 67668 1400 67720
rect 1452 67668 1458 67720
rect 12636 67717 12664 67748
rect 13265 67745 13277 67779
rect 13311 67776 13323 67779
rect 26142 67776 26148 67788
rect 13311 67748 26148 67776
rect 13311 67745 13323 67748
rect 13265 67739 13323 67745
rect 26142 67736 26148 67748
rect 26200 67736 26206 67788
rect 12529 67711 12587 67717
rect 12529 67677 12541 67711
rect 12575 67677 12587 67711
rect 12529 67671 12587 67677
rect 12621 67711 12679 67717
rect 12621 67677 12633 67711
rect 12667 67708 12679 67711
rect 13078 67708 13084 67720
rect 12667 67680 13084 67708
rect 12667 67677 12679 67680
rect 12621 67671 12679 67677
rect 2225 67643 2283 67649
rect 2225 67609 2237 67643
rect 2271 67640 2283 67643
rect 6546 67640 6552 67652
rect 2271 67612 6552 67640
rect 2271 67609 2283 67612
rect 2225 67603 2283 67609
rect 6546 67600 6552 67612
rect 6604 67600 6610 67652
rect 12544 67640 12572 67671
rect 13078 67668 13084 67680
rect 13136 67668 13142 67720
rect 13446 67668 13452 67720
rect 13504 67668 13510 67720
rect 13538 67668 13544 67720
rect 13596 67668 13602 67720
rect 35250 67668 35256 67720
rect 35308 67668 35314 67720
rect 36188 67717 36216 67816
rect 37936 67776 37964 67816
rect 38010 67804 38016 67856
rect 38068 67804 38074 67856
rect 38102 67776 38108 67788
rect 37936 67748 38108 67776
rect 38102 67736 38108 67748
rect 38160 67736 38166 67788
rect 36081 67711 36139 67717
rect 36081 67677 36093 67711
rect 36127 67677 36139 67711
rect 36081 67671 36139 67677
rect 36173 67711 36231 67717
rect 36173 67677 36185 67711
rect 36219 67677 36231 67711
rect 36173 67671 36231 67677
rect 12986 67640 12992 67652
rect 12544 67612 12992 67640
rect 12986 67600 12992 67612
rect 13044 67600 13050 67652
rect 33134 67600 33140 67652
rect 33192 67640 33198 67652
rect 35345 67643 35403 67649
rect 35345 67640 35357 67643
rect 33192 67612 35357 67640
rect 33192 67600 33198 67612
rect 35345 67609 35357 67612
rect 35391 67609 35403 67643
rect 36096 67640 36124 67671
rect 37090 67668 37096 67720
rect 37148 67708 37154 67720
rect 37461 67711 37519 67717
rect 37461 67708 37473 67711
rect 37148 67680 37473 67708
rect 37148 67668 37154 67680
rect 37461 67677 37473 67680
rect 37507 67677 37519 67711
rect 37461 67671 37519 67677
rect 37829 67711 37887 67717
rect 37829 67677 37841 67711
rect 37875 67708 37887 67711
rect 38212 67708 38240 67884
rect 37875 67680 38240 67708
rect 37875 67677 37887 67680
rect 37829 67671 37887 67677
rect 36354 67640 36360 67652
rect 36096 67612 36360 67640
rect 35345 67603 35403 67609
rect 36354 67600 36360 67612
rect 36412 67600 36418 67652
rect 38378 67640 38384 67652
rect 37016 67612 37228 67640
rect 20530 67532 20536 67584
rect 20588 67572 20594 67584
rect 37016 67572 37044 67612
rect 20588 67544 37044 67572
rect 37200 67572 37228 67612
rect 37752 67612 38384 67640
rect 37752 67581 37780 67612
rect 38378 67600 38384 67612
rect 38436 67600 38442 67652
rect 37645 67575 37703 67581
rect 37645 67572 37657 67575
rect 37200 67544 37657 67572
rect 20588 67532 20594 67544
rect 37645 67541 37657 67544
rect 37691 67541 37703 67575
rect 37645 67535 37703 67541
rect 37737 67575 37795 67581
rect 37737 67541 37749 67575
rect 37783 67541 37795 67575
rect 37737 67535 37795 67541
rect 1104 67482 40848 67504
rect 1104 67430 2610 67482
rect 2662 67430 2674 67482
rect 2726 67430 2738 67482
rect 2790 67430 2802 67482
rect 2854 67430 2866 67482
rect 2918 67430 7610 67482
rect 7662 67430 7674 67482
rect 7726 67430 7738 67482
rect 7790 67430 7802 67482
rect 7854 67430 7866 67482
rect 7918 67430 12610 67482
rect 12662 67430 12674 67482
rect 12726 67430 12738 67482
rect 12790 67430 12802 67482
rect 12854 67430 12866 67482
rect 12918 67430 17610 67482
rect 17662 67430 17674 67482
rect 17726 67430 17738 67482
rect 17790 67430 17802 67482
rect 17854 67430 17866 67482
rect 17918 67430 22610 67482
rect 22662 67430 22674 67482
rect 22726 67430 22738 67482
rect 22790 67430 22802 67482
rect 22854 67430 22866 67482
rect 22918 67430 27610 67482
rect 27662 67430 27674 67482
rect 27726 67430 27738 67482
rect 27790 67430 27802 67482
rect 27854 67430 27866 67482
rect 27918 67430 32610 67482
rect 32662 67430 32674 67482
rect 32726 67430 32738 67482
rect 32790 67430 32802 67482
rect 32854 67430 32866 67482
rect 32918 67430 37610 67482
rect 37662 67430 37674 67482
rect 37726 67430 37738 67482
rect 37790 67430 37802 67482
rect 37854 67430 37866 67482
rect 37918 67430 40848 67482
rect 1104 67408 40848 67430
rect 18138 67300 18144 67312
rect 9968 67272 18144 67300
rect 9968 67241 9996 67272
rect 18138 67260 18144 67272
rect 18196 67260 18202 67312
rect 37274 67260 37280 67312
rect 37332 67300 37338 67312
rect 37332 67272 37674 67300
rect 37332 67260 37338 67272
rect 38838 67260 38844 67312
rect 38896 67300 38902 67312
rect 39669 67303 39727 67309
rect 39669 67300 39681 67303
rect 38896 67272 39681 67300
rect 38896 67260 38902 67272
rect 39669 67269 39681 67272
rect 39715 67269 39727 67303
rect 39669 67263 39727 67269
rect 9953 67235 10011 67241
rect 9953 67201 9965 67235
rect 9999 67201 10011 67235
rect 9953 67195 10011 67201
rect 10229 67235 10287 67241
rect 10229 67201 10241 67235
rect 10275 67232 10287 67235
rect 10781 67235 10839 67241
rect 10275 67204 10640 67232
rect 10275 67201 10287 67204
rect 10229 67195 10287 67201
rect 10502 67056 10508 67108
rect 10560 67056 10566 67108
rect 10612 67028 10640 67204
rect 10781 67201 10793 67235
rect 10827 67201 10839 67235
rect 10781 67195 10839 67201
rect 10796 67164 10824 67195
rect 13170 67192 13176 67244
rect 13228 67232 13234 67244
rect 18049 67235 18107 67241
rect 18049 67232 18061 67235
rect 13228 67204 18061 67232
rect 13228 67192 13234 67204
rect 18049 67201 18061 67204
rect 18095 67201 18107 67235
rect 18049 67195 18107 67201
rect 18598 67192 18604 67244
rect 18656 67192 18662 67244
rect 18969 67235 19027 67241
rect 18969 67201 18981 67235
rect 19015 67232 19027 67235
rect 23290 67232 23296 67244
rect 19015 67204 23296 67232
rect 19015 67201 19027 67204
rect 18969 67195 19027 67201
rect 23290 67192 23296 67204
rect 23348 67192 23354 67244
rect 24118 67192 24124 67244
rect 24176 67232 24182 67244
rect 24176 67204 26234 67232
rect 24176 67192 24182 67204
rect 18230 67164 18236 67176
rect 10796 67136 18236 67164
rect 18230 67124 18236 67136
rect 18288 67124 18294 67176
rect 18141 67099 18199 67105
rect 18141 67065 18153 67099
rect 18187 67096 18199 67099
rect 18322 67096 18328 67108
rect 18187 67068 18328 67096
rect 18187 67065 18199 67068
rect 18141 67059 18199 67065
rect 18322 67056 18328 67068
rect 18380 67056 18386 67108
rect 26206 67096 26234 67204
rect 38010 67192 38016 67244
rect 38068 67192 38074 67244
rect 38286 67192 38292 67244
rect 38344 67192 38350 67244
rect 40494 67192 40500 67244
rect 40552 67192 40558 67244
rect 38286 67096 38292 67108
rect 26206 67068 38292 67096
rect 38286 67056 38292 67068
rect 38344 67056 38350 67108
rect 20070 67028 20076 67040
rect 10612 67000 20076 67028
rect 20070 66988 20076 67000
rect 20128 66988 20134 67040
rect 1104 66938 40848 66960
rect 1104 66886 1950 66938
rect 2002 66886 2014 66938
rect 2066 66886 2078 66938
rect 2130 66886 2142 66938
rect 2194 66886 2206 66938
rect 2258 66886 6950 66938
rect 7002 66886 7014 66938
rect 7066 66886 7078 66938
rect 7130 66886 7142 66938
rect 7194 66886 7206 66938
rect 7258 66886 11950 66938
rect 12002 66886 12014 66938
rect 12066 66886 12078 66938
rect 12130 66886 12142 66938
rect 12194 66886 12206 66938
rect 12258 66886 16950 66938
rect 17002 66886 17014 66938
rect 17066 66886 17078 66938
rect 17130 66886 17142 66938
rect 17194 66886 17206 66938
rect 17258 66886 21950 66938
rect 22002 66886 22014 66938
rect 22066 66886 22078 66938
rect 22130 66886 22142 66938
rect 22194 66886 22206 66938
rect 22258 66886 26950 66938
rect 27002 66886 27014 66938
rect 27066 66886 27078 66938
rect 27130 66886 27142 66938
rect 27194 66886 27206 66938
rect 27258 66886 31950 66938
rect 32002 66886 32014 66938
rect 32066 66886 32078 66938
rect 32130 66886 32142 66938
rect 32194 66886 32206 66938
rect 32258 66886 36950 66938
rect 37002 66886 37014 66938
rect 37066 66886 37078 66938
rect 37130 66886 37142 66938
rect 37194 66886 37206 66938
rect 37258 66886 40848 66938
rect 1104 66864 40848 66886
rect 8110 66716 8116 66768
rect 8168 66716 8174 66768
rect 7466 66580 7472 66632
rect 7524 66580 7530 66632
rect 8205 66623 8263 66629
rect 8205 66589 8217 66623
rect 8251 66620 8263 66623
rect 10410 66620 10416 66632
rect 8251 66592 10416 66620
rect 8251 66589 8263 66592
rect 8205 66583 8263 66589
rect 10410 66580 10416 66592
rect 10468 66580 10474 66632
rect 26142 66580 26148 66632
rect 26200 66580 26206 66632
rect 26326 66580 26332 66632
rect 26384 66580 26390 66632
rect 26418 66580 26424 66632
rect 26476 66580 26482 66632
rect 26513 66623 26571 66629
rect 26513 66589 26525 66623
rect 26559 66589 26571 66623
rect 26513 66583 26571 66589
rect 26605 66623 26663 66629
rect 26605 66589 26617 66623
rect 26651 66589 26663 66623
rect 26605 66583 26663 66589
rect 18966 66512 18972 66564
rect 19024 66552 19030 66564
rect 26528 66552 26556 66583
rect 19024 66524 26556 66552
rect 26620 66552 26648 66583
rect 29638 66580 29644 66632
rect 29696 66580 29702 66632
rect 30098 66580 30104 66632
rect 30156 66580 30162 66632
rect 30282 66580 30288 66632
rect 30340 66620 30346 66632
rect 30377 66623 30435 66629
rect 30377 66620 30389 66623
rect 30340 66592 30389 66620
rect 30340 66580 30346 66592
rect 30377 66589 30389 66592
rect 30423 66589 30435 66623
rect 30377 66583 30435 66589
rect 34698 66552 34704 66564
rect 26620 66524 34704 66552
rect 19024 66512 19030 66524
rect 34698 66512 34704 66524
rect 34756 66512 34762 66564
rect 20622 66444 20628 66496
rect 20680 66484 20686 66496
rect 26789 66487 26847 66493
rect 26789 66484 26801 66487
rect 20680 66456 26801 66484
rect 20680 66444 20686 66456
rect 26789 66453 26801 66456
rect 26835 66453 26847 66487
rect 26789 66447 26847 66453
rect 29362 66444 29368 66496
rect 29420 66484 29426 66496
rect 29641 66487 29699 66493
rect 29641 66484 29653 66487
rect 29420 66456 29653 66484
rect 29420 66444 29426 66456
rect 29641 66453 29653 66456
rect 29687 66453 29699 66487
rect 29641 66447 29699 66453
rect 1104 66394 40848 66416
rect 1104 66342 2610 66394
rect 2662 66342 2674 66394
rect 2726 66342 2738 66394
rect 2790 66342 2802 66394
rect 2854 66342 2866 66394
rect 2918 66342 7610 66394
rect 7662 66342 7674 66394
rect 7726 66342 7738 66394
rect 7790 66342 7802 66394
rect 7854 66342 7866 66394
rect 7918 66342 12610 66394
rect 12662 66342 12674 66394
rect 12726 66342 12738 66394
rect 12790 66342 12802 66394
rect 12854 66342 12866 66394
rect 12918 66342 17610 66394
rect 17662 66342 17674 66394
rect 17726 66342 17738 66394
rect 17790 66342 17802 66394
rect 17854 66342 17866 66394
rect 17918 66342 22610 66394
rect 22662 66342 22674 66394
rect 22726 66342 22738 66394
rect 22790 66342 22802 66394
rect 22854 66342 22866 66394
rect 22918 66342 27610 66394
rect 27662 66342 27674 66394
rect 27726 66342 27738 66394
rect 27790 66342 27802 66394
rect 27854 66342 27866 66394
rect 27918 66342 32610 66394
rect 32662 66342 32674 66394
rect 32726 66342 32738 66394
rect 32790 66342 32802 66394
rect 32854 66342 32866 66394
rect 32918 66342 37610 66394
rect 37662 66342 37674 66394
rect 37726 66342 37738 66394
rect 37790 66342 37802 66394
rect 37854 66342 37866 66394
rect 37918 66342 40848 66394
rect 1104 66320 40848 66342
rect 39574 66212 39580 66224
rect 36464 66184 39580 66212
rect 4157 66147 4215 66153
rect 4157 66113 4169 66147
rect 4203 66113 4215 66147
rect 4157 66107 4215 66113
rect 4341 66147 4399 66153
rect 4341 66113 4353 66147
rect 4387 66113 4399 66147
rect 4341 66107 4399 66113
rect 4172 66008 4200 66107
rect 4356 66076 4384 66107
rect 4522 66104 4528 66156
rect 4580 66104 4586 66156
rect 4985 66147 5043 66153
rect 4985 66113 4997 66147
rect 5031 66144 5043 66147
rect 6454 66144 6460 66156
rect 5031 66116 6460 66144
rect 5031 66113 5043 66116
rect 4985 66107 5043 66113
rect 6454 66104 6460 66116
rect 6512 66104 6518 66156
rect 23382 66104 23388 66156
rect 23440 66144 23446 66156
rect 36464 66153 36492 66184
rect 39574 66172 39580 66184
rect 39632 66172 39638 66224
rect 35437 66147 35495 66153
rect 35437 66144 35449 66147
rect 23440 66116 35449 66144
rect 23440 66104 23446 66116
rect 35437 66113 35449 66116
rect 35483 66113 35495 66147
rect 35437 66107 35495 66113
rect 35805 66147 35863 66153
rect 35805 66113 35817 66147
rect 35851 66113 35863 66147
rect 35805 66107 35863 66113
rect 36449 66147 36507 66153
rect 36449 66113 36461 66147
rect 36495 66113 36507 66147
rect 36449 66107 36507 66113
rect 36725 66147 36783 66153
rect 36725 66113 36737 66147
rect 36771 66113 36783 66147
rect 36725 66107 36783 66113
rect 13170 66076 13176 66088
rect 4356 66048 13176 66076
rect 13170 66036 13176 66048
rect 13228 66036 13234 66088
rect 31018 66036 31024 66088
rect 31076 66076 31082 66088
rect 35820 66076 35848 66107
rect 31076 66048 35848 66076
rect 31076 66036 31082 66048
rect 35986 66036 35992 66088
rect 36044 66076 36050 66088
rect 36740 66076 36768 66107
rect 36044 66048 36768 66076
rect 36044 66036 36050 66048
rect 4982 66008 4988 66020
rect 4172 65980 4988 66008
rect 4982 65968 4988 65980
rect 5040 65968 5046 66020
rect 18874 65968 18880 66020
rect 18932 66008 18938 66020
rect 26418 66008 26424 66020
rect 18932 65980 26424 66008
rect 18932 65968 18938 65980
rect 26418 65968 26424 65980
rect 26476 65968 26482 66020
rect 24670 65900 24676 65952
rect 24728 65940 24734 65952
rect 35529 65943 35587 65949
rect 35529 65940 35541 65943
rect 24728 65912 35541 65940
rect 24728 65900 24734 65912
rect 35529 65909 35541 65912
rect 35575 65909 35587 65943
rect 35529 65903 35587 65909
rect 1104 65850 40848 65872
rect 1104 65798 1950 65850
rect 2002 65798 2014 65850
rect 2066 65798 2078 65850
rect 2130 65798 2142 65850
rect 2194 65798 2206 65850
rect 2258 65798 6950 65850
rect 7002 65798 7014 65850
rect 7066 65798 7078 65850
rect 7130 65798 7142 65850
rect 7194 65798 7206 65850
rect 7258 65798 11950 65850
rect 12002 65798 12014 65850
rect 12066 65798 12078 65850
rect 12130 65798 12142 65850
rect 12194 65798 12206 65850
rect 12258 65798 16950 65850
rect 17002 65798 17014 65850
rect 17066 65798 17078 65850
rect 17130 65798 17142 65850
rect 17194 65798 17206 65850
rect 17258 65798 21950 65850
rect 22002 65798 22014 65850
rect 22066 65798 22078 65850
rect 22130 65798 22142 65850
rect 22194 65798 22206 65850
rect 22258 65798 26950 65850
rect 27002 65798 27014 65850
rect 27066 65798 27078 65850
rect 27130 65798 27142 65850
rect 27194 65798 27206 65850
rect 27258 65798 31950 65850
rect 32002 65798 32014 65850
rect 32066 65798 32078 65850
rect 32130 65798 32142 65850
rect 32194 65798 32206 65850
rect 32258 65798 36950 65850
rect 37002 65798 37014 65850
rect 37066 65798 37078 65850
rect 37130 65798 37142 65850
rect 37194 65798 37206 65850
rect 37258 65798 40848 65850
rect 1104 65776 40848 65798
rect 14550 65696 14556 65748
rect 14608 65736 14614 65748
rect 26326 65736 26332 65748
rect 14608 65708 26332 65736
rect 14608 65696 14614 65708
rect 26326 65696 26332 65708
rect 26384 65696 26390 65748
rect 30558 65696 30564 65748
rect 30616 65736 30622 65748
rect 33134 65736 33140 65748
rect 30616 65708 33140 65736
rect 30616 65696 30622 65708
rect 33134 65696 33140 65708
rect 33192 65696 33198 65748
rect 1949 65671 2007 65677
rect 1949 65637 1961 65671
rect 1995 65668 2007 65671
rect 1995 65640 3096 65668
rect 1995 65637 2007 65640
rect 1949 65631 2007 65637
rect 2777 65603 2835 65609
rect 2777 65569 2789 65603
rect 2823 65600 2835 65603
rect 2958 65600 2964 65612
rect 2823 65572 2964 65600
rect 2823 65569 2835 65572
rect 2777 65563 2835 65569
rect 2958 65560 2964 65572
rect 3016 65560 3022 65612
rect 2467 65535 2525 65541
rect 2467 65501 2479 65535
rect 2513 65532 2525 65535
rect 2869 65535 2927 65541
rect 2513 65504 2820 65532
rect 2513 65501 2525 65504
rect 2467 65495 2525 65501
rect 1578 65424 1584 65476
rect 1636 65464 1642 65476
rect 2225 65467 2283 65473
rect 2225 65464 2237 65467
rect 1636 65436 2237 65464
rect 1636 65424 1642 65436
rect 2225 65433 2237 65436
rect 2271 65433 2283 65467
rect 2792 65464 2820 65504
rect 2869 65501 2881 65535
rect 2915 65532 2927 65535
rect 3068 65532 3096 65640
rect 13078 65628 13084 65680
rect 13136 65668 13142 65680
rect 25498 65668 25504 65680
rect 13136 65640 25504 65668
rect 13136 65628 13142 65640
rect 25498 65628 25504 65640
rect 25556 65628 25562 65680
rect 25590 65628 25596 65680
rect 25648 65668 25654 65680
rect 30098 65668 30104 65680
rect 25648 65640 30104 65668
rect 25648 65628 25654 65640
rect 30098 65628 30104 65640
rect 30156 65628 30162 65680
rect 6362 65560 6368 65612
rect 6420 65600 6426 65612
rect 20530 65600 20536 65612
rect 6420 65572 20536 65600
rect 6420 65560 6426 65572
rect 20530 65560 20536 65572
rect 20588 65560 20594 65612
rect 21726 65560 21732 65612
rect 21784 65600 21790 65612
rect 37274 65600 37280 65612
rect 21784 65572 37280 65600
rect 21784 65560 21790 65572
rect 37274 65560 37280 65572
rect 37332 65560 37338 65612
rect 2915 65504 6914 65532
rect 2915 65501 2927 65504
rect 2869 65495 2927 65501
rect 6886 65464 6914 65504
rect 9582 65492 9588 65544
rect 9640 65532 9646 65544
rect 11882 65532 11888 65544
rect 9640 65504 11888 65532
rect 9640 65492 9646 65504
rect 11882 65492 11888 65504
rect 11940 65492 11946 65544
rect 11992 65504 16574 65532
rect 11992 65464 12020 65504
rect 2792 65436 3280 65464
rect 6886 65436 12020 65464
rect 12253 65467 12311 65473
rect 2225 65427 2283 65433
rect 3252 65405 3280 65436
rect 12253 65433 12265 65467
rect 12299 65464 12311 65467
rect 12342 65464 12348 65476
rect 12299 65436 12348 65464
rect 12299 65433 12311 65436
rect 12253 65427 12311 65433
rect 12342 65424 12348 65436
rect 12400 65424 12406 65476
rect 16546 65464 16574 65504
rect 30466 65464 30472 65476
rect 16546 65436 30472 65464
rect 30466 65424 30472 65436
rect 30524 65424 30530 65476
rect 3237 65399 3295 65405
rect 3237 65365 3249 65399
rect 3283 65396 3295 65399
rect 19610 65396 19616 65408
rect 3283 65368 19616 65396
rect 3283 65365 3295 65368
rect 3237 65359 3295 65365
rect 19610 65356 19616 65368
rect 19668 65356 19674 65408
rect 1104 65306 40848 65328
rect 1104 65254 2610 65306
rect 2662 65254 2674 65306
rect 2726 65254 2738 65306
rect 2790 65254 2802 65306
rect 2854 65254 2866 65306
rect 2918 65254 7610 65306
rect 7662 65254 7674 65306
rect 7726 65254 7738 65306
rect 7790 65254 7802 65306
rect 7854 65254 7866 65306
rect 7918 65254 12610 65306
rect 12662 65254 12674 65306
rect 12726 65254 12738 65306
rect 12790 65254 12802 65306
rect 12854 65254 12866 65306
rect 12918 65254 17610 65306
rect 17662 65254 17674 65306
rect 17726 65254 17738 65306
rect 17790 65254 17802 65306
rect 17854 65254 17866 65306
rect 17918 65254 22610 65306
rect 22662 65254 22674 65306
rect 22726 65254 22738 65306
rect 22790 65254 22802 65306
rect 22854 65254 22866 65306
rect 22918 65254 27610 65306
rect 27662 65254 27674 65306
rect 27726 65254 27738 65306
rect 27790 65254 27802 65306
rect 27854 65254 27866 65306
rect 27918 65254 32610 65306
rect 32662 65254 32674 65306
rect 32726 65254 32738 65306
rect 32790 65254 32802 65306
rect 32854 65254 32866 65306
rect 32918 65254 37610 65306
rect 37662 65254 37674 65306
rect 37726 65254 37738 65306
rect 37790 65254 37802 65306
rect 37854 65254 37866 65306
rect 37918 65254 40848 65306
rect 1104 65232 40848 65254
rect 11882 65152 11888 65204
rect 11940 65192 11946 65204
rect 16390 65192 16396 65204
rect 11940 65164 16396 65192
rect 11940 65152 11946 65164
rect 16390 65152 16396 65164
rect 16448 65152 16454 65204
rect 7834 64812 7840 64864
rect 7892 64852 7898 64864
rect 31110 64852 31116 64864
rect 7892 64824 31116 64852
rect 7892 64812 7898 64824
rect 31110 64812 31116 64824
rect 31168 64812 31174 64864
rect 1104 64762 40848 64784
rect 1104 64710 1950 64762
rect 2002 64710 2014 64762
rect 2066 64710 2078 64762
rect 2130 64710 2142 64762
rect 2194 64710 2206 64762
rect 2258 64710 6950 64762
rect 7002 64710 7014 64762
rect 7066 64710 7078 64762
rect 7130 64710 7142 64762
rect 7194 64710 7206 64762
rect 7258 64710 11950 64762
rect 12002 64710 12014 64762
rect 12066 64710 12078 64762
rect 12130 64710 12142 64762
rect 12194 64710 12206 64762
rect 12258 64710 16950 64762
rect 17002 64710 17014 64762
rect 17066 64710 17078 64762
rect 17130 64710 17142 64762
rect 17194 64710 17206 64762
rect 17258 64710 21950 64762
rect 22002 64710 22014 64762
rect 22066 64710 22078 64762
rect 22130 64710 22142 64762
rect 22194 64710 22206 64762
rect 22258 64710 26950 64762
rect 27002 64710 27014 64762
rect 27066 64710 27078 64762
rect 27130 64710 27142 64762
rect 27194 64710 27206 64762
rect 27258 64710 31950 64762
rect 32002 64710 32014 64762
rect 32066 64710 32078 64762
rect 32130 64710 32142 64762
rect 32194 64710 32206 64762
rect 32258 64710 36950 64762
rect 37002 64710 37014 64762
rect 37066 64710 37078 64762
rect 37130 64710 37142 64762
rect 37194 64710 37206 64762
rect 37258 64710 40848 64762
rect 1104 64688 40848 64710
rect 13998 64608 14004 64660
rect 14056 64648 14062 64660
rect 20622 64648 20628 64660
rect 14056 64620 20628 64648
rect 14056 64608 14062 64620
rect 20622 64608 20628 64620
rect 20680 64608 20686 64660
rect 20806 64608 20812 64660
rect 20864 64608 20870 64660
rect 7653 64583 7711 64589
rect 7653 64549 7665 64583
rect 7699 64580 7711 64583
rect 8110 64580 8116 64592
rect 7699 64552 8116 64580
rect 7699 64549 7711 64552
rect 7653 64543 7711 64549
rect 8110 64540 8116 64552
rect 8168 64540 8174 64592
rect 32398 64580 32404 64592
rect 16546 64552 32404 64580
rect 8297 64515 8355 64521
rect 8297 64481 8309 64515
rect 8343 64512 8355 64515
rect 13446 64512 13452 64524
rect 8343 64484 13452 64512
rect 8343 64481 8355 64484
rect 8297 64475 8355 64481
rect 13446 64472 13452 64484
rect 13504 64512 13510 64524
rect 16546 64512 16574 64552
rect 32398 64540 32404 64552
rect 32456 64540 32462 64592
rect 13504 64484 16574 64512
rect 13504 64472 13510 64484
rect 20162 64472 20168 64524
rect 20220 64472 20226 64524
rect 31478 64512 31484 64524
rect 20272 64484 31484 64512
rect 7834 64404 7840 64456
rect 7892 64404 7898 64456
rect 8205 64447 8263 64453
rect 8205 64413 8217 64447
rect 8251 64444 8263 64447
rect 13538 64444 13544 64456
rect 8251 64416 13544 64444
rect 8251 64413 8263 64416
rect 8205 64407 8263 64413
rect 13538 64404 13544 64416
rect 13596 64444 13602 64456
rect 13596 64416 16574 64444
rect 13596 64404 13602 64416
rect 16546 64308 16574 64416
rect 19242 64404 19248 64456
rect 19300 64444 19306 64456
rect 20073 64447 20131 64453
rect 20073 64444 20085 64447
rect 19300 64416 20085 64444
rect 19300 64404 19306 64416
rect 20073 64413 20085 64416
rect 20119 64444 20131 64447
rect 20272 64444 20300 64484
rect 31478 64472 31484 64484
rect 31536 64472 31542 64524
rect 20119 64416 20300 64444
rect 20119 64413 20131 64416
rect 20073 64407 20131 64413
rect 20346 64404 20352 64456
rect 20404 64404 20410 64456
rect 20441 64447 20499 64453
rect 20441 64413 20453 64447
rect 20487 64413 20499 64447
rect 20441 64407 20499 64413
rect 17310 64336 17316 64388
rect 17368 64376 17374 64388
rect 20456 64376 20484 64407
rect 20714 64404 20720 64456
rect 20772 64404 20778 64456
rect 21082 64404 21088 64456
rect 21140 64404 21146 64456
rect 21726 64404 21732 64456
rect 21784 64404 21790 64456
rect 33686 64404 33692 64456
rect 33744 64404 33750 64456
rect 33965 64447 34023 64453
rect 33965 64413 33977 64447
rect 34011 64444 34023 64447
rect 36722 64444 36728 64456
rect 34011 64416 36728 64444
rect 34011 64413 34023 64416
rect 33965 64407 34023 64413
rect 36722 64404 36728 64416
rect 36780 64404 36786 64456
rect 17368 64348 20484 64376
rect 17368 64336 17374 64348
rect 33594 64336 33600 64388
rect 33652 64336 33658 64388
rect 20254 64308 20260 64320
rect 16546 64280 20260 64308
rect 20254 64268 20260 64280
rect 20312 64268 20318 64320
rect 20625 64311 20683 64317
rect 20625 64277 20637 64311
rect 20671 64308 20683 64311
rect 24394 64308 24400 64320
rect 20671 64280 24400 64308
rect 20671 64277 20683 64280
rect 20625 64271 20683 64277
rect 24394 64268 24400 64280
rect 24452 64268 24458 64320
rect 1104 64218 40848 64240
rect 1104 64166 2610 64218
rect 2662 64166 2674 64218
rect 2726 64166 2738 64218
rect 2790 64166 2802 64218
rect 2854 64166 2866 64218
rect 2918 64166 7610 64218
rect 7662 64166 7674 64218
rect 7726 64166 7738 64218
rect 7790 64166 7802 64218
rect 7854 64166 7866 64218
rect 7918 64166 12610 64218
rect 12662 64166 12674 64218
rect 12726 64166 12738 64218
rect 12790 64166 12802 64218
rect 12854 64166 12866 64218
rect 12918 64166 17610 64218
rect 17662 64166 17674 64218
rect 17726 64166 17738 64218
rect 17790 64166 17802 64218
rect 17854 64166 17866 64218
rect 17918 64166 22610 64218
rect 22662 64166 22674 64218
rect 22726 64166 22738 64218
rect 22790 64166 22802 64218
rect 22854 64166 22866 64218
rect 22918 64166 27610 64218
rect 27662 64166 27674 64218
rect 27726 64166 27738 64218
rect 27790 64166 27802 64218
rect 27854 64166 27866 64218
rect 27918 64166 32610 64218
rect 32662 64166 32674 64218
rect 32726 64166 32738 64218
rect 32790 64166 32802 64218
rect 32854 64166 32866 64218
rect 32918 64166 37610 64218
rect 37662 64166 37674 64218
rect 37726 64166 37738 64218
rect 37790 64166 37802 64218
rect 37854 64166 37866 64218
rect 37918 64166 40848 64218
rect 1104 64144 40848 64166
rect 15102 63996 15108 64048
rect 15160 64036 15166 64048
rect 20714 64036 20720 64048
rect 15160 64008 20720 64036
rect 15160 63996 15166 64008
rect 20714 63996 20720 64008
rect 20772 63996 20778 64048
rect 35250 63996 35256 64048
rect 35308 64036 35314 64048
rect 35308 64008 37964 64036
rect 35308 63996 35314 64008
rect 36354 63928 36360 63980
rect 36412 63968 36418 63980
rect 37936 63977 37964 64008
rect 37737 63971 37795 63977
rect 37737 63968 37749 63971
rect 36412 63940 37749 63968
rect 36412 63928 36418 63940
rect 37737 63937 37749 63940
rect 37783 63937 37795 63971
rect 37737 63931 37795 63937
rect 37921 63971 37979 63977
rect 37921 63937 37933 63971
rect 37967 63937 37979 63971
rect 37921 63931 37979 63937
rect 38102 63928 38108 63980
rect 38160 63928 38166 63980
rect 37277 63903 37335 63909
rect 37277 63869 37289 63903
rect 37323 63869 37335 63903
rect 37277 63863 37335 63869
rect 30190 63792 30196 63844
rect 30248 63832 30254 63844
rect 37292 63832 37320 63863
rect 37366 63860 37372 63912
rect 37424 63900 37430 63912
rect 38120 63900 38148 63928
rect 37424 63872 38148 63900
rect 37424 63860 37430 63872
rect 30248 63804 37320 63832
rect 30248 63792 30254 63804
rect 1104 63674 40848 63696
rect 1104 63622 1950 63674
rect 2002 63622 2014 63674
rect 2066 63622 2078 63674
rect 2130 63622 2142 63674
rect 2194 63622 2206 63674
rect 2258 63622 6950 63674
rect 7002 63622 7014 63674
rect 7066 63622 7078 63674
rect 7130 63622 7142 63674
rect 7194 63622 7206 63674
rect 7258 63622 11950 63674
rect 12002 63622 12014 63674
rect 12066 63622 12078 63674
rect 12130 63622 12142 63674
rect 12194 63622 12206 63674
rect 12258 63622 16950 63674
rect 17002 63622 17014 63674
rect 17066 63622 17078 63674
rect 17130 63622 17142 63674
rect 17194 63622 17206 63674
rect 17258 63622 21950 63674
rect 22002 63622 22014 63674
rect 22066 63622 22078 63674
rect 22130 63622 22142 63674
rect 22194 63622 22206 63674
rect 22258 63622 26950 63674
rect 27002 63622 27014 63674
rect 27066 63622 27078 63674
rect 27130 63622 27142 63674
rect 27194 63622 27206 63674
rect 27258 63622 31950 63674
rect 32002 63622 32014 63674
rect 32066 63622 32078 63674
rect 32130 63622 32142 63674
rect 32194 63622 32206 63674
rect 32258 63622 36950 63674
rect 37002 63622 37014 63674
rect 37066 63622 37078 63674
rect 37130 63622 37142 63674
rect 37194 63622 37206 63674
rect 37258 63622 40848 63674
rect 1104 63600 40848 63622
rect 16390 63520 16396 63572
rect 16448 63560 16454 63572
rect 26973 63563 27031 63569
rect 26973 63560 26985 63563
rect 16448 63532 26985 63560
rect 16448 63520 16454 63532
rect 26973 63529 26985 63532
rect 27019 63560 27031 63563
rect 27341 63563 27399 63569
rect 27341 63560 27353 63563
rect 27019 63532 27353 63560
rect 27019 63529 27031 63532
rect 26973 63523 27031 63529
rect 27341 63529 27353 63532
rect 27387 63529 27399 63563
rect 27341 63523 27399 63529
rect 34790 63520 34796 63572
rect 34848 63560 34854 63572
rect 35250 63560 35256 63572
rect 34848 63532 35256 63560
rect 34848 63520 34854 63532
rect 35250 63520 35256 63532
rect 35308 63520 35314 63572
rect 22370 63384 22376 63436
rect 22428 63424 22434 63436
rect 22428 63396 27936 63424
rect 22428 63384 22434 63396
rect 27908 63365 27936 63396
rect 27525 63359 27583 63365
rect 27525 63325 27537 63359
rect 27571 63325 27583 63359
rect 27525 63319 27583 63325
rect 27893 63359 27951 63365
rect 27893 63325 27905 63359
rect 27939 63356 27951 63359
rect 29730 63356 29736 63368
rect 27939 63328 29736 63356
rect 27939 63325 27951 63328
rect 27893 63319 27951 63325
rect 26694 63248 26700 63300
rect 26752 63288 26758 63300
rect 27540 63288 27568 63319
rect 29730 63316 29736 63328
rect 29788 63316 29794 63368
rect 35434 63288 35440 63300
rect 26752 63260 35440 63288
rect 26752 63248 26758 63260
rect 35434 63248 35440 63260
rect 35492 63248 35498 63300
rect 17865 63223 17923 63229
rect 17865 63189 17877 63223
rect 17911 63220 17923 63223
rect 17954 63220 17960 63232
rect 17911 63192 17960 63220
rect 17911 63189 17923 63192
rect 17865 63183 17923 63189
rect 17954 63180 17960 63192
rect 18012 63180 18018 63232
rect 27709 63223 27767 63229
rect 27709 63189 27721 63223
rect 27755 63220 27767 63223
rect 27982 63220 27988 63232
rect 27755 63192 27988 63220
rect 27755 63189 27767 63192
rect 27709 63183 27767 63189
rect 27982 63180 27988 63192
rect 28040 63180 28046 63232
rect 1104 63130 40848 63152
rect 1104 63078 2610 63130
rect 2662 63078 2674 63130
rect 2726 63078 2738 63130
rect 2790 63078 2802 63130
rect 2854 63078 2866 63130
rect 2918 63078 7610 63130
rect 7662 63078 7674 63130
rect 7726 63078 7738 63130
rect 7790 63078 7802 63130
rect 7854 63078 7866 63130
rect 7918 63078 12610 63130
rect 12662 63078 12674 63130
rect 12726 63078 12738 63130
rect 12790 63078 12802 63130
rect 12854 63078 12866 63130
rect 12918 63078 17610 63130
rect 17662 63078 17674 63130
rect 17726 63078 17738 63130
rect 17790 63078 17802 63130
rect 17854 63078 17866 63130
rect 17918 63078 22610 63130
rect 22662 63078 22674 63130
rect 22726 63078 22738 63130
rect 22790 63078 22802 63130
rect 22854 63078 22866 63130
rect 22918 63078 27610 63130
rect 27662 63078 27674 63130
rect 27726 63078 27738 63130
rect 27790 63078 27802 63130
rect 27854 63078 27866 63130
rect 27918 63078 32610 63130
rect 32662 63078 32674 63130
rect 32726 63078 32738 63130
rect 32790 63078 32802 63130
rect 32854 63078 32866 63130
rect 32918 63078 37610 63130
rect 37662 63078 37674 63130
rect 37726 63078 37738 63130
rect 37790 63078 37802 63130
rect 37854 63078 37866 63130
rect 37918 63078 40848 63130
rect 1104 63056 40848 63078
rect 16298 62976 16304 63028
rect 16356 63016 16362 63028
rect 18233 63019 18291 63025
rect 18233 63016 18245 63019
rect 16356 62988 18245 63016
rect 16356 62976 16362 62988
rect 18233 62985 18245 62988
rect 18279 62985 18291 63019
rect 18233 62979 18291 62985
rect 14642 62908 14648 62960
rect 14700 62948 14706 62960
rect 30282 62948 30288 62960
rect 14700 62920 30288 62948
rect 14700 62908 14706 62920
rect 30282 62908 30288 62920
rect 30340 62908 30346 62960
rect 6822 62840 6828 62892
rect 6880 62880 6886 62892
rect 8113 62883 8171 62889
rect 8113 62880 8125 62883
rect 6880 62852 8125 62880
rect 6880 62840 6886 62852
rect 8113 62849 8125 62852
rect 8159 62849 8171 62883
rect 8113 62843 8171 62849
rect 8297 62883 8355 62889
rect 8297 62849 8309 62883
rect 8343 62880 8355 62883
rect 10870 62880 10876 62892
rect 8343 62852 10876 62880
rect 8343 62849 8355 62852
rect 8297 62843 8355 62849
rect 10870 62840 10876 62852
rect 10928 62840 10934 62892
rect 18295 62883 18353 62889
rect 18295 62849 18307 62883
rect 18341 62880 18353 62883
rect 19978 62880 19984 62892
rect 18341 62852 19984 62880
rect 18341 62849 18353 62852
rect 18295 62843 18353 62849
rect 19978 62840 19984 62852
rect 20036 62840 20042 62892
rect 1854 62772 1860 62824
rect 1912 62812 1918 62824
rect 8938 62812 8944 62824
rect 1912 62784 8944 62812
rect 1912 62772 1918 62784
rect 8938 62772 8944 62784
rect 8996 62772 9002 62824
rect 16574 62772 16580 62824
rect 16632 62812 16638 62824
rect 17773 62815 17831 62821
rect 17773 62812 17785 62815
rect 16632 62784 17785 62812
rect 16632 62772 16638 62784
rect 17773 62781 17785 62784
rect 17819 62781 17831 62815
rect 17773 62775 17831 62781
rect 4890 62704 4896 62756
rect 4948 62744 4954 62756
rect 4948 62716 11744 62744
rect 4948 62704 4954 62716
rect 8481 62679 8539 62685
rect 8481 62645 8493 62679
rect 8527 62676 8539 62679
rect 9582 62676 9588 62688
rect 8527 62648 9588 62676
rect 8527 62645 8539 62648
rect 8481 62639 8539 62645
rect 9582 62636 9588 62648
rect 9640 62636 9646 62688
rect 11716 62676 11744 62716
rect 13354 62704 13360 62756
rect 13412 62744 13418 62756
rect 25038 62744 25044 62756
rect 13412 62716 25044 62744
rect 13412 62704 13418 62716
rect 25038 62704 25044 62716
rect 25096 62704 25102 62756
rect 17865 62679 17923 62685
rect 17865 62676 17877 62679
rect 11716 62648 17877 62676
rect 17865 62645 17877 62648
rect 17911 62645 17923 62679
rect 17865 62639 17923 62645
rect 17954 62636 17960 62688
rect 18012 62676 18018 62688
rect 18417 62679 18475 62685
rect 18417 62676 18429 62679
rect 18012 62648 18429 62676
rect 18012 62636 18018 62648
rect 18417 62645 18429 62648
rect 18463 62645 18475 62679
rect 18417 62639 18475 62645
rect 1104 62586 40848 62608
rect 1104 62534 1950 62586
rect 2002 62534 2014 62586
rect 2066 62534 2078 62586
rect 2130 62534 2142 62586
rect 2194 62534 2206 62586
rect 2258 62534 6950 62586
rect 7002 62534 7014 62586
rect 7066 62534 7078 62586
rect 7130 62534 7142 62586
rect 7194 62534 7206 62586
rect 7258 62534 11950 62586
rect 12002 62534 12014 62586
rect 12066 62534 12078 62586
rect 12130 62534 12142 62586
rect 12194 62534 12206 62586
rect 12258 62534 16950 62586
rect 17002 62534 17014 62586
rect 17066 62534 17078 62586
rect 17130 62534 17142 62586
rect 17194 62534 17206 62586
rect 17258 62534 21950 62586
rect 22002 62534 22014 62586
rect 22066 62534 22078 62586
rect 22130 62534 22142 62586
rect 22194 62534 22206 62586
rect 22258 62534 26950 62586
rect 27002 62534 27014 62586
rect 27066 62534 27078 62586
rect 27130 62534 27142 62586
rect 27194 62534 27206 62586
rect 27258 62534 31950 62586
rect 32002 62534 32014 62586
rect 32066 62534 32078 62586
rect 32130 62534 32142 62586
rect 32194 62534 32206 62586
rect 32258 62534 36950 62586
rect 37002 62534 37014 62586
rect 37066 62534 37078 62586
rect 37130 62534 37142 62586
rect 37194 62534 37206 62586
rect 37258 62534 40848 62586
rect 1104 62512 40848 62534
rect 12894 62432 12900 62484
rect 12952 62472 12958 62484
rect 27430 62472 27436 62484
rect 12952 62444 27436 62472
rect 12952 62432 12958 62444
rect 27430 62432 27436 62444
rect 27488 62432 27494 62484
rect 7576 62376 18092 62404
rect 7374 62228 7380 62280
rect 7432 62228 7438 62280
rect 7576 62277 7604 62376
rect 13265 62339 13323 62345
rect 13265 62305 13277 62339
rect 13311 62336 13323 62339
rect 15102 62336 15108 62348
rect 13311 62308 15108 62336
rect 13311 62305 13323 62308
rect 13265 62299 13323 62305
rect 15102 62296 15108 62308
rect 15160 62296 15166 62348
rect 7561 62271 7619 62277
rect 7561 62237 7573 62271
rect 7607 62237 7619 62271
rect 7561 62231 7619 62237
rect 12161 62271 12219 62277
rect 12161 62237 12173 62271
rect 12207 62237 12219 62271
rect 12161 62231 12219 62237
rect 4430 62092 4436 62144
rect 4488 62132 4494 62144
rect 7469 62135 7527 62141
rect 7469 62132 7481 62135
rect 4488 62104 7481 62132
rect 4488 62092 4494 62104
rect 7469 62101 7481 62104
rect 7515 62101 7527 62135
rect 12176 62132 12204 62231
rect 12526 62228 12532 62280
rect 12584 62228 12590 62280
rect 12894 62228 12900 62280
rect 12952 62228 12958 62280
rect 13354 62228 13360 62280
rect 13412 62228 13418 62280
rect 13262 62132 13268 62144
rect 12176 62104 13268 62132
rect 7469 62095 7527 62101
rect 13262 62092 13268 62104
rect 13320 62132 13326 62144
rect 13906 62132 13912 62144
rect 13320 62104 13912 62132
rect 13320 62092 13326 62104
rect 13906 62092 13912 62104
rect 13964 62092 13970 62144
rect 17865 62135 17923 62141
rect 17865 62101 17877 62135
rect 17911 62132 17923 62135
rect 17954 62132 17960 62144
rect 17911 62104 17960 62132
rect 17911 62101 17923 62104
rect 17865 62095 17923 62101
rect 17954 62092 17960 62104
rect 18012 62092 18018 62144
rect 18064 62132 18092 62376
rect 18138 62364 18144 62416
rect 18196 62404 18202 62416
rect 20165 62407 20223 62413
rect 20165 62404 20177 62407
rect 18196 62376 20177 62404
rect 18196 62364 18202 62376
rect 20165 62373 20177 62376
rect 20211 62404 20223 62407
rect 28994 62404 29000 62416
rect 20211 62376 29000 62404
rect 20211 62373 20223 62376
rect 20165 62367 20223 62373
rect 28994 62364 29000 62376
rect 29052 62404 29058 62416
rect 30190 62404 30196 62416
rect 29052 62376 30196 62404
rect 29052 62364 29058 62376
rect 30190 62364 30196 62376
rect 30248 62364 30254 62416
rect 18230 62296 18236 62348
rect 18288 62336 18294 62348
rect 18288 62308 20484 62336
rect 18288 62296 18294 62308
rect 20456 62277 20484 62308
rect 30282 62296 30288 62348
rect 30340 62336 30346 62348
rect 34701 62339 34759 62345
rect 34701 62336 34713 62339
rect 30340 62308 34713 62336
rect 30340 62296 30346 62308
rect 34701 62305 34713 62308
rect 34747 62305 34759 62339
rect 34701 62299 34759 62305
rect 20441 62271 20499 62277
rect 20441 62237 20453 62271
rect 20487 62268 20499 62271
rect 28258 62268 28264 62280
rect 20487 62240 28264 62268
rect 20487 62237 20499 62240
rect 20441 62231 20499 62237
rect 28258 62228 28264 62240
rect 28316 62228 28322 62280
rect 30650 62228 30656 62280
rect 30708 62268 30714 62280
rect 34885 62271 34943 62277
rect 34885 62268 34897 62271
rect 30708 62240 34897 62268
rect 30708 62228 30714 62240
rect 34885 62237 34897 62240
rect 34931 62237 34943 62271
rect 34885 62231 34943 62237
rect 35250 62228 35256 62280
rect 35308 62228 35314 62280
rect 35618 62228 35624 62280
rect 35676 62228 35682 62280
rect 20070 62160 20076 62212
rect 20128 62200 20134 62212
rect 20346 62200 20352 62212
rect 20128 62172 20352 62200
rect 20128 62160 20134 62172
rect 20346 62160 20352 62172
rect 20404 62160 20410 62212
rect 20898 62160 20904 62212
rect 20956 62160 20962 62212
rect 23198 62132 23204 62144
rect 18064 62104 23204 62132
rect 23198 62092 23204 62104
rect 23256 62132 23262 62144
rect 23382 62132 23388 62144
rect 23256 62104 23388 62132
rect 23256 62092 23262 62104
rect 23382 62092 23388 62104
rect 23440 62092 23446 62144
rect 1104 62042 40848 62064
rect 1104 61990 2610 62042
rect 2662 61990 2674 62042
rect 2726 61990 2738 62042
rect 2790 61990 2802 62042
rect 2854 61990 2866 62042
rect 2918 61990 7610 62042
rect 7662 61990 7674 62042
rect 7726 61990 7738 62042
rect 7790 61990 7802 62042
rect 7854 61990 7866 62042
rect 7918 61990 12610 62042
rect 12662 61990 12674 62042
rect 12726 61990 12738 62042
rect 12790 61990 12802 62042
rect 12854 61990 12866 62042
rect 12918 61990 17610 62042
rect 17662 61990 17674 62042
rect 17726 61990 17738 62042
rect 17790 61990 17802 62042
rect 17854 61990 17866 62042
rect 17918 61990 22610 62042
rect 22662 61990 22674 62042
rect 22726 61990 22738 62042
rect 22790 61990 22802 62042
rect 22854 61990 22866 62042
rect 22918 61990 27610 62042
rect 27662 61990 27674 62042
rect 27726 61990 27738 62042
rect 27790 61990 27802 62042
rect 27854 61990 27866 62042
rect 27918 61990 32610 62042
rect 32662 61990 32674 62042
rect 32726 61990 32738 62042
rect 32790 61990 32802 62042
rect 32854 61990 32866 62042
rect 32918 61990 37610 62042
rect 37662 61990 37674 62042
rect 37726 61990 37738 62042
rect 37790 61990 37802 62042
rect 37854 61990 37866 62042
rect 37918 61990 40848 62042
rect 1104 61968 40848 61990
rect 13265 61795 13323 61801
rect 13265 61761 13277 61795
rect 13311 61792 13323 61795
rect 13814 61792 13820 61804
rect 13311 61764 13820 61792
rect 13311 61761 13323 61764
rect 13265 61755 13323 61761
rect 13814 61752 13820 61764
rect 13872 61752 13878 61804
rect 11790 61684 11796 61736
rect 11848 61724 11854 61736
rect 13173 61727 13231 61733
rect 13173 61724 13185 61727
rect 11848 61696 13185 61724
rect 11848 61684 11854 61696
rect 13173 61693 13185 61696
rect 13219 61693 13231 61727
rect 13173 61687 13231 61693
rect 13722 61684 13728 61736
rect 13780 61684 13786 61736
rect 17865 61591 17923 61597
rect 17865 61557 17877 61591
rect 17911 61588 17923 61591
rect 17954 61588 17960 61600
rect 17911 61560 17960 61588
rect 17911 61557 17923 61560
rect 17865 61551 17923 61557
rect 17954 61548 17960 61560
rect 18012 61588 18018 61600
rect 18782 61588 18788 61600
rect 18012 61560 18788 61588
rect 18012 61548 18018 61560
rect 18782 61548 18788 61560
rect 18840 61548 18846 61600
rect 1104 61498 40848 61520
rect 1104 61446 1950 61498
rect 2002 61446 2014 61498
rect 2066 61446 2078 61498
rect 2130 61446 2142 61498
rect 2194 61446 2206 61498
rect 2258 61446 6950 61498
rect 7002 61446 7014 61498
rect 7066 61446 7078 61498
rect 7130 61446 7142 61498
rect 7194 61446 7206 61498
rect 7258 61446 11950 61498
rect 12002 61446 12014 61498
rect 12066 61446 12078 61498
rect 12130 61446 12142 61498
rect 12194 61446 12206 61498
rect 12258 61446 16950 61498
rect 17002 61446 17014 61498
rect 17066 61446 17078 61498
rect 17130 61446 17142 61498
rect 17194 61446 17206 61498
rect 17258 61446 21950 61498
rect 22002 61446 22014 61498
rect 22066 61446 22078 61498
rect 22130 61446 22142 61498
rect 22194 61446 22206 61498
rect 22258 61446 26950 61498
rect 27002 61446 27014 61498
rect 27066 61446 27078 61498
rect 27130 61446 27142 61498
rect 27194 61446 27206 61498
rect 27258 61446 31950 61498
rect 32002 61446 32014 61498
rect 32066 61446 32078 61498
rect 32130 61446 32142 61498
rect 32194 61446 32206 61498
rect 32258 61446 36950 61498
rect 37002 61446 37014 61498
rect 37066 61446 37078 61498
rect 37130 61446 37142 61498
rect 37194 61446 37206 61498
rect 37258 61446 40848 61498
rect 1104 61424 40848 61446
rect 13906 61344 13912 61396
rect 13964 61384 13970 61396
rect 36538 61384 36544 61396
rect 13964 61356 36544 61384
rect 13964 61344 13970 61356
rect 36538 61344 36544 61356
rect 36596 61344 36602 61396
rect 1412 61288 16574 61316
rect 1412 61180 1440 61288
rect 1489 61251 1547 61257
rect 1489 61217 1501 61251
rect 1535 61248 1547 61251
rect 16546 61248 16574 61288
rect 17954 61248 17960 61260
rect 1535 61220 9536 61248
rect 16546 61220 17960 61248
rect 1535 61217 1547 61220
rect 1489 61211 1547 61217
rect 1581 61183 1639 61189
rect 1581 61180 1593 61183
rect 1412 61152 1593 61180
rect 1581 61149 1593 61152
rect 1627 61149 1639 61183
rect 1581 61143 1639 61149
rect 2409 61183 2467 61189
rect 2409 61149 2421 61183
rect 2455 61180 2467 61183
rect 2498 61180 2504 61192
rect 2455 61152 2504 61180
rect 2455 61149 2467 61152
rect 2409 61143 2467 61149
rect 2498 61140 2504 61152
rect 2556 61140 2562 61192
rect 4249 61183 4307 61189
rect 4249 61149 4261 61183
rect 4295 61180 4307 61183
rect 5534 61180 5540 61192
rect 4295 61152 5540 61180
rect 4295 61149 4307 61152
rect 4249 61143 4307 61149
rect 5534 61140 5540 61152
rect 5592 61140 5598 61192
rect 8938 61140 8944 61192
rect 8996 61140 9002 61192
rect 9214 61140 9220 61192
rect 9272 61140 9278 61192
rect 9508 61180 9536 61220
rect 17954 61208 17960 61220
rect 18012 61248 18018 61260
rect 19242 61248 19248 61260
rect 18012 61220 19248 61248
rect 18012 61208 18018 61220
rect 19242 61208 19248 61220
rect 19300 61208 19306 61260
rect 33870 61180 33876 61192
rect 9508 61152 33876 61180
rect 33870 61140 33876 61152
rect 33928 61140 33934 61192
rect 2314 61072 2320 61124
rect 2372 61072 2378 61124
rect 3694 61072 3700 61124
rect 3752 61112 3758 61124
rect 4065 61115 4123 61121
rect 4065 61112 4077 61115
rect 3752 61084 4077 61112
rect 3752 61072 3758 61084
rect 4065 61081 4077 61084
rect 4111 61081 4123 61115
rect 4065 61075 4123 61081
rect 4157 61115 4215 61121
rect 4157 61081 4169 61115
rect 4203 61112 4215 61115
rect 4433 61115 4491 61121
rect 4203 61084 4384 61112
rect 4203 61081 4215 61084
rect 4157 61075 4215 61081
rect 3878 61004 3884 61056
rect 3936 61004 3942 61056
rect 4356 61044 4384 61084
rect 4433 61081 4445 61115
rect 4479 61112 4491 61115
rect 4706 61112 4712 61124
rect 4479 61084 4712 61112
rect 4479 61081 4491 61084
rect 4433 61075 4491 61081
rect 4706 61072 4712 61084
rect 4764 61072 4770 61124
rect 8018 61072 8024 61124
rect 8076 61112 8082 61124
rect 9125 61115 9183 61121
rect 9125 61112 9137 61115
rect 8076 61084 9137 61112
rect 8076 61072 8082 61084
rect 9125 61081 9137 61084
rect 9171 61081 9183 61115
rect 9125 61075 9183 61081
rect 9677 61115 9735 61121
rect 9677 61081 9689 61115
rect 9723 61112 9735 61115
rect 10318 61112 10324 61124
rect 9723 61084 10324 61112
rect 9723 61081 9735 61084
rect 9677 61075 9735 61081
rect 10318 61072 10324 61084
rect 10376 61072 10382 61124
rect 4798 61044 4804 61056
rect 4356 61016 4804 61044
rect 4798 61004 4804 61016
rect 4856 61004 4862 61056
rect 1104 60954 40848 60976
rect 1104 60902 2610 60954
rect 2662 60902 2674 60954
rect 2726 60902 2738 60954
rect 2790 60902 2802 60954
rect 2854 60902 2866 60954
rect 2918 60902 7610 60954
rect 7662 60902 7674 60954
rect 7726 60902 7738 60954
rect 7790 60902 7802 60954
rect 7854 60902 7866 60954
rect 7918 60902 12610 60954
rect 12662 60902 12674 60954
rect 12726 60902 12738 60954
rect 12790 60902 12802 60954
rect 12854 60902 12866 60954
rect 12918 60902 17610 60954
rect 17662 60902 17674 60954
rect 17726 60902 17738 60954
rect 17790 60902 17802 60954
rect 17854 60902 17866 60954
rect 17918 60902 22610 60954
rect 22662 60902 22674 60954
rect 22726 60902 22738 60954
rect 22790 60902 22802 60954
rect 22854 60902 22866 60954
rect 22918 60902 27610 60954
rect 27662 60902 27674 60954
rect 27726 60902 27738 60954
rect 27790 60902 27802 60954
rect 27854 60902 27866 60954
rect 27918 60902 32610 60954
rect 32662 60902 32674 60954
rect 32726 60902 32738 60954
rect 32790 60902 32802 60954
rect 32854 60902 32866 60954
rect 32918 60902 37610 60954
rect 37662 60902 37674 60954
rect 37726 60902 37738 60954
rect 37790 60902 37802 60954
rect 37854 60902 37866 60954
rect 37918 60902 40848 60954
rect 1104 60880 40848 60902
rect 4798 60732 4804 60784
rect 4856 60772 4862 60784
rect 10686 60772 10692 60784
rect 4856 60744 10692 60772
rect 4856 60732 4862 60744
rect 10686 60732 10692 60744
rect 10744 60732 10750 60784
rect 1670 60664 1676 60716
rect 1728 60704 1734 60716
rect 8113 60707 8171 60713
rect 8113 60704 8125 60707
rect 1728 60676 8125 60704
rect 1728 60664 1734 60676
rect 8113 60673 8125 60676
rect 8159 60673 8171 60707
rect 8113 60667 8171 60673
rect 8478 60664 8484 60716
rect 8536 60664 8542 60716
rect 9030 60704 9036 60716
rect 8588 60676 9036 60704
rect 5534 60596 5540 60648
rect 5592 60636 5598 60648
rect 8205 60639 8263 60645
rect 8205 60636 8217 60639
rect 5592 60608 8217 60636
rect 5592 60596 5598 60608
rect 8205 60605 8217 60608
rect 8251 60636 8263 60639
rect 8588 60636 8616 60676
rect 9030 60664 9036 60676
rect 9088 60664 9094 60716
rect 18598 60664 18604 60716
rect 18656 60704 18662 60716
rect 28997 60707 29055 60713
rect 28997 60704 29009 60707
rect 18656 60676 29009 60704
rect 18656 60664 18662 60676
rect 28997 60673 29009 60676
rect 29043 60673 29055 60707
rect 28997 60667 29055 60673
rect 29546 60664 29552 60716
rect 29604 60664 29610 60716
rect 38654 60664 38660 60716
rect 38712 60664 38718 60716
rect 38746 60664 38752 60716
rect 38804 60664 38810 60716
rect 38933 60707 38991 60713
rect 38933 60673 38945 60707
rect 38979 60673 38991 60707
rect 38933 60667 38991 60673
rect 8251 60608 8616 60636
rect 8665 60639 8723 60645
rect 8251 60605 8263 60608
rect 8205 60599 8263 60605
rect 8665 60605 8677 60639
rect 8711 60636 8723 60639
rect 38838 60636 38844 60648
rect 8711 60608 38844 60636
rect 8711 60605 8723 60608
rect 8665 60599 8723 60605
rect 8680 60568 8708 60599
rect 38838 60596 38844 60608
rect 38896 60596 38902 60648
rect 38289 60571 38347 60577
rect 38289 60568 38301 60571
rect 5552 60540 8708 60568
rect 8772 60540 38301 60568
rect 5552 60512 5580 60540
rect 5534 60460 5540 60512
rect 5592 60460 5598 60512
rect 8110 60460 8116 60512
rect 8168 60500 8174 60512
rect 8772 60500 8800 60540
rect 38289 60537 38301 60540
rect 38335 60568 38347 60571
rect 38948 60568 38976 60667
rect 38335 60540 38976 60568
rect 38335 60537 38347 60540
rect 38289 60531 38347 60537
rect 8168 60472 8800 60500
rect 8168 60460 8174 60472
rect 8846 60460 8852 60512
rect 8904 60460 8910 60512
rect 19337 60503 19395 60509
rect 19337 60469 19349 60503
rect 19383 60500 19395 60503
rect 19702 60500 19708 60512
rect 19383 60472 19708 60500
rect 19383 60469 19395 60472
rect 19337 60463 19395 60469
rect 19702 60460 19708 60472
rect 19760 60460 19766 60512
rect 29086 60460 29092 60512
rect 29144 60460 29150 60512
rect 39114 60460 39120 60512
rect 39172 60460 39178 60512
rect 1104 60410 40848 60432
rect 1104 60358 1950 60410
rect 2002 60358 2014 60410
rect 2066 60358 2078 60410
rect 2130 60358 2142 60410
rect 2194 60358 2206 60410
rect 2258 60358 6950 60410
rect 7002 60358 7014 60410
rect 7066 60358 7078 60410
rect 7130 60358 7142 60410
rect 7194 60358 7206 60410
rect 7258 60358 11950 60410
rect 12002 60358 12014 60410
rect 12066 60358 12078 60410
rect 12130 60358 12142 60410
rect 12194 60358 12206 60410
rect 12258 60358 16950 60410
rect 17002 60358 17014 60410
rect 17066 60358 17078 60410
rect 17130 60358 17142 60410
rect 17194 60358 17206 60410
rect 17258 60358 21950 60410
rect 22002 60358 22014 60410
rect 22066 60358 22078 60410
rect 22130 60358 22142 60410
rect 22194 60358 22206 60410
rect 22258 60358 26950 60410
rect 27002 60358 27014 60410
rect 27066 60358 27078 60410
rect 27130 60358 27142 60410
rect 27194 60358 27206 60410
rect 27258 60358 31950 60410
rect 32002 60358 32014 60410
rect 32066 60358 32078 60410
rect 32130 60358 32142 60410
rect 32194 60358 32206 60410
rect 32258 60358 36950 60410
rect 37002 60358 37014 60410
rect 37066 60358 37078 60410
rect 37130 60358 37142 60410
rect 37194 60358 37206 60410
rect 37258 60358 40848 60410
rect 1104 60336 40848 60358
rect 19610 60256 19616 60308
rect 19668 60256 19674 60308
rect 34698 60256 34704 60308
rect 34756 60256 34762 60308
rect 39114 60296 39120 60308
rect 35866 60268 39120 60296
rect 26206 60200 35020 60228
rect 6886 60132 21772 60160
rect 5994 60052 6000 60104
rect 6052 60092 6058 60104
rect 6886 60092 6914 60132
rect 6052 60064 6914 60092
rect 6052 60052 6058 60064
rect 19242 60052 19248 60104
rect 19300 60052 19306 60104
rect 21744 60101 21772 60132
rect 23842 60120 23848 60172
rect 23900 60160 23906 60172
rect 26206 60160 26234 60200
rect 23900 60132 26234 60160
rect 23900 60120 23906 60132
rect 29638 60120 29644 60172
rect 29696 60120 29702 60172
rect 21729 60095 21787 60101
rect 21729 60061 21741 60095
rect 21775 60061 21787 60095
rect 21729 60055 21787 60061
rect 22094 60052 22100 60104
rect 22152 60052 22158 60104
rect 22189 60095 22247 60101
rect 22189 60061 22201 60095
rect 22235 60092 22247 60095
rect 23106 60092 23112 60104
rect 22235 60064 23112 60092
rect 22235 60061 22247 60064
rect 22189 60055 22247 60061
rect 23106 60052 23112 60064
rect 23164 60052 23170 60104
rect 28902 60052 28908 60104
rect 28960 60092 28966 60104
rect 30193 60095 30251 60101
rect 30193 60092 30205 60095
rect 28960 60064 30205 60092
rect 28960 60052 28966 60064
rect 30193 60061 30205 60064
rect 30239 60061 30251 60095
rect 30193 60055 30251 60061
rect 21266 59984 21272 60036
rect 21324 59984 21330 60036
rect 30208 60024 30236 60055
rect 30926 60052 30932 60104
rect 30984 60092 30990 60104
rect 32677 60095 32735 60101
rect 32677 60092 32689 60095
rect 30984 60064 32689 60092
rect 30984 60052 30990 60064
rect 32677 60061 32689 60064
rect 32723 60061 32735 60095
rect 32677 60055 32735 60061
rect 33134 60052 33140 60104
rect 33192 60052 33198 60104
rect 33410 60052 33416 60104
rect 33468 60052 33474 60104
rect 33778 60052 33784 60104
rect 33836 60052 33842 60104
rect 34146 60052 34152 60104
rect 34204 60052 34210 60104
rect 34992 60101 35020 60200
rect 34977 60095 35035 60101
rect 34977 60061 34989 60095
rect 35023 60061 35035 60095
rect 34977 60055 35035 60061
rect 32585 60027 32643 60033
rect 32585 60024 32597 60027
rect 30208 59996 32597 60024
rect 32585 59993 32597 59996
rect 32631 59993 32643 60027
rect 32585 59987 32643 59993
rect 34698 59984 34704 60036
rect 34756 59984 34762 60036
rect 35866 60024 35894 60268
rect 39114 60256 39120 60268
rect 39172 60256 39178 60308
rect 34808 59996 35894 60024
rect 19613 59959 19671 59965
rect 19613 59925 19625 59959
rect 19659 59956 19671 59959
rect 19702 59956 19708 59968
rect 19659 59928 19708 59956
rect 19659 59925 19671 59928
rect 19613 59919 19671 59925
rect 19702 59916 19708 59928
rect 19760 59916 19766 59968
rect 19797 59959 19855 59965
rect 19797 59925 19809 59959
rect 19843 59956 19855 59959
rect 22462 59956 22468 59968
rect 19843 59928 22468 59956
rect 19843 59925 19855 59928
rect 19797 59919 19855 59925
rect 22462 59916 22468 59928
rect 22520 59916 22526 59968
rect 27522 59916 27528 59968
rect 27580 59956 27586 59968
rect 34808 59956 34836 59996
rect 27580 59928 34836 59956
rect 27580 59916 27586 59928
rect 34882 59916 34888 59968
rect 34940 59916 34946 59968
rect 1104 59866 40848 59888
rect 1104 59814 2610 59866
rect 2662 59814 2674 59866
rect 2726 59814 2738 59866
rect 2790 59814 2802 59866
rect 2854 59814 2866 59866
rect 2918 59814 7610 59866
rect 7662 59814 7674 59866
rect 7726 59814 7738 59866
rect 7790 59814 7802 59866
rect 7854 59814 7866 59866
rect 7918 59814 12610 59866
rect 12662 59814 12674 59866
rect 12726 59814 12738 59866
rect 12790 59814 12802 59866
rect 12854 59814 12866 59866
rect 12918 59814 17610 59866
rect 17662 59814 17674 59866
rect 17726 59814 17738 59866
rect 17790 59814 17802 59866
rect 17854 59814 17866 59866
rect 17918 59814 22610 59866
rect 22662 59814 22674 59866
rect 22726 59814 22738 59866
rect 22790 59814 22802 59866
rect 22854 59814 22866 59866
rect 22918 59814 27610 59866
rect 27662 59814 27674 59866
rect 27726 59814 27738 59866
rect 27790 59814 27802 59866
rect 27854 59814 27866 59866
rect 27918 59814 32610 59866
rect 32662 59814 32674 59866
rect 32726 59814 32738 59866
rect 32790 59814 32802 59866
rect 32854 59814 32866 59866
rect 32918 59814 37610 59866
rect 37662 59814 37674 59866
rect 37726 59814 37738 59866
rect 37790 59814 37802 59866
rect 37854 59814 37866 59866
rect 37918 59814 40848 59866
rect 1104 59792 40848 59814
rect 21266 59644 21272 59696
rect 21324 59684 21330 59696
rect 34882 59684 34888 59696
rect 21324 59656 34888 59684
rect 21324 59644 21330 59656
rect 34882 59644 34888 59656
rect 34940 59644 34946 59696
rect 39942 59576 39948 59628
rect 40000 59616 40006 59628
rect 40313 59619 40371 59625
rect 40313 59616 40325 59619
rect 40000 59588 40325 59616
rect 40000 59576 40006 59588
rect 40313 59585 40325 59588
rect 40359 59585 40371 59619
rect 40313 59579 40371 59585
rect 39666 59508 39672 59560
rect 39724 59508 39730 59560
rect 12526 59440 12532 59492
rect 12584 59480 12590 59492
rect 18506 59480 18512 59492
rect 12584 59452 18512 59480
rect 12584 59440 12590 59452
rect 18506 59440 18512 59452
rect 18564 59440 18570 59492
rect 18598 59372 18604 59424
rect 18656 59412 18662 59424
rect 19058 59412 19064 59424
rect 18656 59384 19064 59412
rect 18656 59372 18662 59384
rect 19058 59372 19064 59384
rect 19116 59372 19122 59424
rect 19337 59415 19395 59421
rect 19337 59381 19349 59415
rect 19383 59412 19395 59415
rect 19702 59412 19708 59424
rect 19383 59384 19708 59412
rect 19383 59381 19395 59384
rect 19337 59375 19395 59381
rect 19702 59372 19708 59384
rect 19760 59412 19766 59424
rect 21358 59412 21364 59424
rect 19760 59384 21364 59412
rect 19760 59372 19766 59384
rect 21358 59372 21364 59384
rect 21416 59372 21422 59424
rect 1104 59322 40848 59344
rect 1104 59270 1950 59322
rect 2002 59270 2014 59322
rect 2066 59270 2078 59322
rect 2130 59270 2142 59322
rect 2194 59270 2206 59322
rect 2258 59270 6950 59322
rect 7002 59270 7014 59322
rect 7066 59270 7078 59322
rect 7130 59270 7142 59322
rect 7194 59270 7206 59322
rect 7258 59270 11950 59322
rect 12002 59270 12014 59322
rect 12066 59270 12078 59322
rect 12130 59270 12142 59322
rect 12194 59270 12206 59322
rect 12258 59270 16950 59322
rect 17002 59270 17014 59322
rect 17066 59270 17078 59322
rect 17130 59270 17142 59322
rect 17194 59270 17206 59322
rect 17258 59270 21950 59322
rect 22002 59270 22014 59322
rect 22066 59270 22078 59322
rect 22130 59270 22142 59322
rect 22194 59270 22206 59322
rect 22258 59270 26950 59322
rect 27002 59270 27014 59322
rect 27066 59270 27078 59322
rect 27130 59270 27142 59322
rect 27194 59270 27206 59322
rect 27258 59270 31950 59322
rect 32002 59270 32014 59322
rect 32066 59270 32078 59322
rect 32130 59270 32142 59322
rect 32194 59270 32206 59322
rect 32258 59270 36950 59322
rect 37002 59270 37014 59322
rect 37066 59270 37078 59322
rect 37130 59270 37142 59322
rect 37194 59270 37206 59322
rect 37258 59270 40848 59322
rect 1104 59248 40848 59270
rect 26694 59208 26700 59220
rect 6886 59180 26700 59208
rect 6886 59140 6914 59180
rect 26694 59168 26700 59180
rect 26752 59168 26758 59220
rect 4356 59112 6914 59140
rect 7193 59143 7251 59149
rect 4356 59016 4384 59112
rect 7193 59109 7205 59143
rect 7239 59140 7251 59143
rect 7466 59140 7472 59152
rect 7239 59112 7472 59140
rect 7239 59109 7251 59112
rect 7193 59103 7251 59109
rect 7466 59100 7472 59112
rect 7524 59100 7530 59152
rect 4709 59075 4767 59081
rect 4709 59041 4721 59075
rect 4755 59072 4767 59075
rect 6362 59072 6368 59084
rect 4755 59044 6368 59072
rect 4755 59041 4767 59044
rect 4709 59035 4767 59041
rect 6362 59032 6368 59044
rect 6420 59032 6426 59084
rect 22370 59072 22376 59084
rect 6886 59044 22376 59072
rect 4338 58964 4344 59016
rect 4396 58964 4402 59016
rect 6730 58964 6736 59016
rect 6788 58964 6794 59016
rect 4157 58939 4215 58945
rect 4157 58905 4169 58939
rect 4203 58936 4215 58939
rect 4614 58936 4620 58948
rect 4203 58908 4620 58936
rect 4203 58905 4215 58908
rect 4157 58899 4215 58905
rect 4614 58896 4620 58908
rect 4672 58936 4678 58948
rect 6886 58936 6914 59044
rect 22370 59032 22376 59044
rect 22428 59032 22434 59084
rect 30929 59075 30987 59081
rect 30929 59072 30941 59075
rect 26206 59044 30941 59072
rect 22278 58964 22284 59016
rect 22336 59004 22342 59016
rect 22925 59007 22983 59013
rect 22925 59004 22937 59007
rect 22336 58976 22937 59004
rect 22336 58964 22342 58976
rect 22925 58973 22937 58976
rect 22971 58973 22983 59007
rect 22925 58967 22983 58973
rect 23201 59007 23259 59013
rect 23201 58973 23213 59007
rect 23247 59004 23259 59007
rect 23382 59004 23388 59016
rect 23247 58976 23388 59004
rect 23247 58973 23259 58976
rect 23201 58967 23259 58973
rect 23382 58964 23388 58976
rect 23440 58964 23446 59016
rect 4672 58908 6914 58936
rect 4672 58896 4678 58908
rect 20806 58896 20812 58948
rect 20864 58936 20870 58948
rect 23109 58939 23167 58945
rect 23109 58936 23121 58939
rect 20864 58908 23121 58936
rect 20864 58896 20870 58908
rect 23109 58905 23121 58908
rect 23155 58905 23167 58939
rect 23109 58899 23167 58905
rect 23658 58896 23664 58948
rect 23716 58896 23722 58948
rect 25682 58896 25688 58948
rect 25740 58936 25746 58948
rect 26206 58936 26234 59044
rect 30929 59041 30941 59044
rect 30975 59072 30987 59075
rect 31018 59072 31024 59084
rect 30975 59044 31024 59072
rect 30975 59041 30987 59044
rect 30929 59035 30987 59041
rect 31018 59032 31024 59044
rect 31076 59032 31082 59084
rect 38010 59032 38016 59084
rect 38068 59072 38074 59084
rect 38105 59075 38163 59081
rect 38105 59072 38117 59075
rect 38068 59044 38117 59072
rect 38068 59032 38074 59044
rect 38105 59041 38117 59044
rect 38151 59041 38163 59075
rect 38105 59035 38163 59041
rect 29914 58964 29920 59016
rect 29972 58964 29978 59016
rect 30469 59007 30527 59013
rect 30469 58973 30481 59007
rect 30515 58973 30527 59007
rect 30469 58967 30527 58973
rect 25740 58908 26234 58936
rect 25740 58896 25746 58908
rect 27430 58896 27436 58948
rect 27488 58936 27494 58948
rect 30484 58936 30512 58967
rect 31478 58964 31484 59016
rect 31536 59004 31542 59016
rect 38197 59007 38255 59013
rect 38197 59004 38209 59007
rect 31536 58976 38209 59004
rect 31536 58964 31542 58976
rect 38197 58973 38209 58976
rect 38243 58973 38255 59007
rect 38197 58967 38255 58973
rect 38381 59007 38439 59013
rect 38381 58973 38393 59007
rect 38427 58973 38439 59007
rect 38381 58967 38439 58973
rect 27488 58908 30512 58936
rect 27488 58896 27494 58908
rect 35158 58896 35164 58948
rect 35216 58936 35222 58948
rect 38396 58936 38424 58967
rect 35216 58908 38424 58936
rect 35216 58896 35222 58908
rect 30006 58828 30012 58880
rect 30064 58828 30070 58880
rect 1104 58778 40848 58800
rect 1104 58726 2610 58778
rect 2662 58726 2674 58778
rect 2726 58726 2738 58778
rect 2790 58726 2802 58778
rect 2854 58726 2866 58778
rect 2918 58726 7610 58778
rect 7662 58726 7674 58778
rect 7726 58726 7738 58778
rect 7790 58726 7802 58778
rect 7854 58726 7866 58778
rect 7918 58726 12610 58778
rect 12662 58726 12674 58778
rect 12726 58726 12738 58778
rect 12790 58726 12802 58778
rect 12854 58726 12866 58778
rect 12918 58726 17610 58778
rect 17662 58726 17674 58778
rect 17726 58726 17738 58778
rect 17790 58726 17802 58778
rect 17854 58726 17866 58778
rect 17918 58726 22610 58778
rect 22662 58726 22674 58778
rect 22726 58726 22738 58778
rect 22790 58726 22802 58778
rect 22854 58726 22866 58778
rect 22918 58726 27610 58778
rect 27662 58726 27674 58778
rect 27726 58726 27738 58778
rect 27790 58726 27802 58778
rect 27854 58726 27866 58778
rect 27918 58726 32610 58778
rect 32662 58726 32674 58778
rect 32726 58726 32738 58778
rect 32790 58726 32802 58778
rect 32854 58726 32866 58778
rect 32918 58726 37610 58778
rect 37662 58726 37674 58778
rect 37726 58726 37738 58778
rect 37790 58726 37802 58778
rect 37854 58726 37866 58778
rect 37918 58726 40848 58778
rect 1104 58704 40848 58726
rect 19242 58624 19248 58676
rect 19300 58664 19306 58676
rect 30098 58664 30104 58676
rect 19300 58636 30104 58664
rect 19300 58624 19306 58636
rect 30098 58624 30104 58636
rect 30156 58624 30162 58676
rect 2593 58599 2651 58605
rect 2593 58565 2605 58599
rect 2639 58596 2651 58599
rect 6730 58596 6736 58608
rect 2639 58568 6736 58596
rect 2639 58565 2651 58568
rect 2593 58559 2651 58565
rect 6730 58556 6736 58568
rect 6788 58556 6794 58608
rect 39298 58556 39304 58608
rect 39356 58556 39362 58608
rect 842 58488 848 58540
rect 900 58528 906 58540
rect 1397 58531 1455 58537
rect 1397 58528 1409 58531
rect 900 58500 1409 58528
rect 900 58488 906 58500
rect 1397 58497 1409 58500
rect 1443 58497 1455 58531
rect 1397 58491 1455 58497
rect 13909 58531 13967 58537
rect 13909 58497 13921 58531
rect 13955 58497 13967 58531
rect 13909 58491 13967 58497
rect 13924 58392 13952 58491
rect 14366 58488 14372 58540
rect 14424 58488 14430 58540
rect 14737 58531 14795 58537
rect 14737 58497 14749 58531
rect 14783 58528 14795 58531
rect 19886 58528 19892 58540
rect 14783 58500 19892 58528
rect 14783 58497 14795 58500
rect 14737 58491 14795 58497
rect 19886 58488 19892 58500
rect 19944 58488 19950 58540
rect 38657 58531 38715 58537
rect 38657 58528 38669 58531
rect 38212 58500 38669 58528
rect 13998 58420 14004 58472
rect 14056 58420 14062 58472
rect 38010 58420 38016 58472
rect 38068 58460 38074 58472
rect 38212 58460 38240 58500
rect 38657 58497 38669 58500
rect 38703 58497 38715 58531
rect 38657 58491 38715 58497
rect 39114 58488 39120 58540
rect 39172 58528 39178 58540
rect 39209 58531 39267 58537
rect 39209 58528 39221 58531
rect 39172 58500 39221 58528
rect 39172 58488 39178 58500
rect 39209 58497 39221 58500
rect 39255 58497 39267 58531
rect 39209 58491 39267 58497
rect 38068 58432 38240 58460
rect 38068 58420 38074 58432
rect 14182 58392 14188 58404
rect 13924 58364 14188 58392
rect 14182 58352 14188 58364
rect 14240 58352 14246 58404
rect 1104 58234 40848 58256
rect 1104 58182 1950 58234
rect 2002 58182 2014 58234
rect 2066 58182 2078 58234
rect 2130 58182 2142 58234
rect 2194 58182 2206 58234
rect 2258 58182 6950 58234
rect 7002 58182 7014 58234
rect 7066 58182 7078 58234
rect 7130 58182 7142 58234
rect 7194 58182 7206 58234
rect 7258 58182 11950 58234
rect 12002 58182 12014 58234
rect 12066 58182 12078 58234
rect 12130 58182 12142 58234
rect 12194 58182 12206 58234
rect 12258 58182 16950 58234
rect 17002 58182 17014 58234
rect 17066 58182 17078 58234
rect 17130 58182 17142 58234
rect 17194 58182 17206 58234
rect 17258 58182 21950 58234
rect 22002 58182 22014 58234
rect 22066 58182 22078 58234
rect 22130 58182 22142 58234
rect 22194 58182 22206 58234
rect 22258 58182 26950 58234
rect 27002 58182 27014 58234
rect 27066 58182 27078 58234
rect 27130 58182 27142 58234
rect 27194 58182 27206 58234
rect 27258 58182 31950 58234
rect 32002 58182 32014 58234
rect 32066 58182 32078 58234
rect 32130 58182 32142 58234
rect 32194 58182 32206 58234
rect 32258 58182 36950 58234
rect 37002 58182 37014 58234
rect 37066 58182 37078 58234
rect 37130 58182 37142 58234
rect 37194 58182 37206 58234
rect 37258 58182 40848 58234
rect 1104 58160 40848 58182
rect 26881 58123 26939 58129
rect 26881 58089 26893 58123
rect 26927 58120 26939 58123
rect 27522 58120 27528 58132
rect 26927 58092 27528 58120
rect 26927 58089 26939 58092
rect 26881 58083 26939 58089
rect 27522 58080 27528 58092
rect 27580 58080 27586 58132
rect 19886 57944 19892 57996
rect 19944 57944 19950 57996
rect 10962 57876 10968 57928
rect 11020 57916 11026 57928
rect 11020 57888 20024 57916
rect 11020 57876 11026 57888
rect 19996 57848 20024 57888
rect 20070 57876 20076 57928
rect 20128 57876 20134 57928
rect 20625 57919 20683 57925
rect 20625 57885 20637 57919
rect 20671 57916 20683 57919
rect 20714 57916 20720 57928
rect 20671 57888 20720 57916
rect 20671 57885 20683 57888
rect 20625 57879 20683 57885
rect 20714 57876 20720 57888
rect 20772 57876 20778 57928
rect 20990 57876 20996 57928
rect 21048 57876 21054 57928
rect 24673 57919 24731 57925
rect 24673 57885 24685 57919
rect 24719 57916 24731 57919
rect 27801 57919 27859 57925
rect 24719 57888 27752 57916
rect 24719 57885 24731 57888
rect 24673 57879 24731 57885
rect 27157 57851 27215 57857
rect 27157 57848 27169 57851
rect 19996 57820 27169 57848
rect 27157 57817 27169 57820
rect 27203 57817 27215 57851
rect 27724 57848 27752 57888
rect 27801 57885 27813 57919
rect 27847 57916 27859 57919
rect 28074 57916 28080 57928
rect 27847 57888 28080 57916
rect 27847 57885 27859 57888
rect 27801 57879 27859 57885
rect 28074 57876 28080 57888
rect 28132 57876 28138 57928
rect 28902 57848 28908 57860
rect 27724 57820 28908 57848
rect 27157 57811 27215 57817
rect 28902 57808 28908 57820
rect 28960 57808 28966 57860
rect 12434 57740 12440 57792
rect 12492 57780 12498 57792
rect 24489 57783 24547 57789
rect 24489 57780 24501 57783
rect 12492 57752 24501 57780
rect 12492 57740 12498 57752
rect 24489 57749 24501 57752
rect 24535 57749 24547 57783
rect 24489 57743 24547 57749
rect 26142 57740 26148 57792
rect 26200 57780 26206 57792
rect 27522 57780 27528 57792
rect 27580 57789 27586 57792
rect 26200 57752 27528 57780
rect 26200 57740 26206 57752
rect 27522 57740 27528 57752
rect 27580 57780 27592 57789
rect 27580 57752 27625 57780
rect 27580 57743 27592 57752
rect 27580 57740 27586 57743
rect 1104 57690 40848 57712
rect 1104 57638 2610 57690
rect 2662 57638 2674 57690
rect 2726 57638 2738 57690
rect 2790 57638 2802 57690
rect 2854 57638 2866 57690
rect 2918 57638 7610 57690
rect 7662 57638 7674 57690
rect 7726 57638 7738 57690
rect 7790 57638 7802 57690
rect 7854 57638 7866 57690
rect 7918 57638 12610 57690
rect 12662 57638 12674 57690
rect 12726 57638 12738 57690
rect 12790 57638 12802 57690
rect 12854 57638 12866 57690
rect 12918 57638 17610 57690
rect 17662 57638 17674 57690
rect 17726 57638 17738 57690
rect 17790 57638 17802 57690
rect 17854 57638 17866 57690
rect 17918 57638 22610 57690
rect 22662 57638 22674 57690
rect 22726 57638 22738 57690
rect 22790 57638 22802 57690
rect 22854 57638 22866 57690
rect 22918 57638 27610 57690
rect 27662 57638 27674 57690
rect 27726 57638 27738 57690
rect 27790 57638 27802 57690
rect 27854 57638 27866 57690
rect 27918 57638 32610 57690
rect 32662 57638 32674 57690
rect 32726 57638 32738 57690
rect 32790 57638 32802 57690
rect 32854 57638 32866 57690
rect 32918 57638 37610 57690
rect 37662 57638 37674 57690
rect 37726 57638 37738 57690
rect 37790 57638 37802 57690
rect 37854 57638 37866 57690
rect 37918 57638 40848 57690
rect 1104 57616 40848 57638
rect 20714 57536 20720 57588
rect 20772 57576 20778 57588
rect 24854 57576 24860 57588
rect 20772 57548 24860 57576
rect 20772 57536 20778 57548
rect 24854 57536 24860 57548
rect 24912 57536 24918 57588
rect 31662 57536 31668 57588
rect 31720 57576 31726 57588
rect 33410 57576 33416 57588
rect 31720 57548 33416 57576
rect 31720 57536 31726 57548
rect 33410 57536 33416 57548
rect 33468 57536 33474 57588
rect 16850 57400 16856 57452
rect 16908 57440 16914 57452
rect 17129 57443 17187 57449
rect 17129 57440 17141 57443
rect 16908 57412 17141 57440
rect 16908 57400 16914 57412
rect 17129 57409 17141 57412
rect 17175 57409 17187 57443
rect 17129 57403 17187 57409
rect 21542 57400 21548 57452
rect 21600 57440 21606 57452
rect 21600 57412 26234 57440
rect 21600 57400 21606 57412
rect 16666 57332 16672 57384
rect 16724 57332 16730 57384
rect 17221 57375 17279 57381
rect 17221 57341 17233 57375
rect 17267 57372 17279 57375
rect 22370 57372 22376 57384
rect 17267 57344 22376 57372
rect 17267 57341 17279 57344
rect 17221 57335 17279 57341
rect 22370 57332 22376 57344
rect 22428 57332 22434 57384
rect 26206 57372 26234 57412
rect 38930 57400 38936 57452
rect 38988 57440 38994 57452
rect 39025 57443 39083 57449
rect 39025 57440 39037 57443
rect 38988 57412 39037 57440
rect 38988 57400 38994 57412
rect 39025 57409 39037 57412
rect 39071 57409 39083 57443
rect 39025 57403 39083 57409
rect 39206 57400 39212 57452
rect 39264 57440 39270 57452
rect 39574 57440 39580 57452
rect 39264 57412 39580 57440
rect 39264 57400 39270 57412
rect 39574 57400 39580 57412
rect 39632 57400 39638 57452
rect 39850 57400 39856 57452
rect 39908 57400 39914 57452
rect 40221 57443 40279 57449
rect 40221 57409 40233 57443
rect 40267 57409 40279 57443
rect 40221 57403 40279 57409
rect 40236 57372 40264 57403
rect 26206 57344 40264 57372
rect 16114 57264 16120 57316
rect 16172 57304 16178 57316
rect 22278 57304 22284 57316
rect 16172 57276 22284 57304
rect 16172 57264 16178 57276
rect 22278 57264 22284 57276
rect 22336 57264 22342 57316
rect 23658 57264 23664 57316
rect 23716 57304 23722 57316
rect 31202 57304 31208 57316
rect 23716 57276 31208 57304
rect 23716 57264 23722 57276
rect 31202 57264 31208 57276
rect 31260 57264 31266 57316
rect 31294 57264 31300 57316
rect 31352 57304 31358 57316
rect 39117 57307 39175 57313
rect 39117 57304 39129 57307
rect 31352 57276 39129 57304
rect 31352 57264 31358 57276
rect 39117 57273 39129 57276
rect 39163 57273 39175 57307
rect 39117 57267 39175 57273
rect 2314 57196 2320 57248
rect 2372 57236 2378 57248
rect 33502 57236 33508 57248
rect 2372 57208 33508 57236
rect 2372 57196 2378 57208
rect 33502 57196 33508 57208
rect 33560 57196 33566 57248
rect 1104 57146 40848 57168
rect 1104 57094 1950 57146
rect 2002 57094 2014 57146
rect 2066 57094 2078 57146
rect 2130 57094 2142 57146
rect 2194 57094 2206 57146
rect 2258 57094 6950 57146
rect 7002 57094 7014 57146
rect 7066 57094 7078 57146
rect 7130 57094 7142 57146
rect 7194 57094 7206 57146
rect 7258 57094 11950 57146
rect 12002 57094 12014 57146
rect 12066 57094 12078 57146
rect 12130 57094 12142 57146
rect 12194 57094 12206 57146
rect 12258 57094 16950 57146
rect 17002 57094 17014 57146
rect 17066 57094 17078 57146
rect 17130 57094 17142 57146
rect 17194 57094 17206 57146
rect 17258 57094 21950 57146
rect 22002 57094 22014 57146
rect 22066 57094 22078 57146
rect 22130 57094 22142 57146
rect 22194 57094 22206 57146
rect 22258 57094 26950 57146
rect 27002 57094 27014 57146
rect 27066 57094 27078 57146
rect 27130 57094 27142 57146
rect 27194 57094 27206 57146
rect 27258 57094 31950 57146
rect 32002 57094 32014 57146
rect 32066 57094 32078 57146
rect 32130 57094 32142 57146
rect 32194 57094 32206 57146
rect 32258 57094 36950 57146
rect 37002 57094 37014 57146
rect 37066 57094 37078 57146
rect 37130 57094 37142 57146
rect 37194 57094 37206 57146
rect 37258 57094 40848 57146
rect 1104 57072 40848 57094
rect 26234 56992 26240 57044
rect 26292 57032 26298 57044
rect 35158 57032 35164 57044
rect 26292 57004 35164 57032
rect 26292 56992 26298 57004
rect 35158 56992 35164 57004
rect 35216 56992 35222 57044
rect 9030 56924 9036 56976
rect 9088 56964 9094 56976
rect 39850 56964 39856 56976
rect 9088 56936 39856 56964
rect 9088 56924 9094 56936
rect 39850 56924 39856 56936
rect 39908 56924 39914 56976
rect 10134 56856 10140 56908
rect 10192 56856 10198 56908
rect 10686 56856 10692 56908
rect 10744 56896 10750 56908
rect 19794 56896 19800 56908
rect 10744 56868 19800 56896
rect 10744 56856 10750 56868
rect 5074 56788 5080 56840
rect 5132 56828 5138 56840
rect 10045 56831 10103 56837
rect 10045 56828 10057 56831
rect 5132 56800 10057 56828
rect 5132 56788 5138 56800
rect 10045 56797 10057 56800
rect 10091 56797 10103 56831
rect 10045 56791 10103 56797
rect 10778 56788 10784 56840
rect 10836 56788 10842 56840
rect 10888 56837 10916 56868
rect 19794 56856 19800 56868
rect 19852 56856 19858 56908
rect 26421 56899 26479 56905
rect 26421 56865 26433 56899
rect 26467 56896 26479 56899
rect 31110 56896 31116 56908
rect 26467 56868 31116 56896
rect 26467 56865 26479 56868
rect 26421 56859 26479 56865
rect 31110 56856 31116 56868
rect 31168 56856 31174 56908
rect 10873 56831 10931 56837
rect 10873 56797 10885 56831
rect 10919 56797 10931 56831
rect 10873 56791 10931 56797
rect 11517 56831 11575 56837
rect 11517 56797 11529 56831
rect 11563 56828 11575 56831
rect 16298 56828 16304 56840
rect 11563 56800 16304 56828
rect 11563 56797 11575 56800
rect 11517 56791 11575 56797
rect 16298 56788 16304 56800
rect 16356 56788 16362 56840
rect 26142 56788 26148 56840
rect 26200 56828 26206 56840
rect 26234 56828 26240 56840
rect 26200 56800 26240 56828
rect 26200 56788 26206 56800
rect 26234 56788 26240 56800
rect 26292 56828 26298 56840
rect 26329 56831 26387 56837
rect 26329 56828 26341 56831
rect 26292 56800 26341 56828
rect 26292 56788 26298 56800
rect 26329 56797 26341 56800
rect 26375 56797 26387 56831
rect 26329 56791 26387 56797
rect 26789 56831 26847 56837
rect 26789 56797 26801 56831
rect 26835 56797 26847 56831
rect 26789 56791 26847 56797
rect 19978 56652 19984 56704
rect 20036 56692 20042 56704
rect 26804 56692 26832 56791
rect 20036 56664 26832 56692
rect 20036 56652 20042 56664
rect 1104 56602 40848 56624
rect 1104 56550 2610 56602
rect 2662 56550 2674 56602
rect 2726 56550 2738 56602
rect 2790 56550 2802 56602
rect 2854 56550 2866 56602
rect 2918 56550 7610 56602
rect 7662 56550 7674 56602
rect 7726 56550 7738 56602
rect 7790 56550 7802 56602
rect 7854 56550 7866 56602
rect 7918 56550 12610 56602
rect 12662 56550 12674 56602
rect 12726 56550 12738 56602
rect 12790 56550 12802 56602
rect 12854 56550 12866 56602
rect 12918 56550 17610 56602
rect 17662 56550 17674 56602
rect 17726 56550 17738 56602
rect 17790 56550 17802 56602
rect 17854 56550 17866 56602
rect 17918 56550 22610 56602
rect 22662 56550 22674 56602
rect 22726 56550 22738 56602
rect 22790 56550 22802 56602
rect 22854 56550 22866 56602
rect 22918 56550 27610 56602
rect 27662 56550 27674 56602
rect 27726 56550 27738 56602
rect 27790 56550 27802 56602
rect 27854 56550 27866 56602
rect 27918 56550 32610 56602
rect 32662 56550 32674 56602
rect 32726 56550 32738 56602
rect 32790 56550 32802 56602
rect 32854 56550 32866 56602
rect 32918 56550 37610 56602
rect 37662 56550 37674 56602
rect 37726 56550 37738 56602
rect 37790 56550 37802 56602
rect 37854 56550 37866 56602
rect 37918 56550 40848 56602
rect 1104 56528 40848 56550
rect 24210 56176 24216 56228
rect 24268 56216 24274 56228
rect 29086 56216 29092 56228
rect 24268 56188 29092 56216
rect 24268 56176 24274 56188
rect 29086 56176 29092 56188
rect 29144 56176 29150 56228
rect 13814 56108 13820 56160
rect 13872 56148 13878 56160
rect 33962 56148 33968 56160
rect 13872 56120 33968 56148
rect 13872 56108 13878 56120
rect 33962 56108 33968 56120
rect 34020 56108 34026 56160
rect 1104 56058 40848 56080
rect 1104 56006 1950 56058
rect 2002 56006 2014 56058
rect 2066 56006 2078 56058
rect 2130 56006 2142 56058
rect 2194 56006 2206 56058
rect 2258 56006 6950 56058
rect 7002 56006 7014 56058
rect 7066 56006 7078 56058
rect 7130 56006 7142 56058
rect 7194 56006 7206 56058
rect 7258 56006 11950 56058
rect 12002 56006 12014 56058
rect 12066 56006 12078 56058
rect 12130 56006 12142 56058
rect 12194 56006 12206 56058
rect 12258 56006 16950 56058
rect 17002 56006 17014 56058
rect 17066 56006 17078 56058
rect 17130 56006 17142 56058
rect 17194 56006 17206 56058
rect 17258 56006 21950 56058
rect 22002 56006 22014 56058
rect 22066 56006 22078 56058
rect 22130 56006 22142 56058
rect 22194 56006 22206 56058
rect 22258 56006 26950 56058
rect 27002 56006 27014 56058
rect 27066 56006 27078 56058
rect 27130 56006 27142 56058
rect 27194 56006 27206 56058
rect 27258 56006 31950 56058
rect 32002 56006 32014 56058
rect 32066 56006 32078 56058
rect 32130 56006 32142 56058
rect 32194 56006 32206 56058
rect 32258 56006 36950 56058
rect 37002 56006 37014 56058
rect 37066 56006 37078 56058
rect 37130 56006 37142 56058
rect 37194 56006 37206 56058
rect 37258 56006 40848 56058
rect 1104 55984 40848 56006
rect 10686 55904 10692 55956
rect 10744 55944 10750 55956
rect 39298 55944 39304 55956
rect 10744 55916 39304 55944
rect 10744 55904 10750 55916
rect 39298 55904 39304 55916
rect 39356 55904 39362 55956
rect 3786 55836 3792 55888
rect 3844 55876 3850 55888
rect 10962 55876 10968 55888
rect 3844 55848 10968 55876
rect 3844 55836 3850 55848
rect 10962 55836 10968 55848
rect 11020 55836 11026 55888
rect 15930 55836 15936 55888
rect 15988 55836 15994 55888
rect 19426 55836 19432 55888
rect 19484 55876 19490 55888
rect 34698 55876 34704 55888
rect 19484 55848 34704 55876
rect 19484 55836 19490 55848
rect 34698 55836 34704 55848
rect 34756 55836 34762 55888
rect 9398 55768 9404 55820
rect 9456 55808 9462 55820
rect 9585 55811 9643 55817
rect 9585 55808 9597 55811
rect 9456 55780 9597 55808
rect 9456 55768 9462 55780
rect 9585 55777 9597 55780
rect 9631 55777 9643 55811
rect 9585 55771 9643 55777
rect 22370 55768 22376 55820
rect 22428 55808 22434 55820
rect 23198 55808 23204 55820
rect 22428 55780 23204 55808
rect 22428 55768 22434 55780
rect 23198 55768 23204 55780
rect 23256 55768 23262 55820
rect 9490 55700 9496 55752
rect 9548 55700 9554 55752
rect 9950 55700 9956 55752
rect 10008 55700 10014 55752
rect 11698 55700 11704 55752
rect 11756 55740 11762 55752
rect 15841 55743 15899 55749
rect 15841 55740 15853 55743
rect 11756 55712 15853 55740
rect 11756 55700 11762 55712
rect 15841 55709 15853 55712
rect 15887 55709 15899 55743
rect 15841 55703 15899 55709
rect 16363 55743 16421 55749
rect 16363 55709 16375 55743
rect 16409 55740 16421 55743
rect 17954 55740 17960 55752
rect 16409 55712 17960 55740
rect 16409 55709 16421 55712
rect 16363 55703 16421 55709
rect 17954 55700 17960 55712
rect 18012 55740 18018 55752
rect 19242 55740 19248 55752
rect 18012 55712 19248 55740
rect 18012 55700 18018 55712
rect 19242 55700 19248 55712
rect 19300 55700 19306 55752
rect 10137 55675 10195 55681
rect 10137 55641 10149 55675
rect 10183 55672 10195 55675
rect 24118 55672 24124 55684
rect 10183 55644 24124 55672
rect 10183 55641 10195 55644
rect 10137 55635 10195 55641
rect 24118 55632 24124 55644
rect 24176 55632 24182 55684
rect 16298 55564 16304 55616
rect 16356 55564 16362 55616
rect 16482 55564 16488 55616
rect 16540 55564 16546 55616
rect 1104 55514 40848 55536
rect 1104 55462 2610 55514
rect 2662 55462 2674 55514
rect 2726 55462 2738 55514
rect 2790 55462 2802 55514
rect 2854 55462 2866 55514
rect 2918 55462 7610 55514
rect 7662 55462 7674 55514
rect 7726 55462 7738 55514
rect 7790 55462 7802 55514
rect 7854 55462 7866 55514
rect 7918 55462 12610 55514
rect 12662 55462 12674 55514
rect 12726 55462 12738 55514
rect 12790 55462 12802 55514
rect 12854 55462 12866 55514
rect 12918 55462 17610 55514
rect 17662 55462 17674 55514
rect 17726 55462 17738 55514
rect 17790 55462 17802 55514
rect 17854 55462 17866 55514
rect 17918 55462 22610 55514
rect 22662 55462 22674 55514
rect 22726 55462 22738 55514
rect 22790 55462 22802 55514
rect 22854 55462 22866 55514
rect 22918 55462 27610 55514
rect 27662 55462 27674 55514
rect 27726 55462 27738 55514
rect 27790 55462 27802 55514
rect 27854 55462 27866 55514
rect 27918 55462 32610 55514
rect 32662 55462 32674 55514
rect 32726 55462 32738 55514
rect 32790 55462 32802 55514
rect 32854 55462 32866 55514
rect 32918 55462 37610 55514
rect 37662 55462 37674 55514
rect 37726 55462 37738 55514
rect 37790 55462 37802 55514
rect 37854 55462 37866 55514
rect 37918 55462 40848 55514
rect 1104 55440 40848 55462
rect 13722 55332 13728 55344
rect 4908 55304 13728 55332
rect 4908 55273 4936 55304
rect 13722 55292 13728 55304
rect 13780 55332 13786 55344
rect 14458 55332 14464 55344
rect 13780 55304 14464 55332
rect 13780 55292 13786 55304
rect 14458 55292 14464 55304
rect 14516 55292 14522 55344
rect 4893 55267 4951 55273
rect 4893 55233 4905 55267
rect 4939 55233 4951 55267
rect 4893 55227 4951 55233
rect 5261 55267 5319 55273
rect 5261 55233 5273 55267
rect 5307 55264 5319 55267
rect 6178 55264 6184 55276
rect 5307 55236 6184 55264
rect 5307 55233 5319 55236
rect 5261 55227 5319 55233
rect 6178 55224 6184 55236
rect 6236 55224 6242 55276
rect 13446 55156 13452 55208
rect 13504 55196 13510 55208
rect 14642 55196 14648 55208
rect 13504 55168 14648 55196
rect 13504 55156 13510 55168
rect 14642 55156 14648 55168
rect 14700 55156 14706 55208
rect 5813 55063 5871 55069
rect 5813 55029 5825 55063
rect 5859 55060 5871 55063
rect 6270 55060 6276 55072
rect 5859 55032 6276 55060
rect 5859 55029 5871 55032
rect 5813 55023 5871 55029
rect 6270 55020 6276 55032
rect 6328 55020 6334 55072
rect 1104 54970 40848 54992
rect 1104 54918 1950 54970
rect 2002 54918 2014 54970
rect 2066 54918 2078 54970
rect 2130 54918 2142 54970
rect 2194 54918 2206 54970
rect 2258 54918 6950 54970
rect 7002 54918 7014 54970
rect 7066 54918 7078 54970
rect 7130 54918 7142 54970
rect 7194 54918 7206 54970
rect 7258 54918 11950 54970
rect 12002 54918 12014 54970
rect 12066 54918 12078 54970
rect 12130 54918 12142 54970
rect 12194 54918 12206 54970
rect 12258 54918 16950 54970
rect 17002 54918 17014 54970
rect 17066 54918 17078 54970
rect 17130 54918 17142 54970
rect 17194 54918 17206 54970
rect 17258 54918 21950 54970
rect 22002 54918 22014 54970
rect 22066 54918 22078 54970
rect 22130 54918 22142 54970
rect 22194 54918 22206 54970
rect 22258 54918 26950 54970
rect 27002 54918 27014 54970
rect 27066 54918 27078 54970
rect 27130 54918 27142 54970
rect 27194 54918 27206 54970
rect 27258 54918 31950 54970
rect 32002 54918 32014 54970
rect 32066 54918 32078 54970
rect 32130 54918 32142 54970
rect 32194 54918 32206 54970
rect 32258 54918 36950 54970
rect 37002 54918 37014 54970
rect 37066 54918 37078 54970
rect 37130 54918 37142 54970
rect 37194 54918 37206 54970
rect 37258 54918 40848 54970
rect 1104 54896 40848 54918
rect 35066 54788 35072 54800
rect 26206 54760 35072 54788
rect 6730 54680 6736 54732
rect 6788 54720 6794 54732
rect 7466 54720 7472 54732
rect 6788 54692 7472 54720
rect 6788 54680 6794 54692
rect 7466 54680 7472 54692
rect 7524 54720 7530 54732
rect 15470 54720 15476 54732
rect 7524 54692 15476 54720
rect 7524 54680 7530 54692
rect 15470 54680 15476 54692
rect 15528 54680 15534 54732
rect 24854 54680 24860 54732
rect 24912 54720 24918 54732
rect 26206 54720 26234 54760
rect 35066 54748 35072 54760
rect 35124 54748 35130 54800
rect 34882 54720 34888 54732
rect 24912 54692 26234 54720
rect 29840 54692 34888 54720
rect 24912 54680 24918 54692
rect 6825 54655 6883 54661
rect 6825 54621 6837 54655
rect 6871 54652 6883 54655
rect 8202 54652 8208 54664
rect 6871 54624 8208 54652
rect 6871 54621 6883 54624
rect 6825 54615 6883 54621
rect 8202 54612 8208 54624
rect 8260 54612 8266 54664
rect 15749 54655 15807 54661
rect 15749 54621 15761 54655
rect 15795 54652 15807 54655
rect 29840 54652 29868 54692
rect 34882 54680 34888 54692
rect 34940 54680 34946 54732
rect 15795 54624 29868 54652
rect 15795 54621 15807 54624
rect 15749 54615 15807 54621
rect 29914 54612 29920 54664
rect 29972 54652 29978 54664
rect 33873 54655 33931 54661
rect 33873 54652 33885 54655
rect 29972 54624 33885 54652
rect 29972 54612 29978 54624
rect 33873 54621 33885 54624
rect 33919 54621 33931 54655
rect 33873 54615 33931 54621
rect 5534 54544 5540 54596
rect 5592 54584 5598 54596
rect 5902 54584 5908 54596
rect 5592 54556 5908 54584
rect 5592 54544 5598 54556
rect 5902 54544 5908 54556
rect 5960 54544 5966 54596
rect 6546 54544 6552 54596
rect 6604 54544 6610 54596
rect 6917 54587 6975 54593
rect 6917 54553 6929 54587
rect 6963 54584 6975 54587
rect 9306 54584 9312 54596
rect 6963 54556 9312 54584
rect 6963 54553 6975 54556
rect 6917 54547 6975 54553
rect 9306 54544 9312 54556
rect 9364 54544 9370 54596
rect 14366 54544 14372 54596
rect 14424 54584 14430 54596
rect 30282 54584 30288 54596
rect 14424 54556 30288 54584
rect 14424 54544 14430 54556
rect 30282 54544 30288 54556
rect 30340 54544 30346 54596
rect 4246 54476 4252 54528
rect 4304 54516 4310 54528
rect 4706 54516 4712 54528
rect 4304 54488 4712 54516
rect 4304 54476 4310 54488
rect 4706 54476 4712 54488
rect 4764 54476 4770 54528
rect 6730 54476 6736 54528
rect 6788 54476 6794 54528
rect 7098 54476 7104 54528
rect 7156 54476 7162 54528
rect 33962 54476 33968 54528
rect 34020 54476 34026 54528
rect 1104 54426 40848 54448
rect 1104 54374 2610 54426
rect 2662 54374 2674 54426
rect 2726 54374 2738 54426
rect 2790 54374 2802 54426
rect 2854 54374 2866 54426
rect 2918 54374 7610 54426
rect 7662 54374 7674 54426
rect 7726 54374 7738 54426
rect 7790 54374 7802 54426
rect 7854 54374 7866 54426
rect 7918 54374 12610 54426
rect 12662 54374 12674 54426
rect 12726 54374 12738 54426
rect 12790 54374 12802 54426
rect 12854 54374 12866 54426
rect 12918 54374 17610 54426
rect 17662 54374 17674 54426
rect 17726 54374 17738 54426
rect 17790 54374 17802 54426
rect 17854 54374 17866 54426
rect 17918 54374 22610 54426
rect 22662 54374 22674 54426
rect 22726 54374 22738 54426
rect 22790 54374 22802 54426
rect 22854 54374 22866 54426
rect 22918 54374 27610 54426
rect 27662 54374 27674 54426
rect 27726 54374 27738 54426
rect 27790 54374 27802 54426
rect 27854 54374 27866 54426
rect 27918 54374 32610 54426
rect 32662 54374 32674 54426
rect 32726 54374 32738 54426
rect 32790 54374 32802 54426
rect 32854 54374 32866 54426
rect 32918 54374 37610 54426
rect 37662 54374 37674 54426
rect 37726 54374 37738 54426
rect 37790 54374 37802 54426
rect 37854 54374 37866 54426
rect 37918 54374 40848 54426
rect 1104 54352 40848 54374
rect 7098 54272 7104 54324
rect 7156 54312 7162 54324
rect 29914 54312 29920 54324
rect 7156 54284 29920 54312
rect 7156 54272 7162 54284
rect 29914 54272 29920 54284
rect 29972 54272 29978 54324
rect 15565 54247 15623 54253
rect 15565 54213 15577 54247
rect 15611 54244 15623 54247
rect 21542 54244 21548 54256
rect 15611 54216 21548 54244
rect 15611 54213 15623 54216
rect 15565 54207 15623 54213
rect 21542 54204 21548 54216
rect 21600 54204 21606 54256
rect 22066 54216 28672 54244
rect 15286 54136 15292 54188
rect 15344 54176 15350 54188
rect 15381 54179 15439 54185
rect 15381 54176 15393 54179
rect 15344 54148 15393 54176
rect 15344 54136 15350 54148
rect 15381 54145 15393 54148
rect 15427 54145 15439 54179
rect 15381 54139 15439 54145
rect 19150 54136 19156 54188
rect 19208 54176 19214 54188
rect 20346 54176 20352 54188
rect 19208 54148 20352 54176
rect 19208 54136 19214 54148
rect 20346 54136 20352 54148
rect 20404 54176 20410 54188
rect 22066 54176 22094 54216
rect 20404 54148 22094 54176
rect 20404 54136 20410 54148
rect 28074 54136 28080 54188
rect 28132 54176 28138 54188
rect 28258 54176 28264 54188
rect 28132 54148 28264 54176
rect 28132 54136 28138 54148
rect 28258 54136 28264 54148
rect 28316 54136 28322 54188
rect 28644 54185 28672 54216
rect 28629 54179 28687 54185
rect 28629 54145 28641 54179
rect 28675 54145 28687 54179
rect 28629 54139 28687 54145
rect 28994 54136 29000 54188
rect 29052 54136 29058 54188
rect 13170 54000 13176 54052
rect 13228 54040 13234 54052
rect 15930 54040 15936 54052
rect 13228 54012 15936 54040
rect 13228 54000 13234 54012
rect 15930 54000 15936 54012
rect 15988 54000 15994 54052
rect 6086 53932 6092 53984
rect 6144 53972 6150 53984
rect 6546 53972 6552 53984
rect 6144 53944 6552 53972
rect 6144 53932 6150 53944
rect 6546 53932 6552 53944
rect 6604 53932 6610 53984
rect 28350 53932 28356 53984
rect 28408 53932 28414 53984
rect 1104 53882 40848 53904
rect 1104 53830 1950 53882
rect 2002 53830 2014 53882
rect 2066 53830 2078 53882
rect 2130 53830 2142 53882
rect 2194 53830 2206 53882
rect 2258 53830 6950 53882
rect 7002 53830 7014 53882
rect 7066 53830 7078 53882
rect 7130 53830 7142 53882
rect 7194 53830 7206 53882
rect 7258 53830 11950 53882
rect 12002 53830 12014 53882
rect 12066 53830 12078 53882
rect 12130 53830 12142 53882
rect 12194 53830 12206 53882
rect 12258 53830 16950 53882
rect 17002 53830 17014 53882
rect 17066 53830 17078 53882
rect 17130 53830 17142 53882
rect 17194 53830 17206 53882
rect 17258 53830 21950 53882
rect 22002 53830 22014 53882
rect 22066 53830 22078 53882
rect 22130 53830 22142 53882
rect 22194 53830 22206 53882
rect 22258 53830 26950 53882
rect 27002 53830 27014 53882
rect 27066 53830 27078 53882
rect 27130 53830 27142 53882
rect 27194 53830 27206 53882
rect 27258 53830 31950 53882
rect 32002 53830 32014 53882
rect 32066 53830 32078 53882
rect 32130 53830 32142 53882
rect 32194 53830 32206 53882
rect 32258 53830 36950 53882
rect 37002 53830 37014 53882
rect 37066 53830 37078 53882
rect 37130 53830 37142 53882
rect 37194 53830 37206 53882
rect 37258 53830 40848 53882
rect 1104 53808 40848 53830
rect 14918 53660 14924 53712
rect 14976 53700 14982 53712
rect 15378 53700 15384 53712
rect 14976 53672 15384 53700
rect 14976 53660 14982 53672
rect 15378 53660 15384 53672
rect 15436 53660 15442 53712
rect 5994 53632 6000 53644
rect 4080 53604 6000 53632
rect 4080 53573 4108 53604
rect 5994 53592 6000 53604
rect 6052 53592 6058 53644
rect 9306 53592 9312 53644
rect 9364 53632 9370 53644
rect 9364 53604 22094 53632
rect 9364 53592 9370 53604
rect 4065 53567 4123 53573
rect 4065 53533 4077 53567
rect 4111 53533 4123 53567
rect 4065 53527 4123 53533
rect 4341 53567 4399 53573
rect 4341 53533 4353 53567
rect 4387 53564 4399 53567
rect 4430 53564 4436 53576
rect 4387 53536 4436 53564
rect 4387 53533 4399 53536
rect 4341 53527 4399 53533
rect 4430 53524 4436 53536
rect 4488 53524 4494 53576
rect 15120 53573 15148 53604
rect 15105 53567 15163 53573
rect 6886 53536 15056 53564
rect 4525 53499 4583 53505
rect 4525 53465 4537 53499
rect 4571 53465 4583 53499
rect 4525 53459 4583 53465
rect 4540 53428 4568 53459
rect 6886 53428 6914 53536
rect 8202 53456 8208 53508
rect 8260 53496 8266 53508
rect 14918 53496 14924 53508
rect 8260 53468 14924 53496
rect 8260 53456 8266 53468
rect 14918 53456 14924 53468
rect 14976 53456 14982 53508
rect 15028 53496 15056 53536
rect 15105 53533 15117 53567
rect 15151 53533 15163 53567
rect 15105 53527 15163 53533
rect 15378 53524 15384 53576
rect 15436 53524 15442 53576
rect 15028 53468 15424 53496
rect 4540 53400 6914 53428
rect 7282 53388 7288 53440
rect 7340 53428 7346 53440
rect 15286 53428 15292 53440
rect 7340 53400 15292 53428
rect 7340 53388 7346 53400
rect 15286 53388 15292 53400
rect 15344 53388 15350 53440
rect 15396 53428 15424 53468
rect 15470 53456 15476 53508
rect 15528 53456 15534 53508
rect 15838 53456 15844 53508
rect 15896 53456 15902 53508
rect 22066 53496 22094 53604
rect 38286 53524 38292 53576
rect 38344 53524 38350 53576
rect 26786 53496 26792 53508
rect 22066 53468 26792 53496
rect 26786 53456 26792 53468
rect 26844 53456 26850 53508
rect 39206 53456 39212 53508
rect 39264 53456 39270 53508
rect 23106 53428 23112 53440
rect 15396 53400 23112 53428
rect 23106 53388 23112 53400
rect 23164 53428 23170 53440
rect 28442 53428 28448 53440
rect 23164 53400 28448 53428
rect 23164 53388 23170 53400
rect 28442 53388 28448 53400
rect 28500 53388 28506 53440
rect 1104 53338 40848 53360
rect 1104 53286 2610 53338
rect 2662 53286 2674 53338
rect 2726 53286 2738 53338
rect 2790 53286 2802 53338
rect 2854 53286 2866 53338
rect 2918 53286 7610 53338
rect 7662 53286 7674 53338
rect 7726 53286 7738 53338
rect 7790 53286 7802 53338
rect 7854 53286 7866 53338
rect 7918 53286 12610 53338
rect 12662 53286 12674 53338
rect 12726 53286 12738 53338
rect 12790 53286 12802 53338
rect 12854 53286 12866 53338
rect 12918 53286 17610 53338
rect 17662 53286 17674 53338
rect 17726 53286 17738 53338
rect 17790 53286 17802 53338
rect 17854 53286 17866 53338
rect 17918 53286 22610 53338
rect 22662 53286 22674 53338
rect 22726 53286 22738 53338
rect 22790 53286 22802 53338
rect 22854 53286 22866 53338
rect 22918 53286 27610 53338
rect 27662 53286 27674 53338
rect 27726 53286 27738 53338
rect 27790 53286 27802 53338
rect 27854 53286 27866 53338
rect 27918 53286 32610 53338
rect 32662 53286 32674 53338
rect 32726 53286 32738 53338
rect 32790 53286 32802 53338
rect 32854 53286 32866 53338
rect 32918 53286 37610 53338
rect 37662 53286 37674 53338
rect 37726 53286 37738 53338
rect 37790 53286 37802 53338
rect 37854 53286 37866 53338
rect 37918 53286 40848 53338
rect 1104 53264 40848 53286
rect 2498 53116 2504 53168
rect 2556 53156 2562 53168
rect 21726 53156 21732 53168
rect 2556 53128 21732 53156
rect 2556 53116 2562 53128
rect 21726 53116 21732 53128
rect 21784 53116 21790 53168
rect 36446 53116 36452 53168
rect 36504 53156 36510 53168
rect 36722 53156 36728 53168
rect 36504 53128 36728 53156
rect 36504 53116 36510 53128
rect 36722 53116 36728 53128
rect 36780 53156 36786 53168
rect 37001 53159 37059 53165
rect 37001 53156 37013 53159
rect 36780 53128 37013 53156
rect 36780 53116 36786 53128
rect 37001 53125 37013 53128
rect 37047 53125 37059 53159
rect 37001 53119 37059 53125
rect 15286 53048 15292 53100
rect 15344 53048 15350 53100
rect 15562 53048 15568 53100
rect 15620 53088 15626 53100
rect 16206 53088 16212 53100
rect 15620 53060 16212 53088
rect 15620 53048 15626 53060
rect 16206 53048 16212 53060
rect 16264 53048 16270 53100
rect 33686 53048 33692 53100
rect 33744 53088 33750 53100
rect 34054 53088 34060 53100
rect 33744 53060 34060 53088
rect 33744 53048 33750 53060
rect 34054 53048 34060 53060
rect 34112 53088 34118 53100
rect 36817 53091 36875 53097
rect 36817 53088 36829 53091
rect 34112 53060 36829 53088
rect 34112 53048 34118 53060
rect 36817 53057 36829 53060
rect 36863 53057 36875 53091
rect 36817 53051 36875 53057
rect 15930 52980 15936 53032
rect 15988 52980 15994 53032
rect 15194 52912 15200 52964
rect 15252 52952 15258 52964
rect 15289 52955 15347 52961
rect 15289 52952 15301 52955
rect 15252 52924 15301 52952
rect 15252 52912 15258 52924
rect 15289 52921 15301 52924
rect 15335 52952 15347 52955
rect 38746 52952 38752 52964
rect 15335 52924 38752 52952
rect 15335 52921 15347 52924
rect 15289 52915 15347 52921
rect 38746 52912 38752 52924
rect 38804 52912 38810 52964
rect 36722 52844 36728 52896
rect 36780 52844 36786 52896
rect 1104 52794 40848 52816
rect 1104 52742 1950 52794
rect 2002 52742 2014 52794
rect 2066 52742 2078 52794
rect 2130 52742 2142 52794
rect 2194 52742 2206 52794
rect 2258 52742 6950 52794
rect 7002 52742 7014 52794
rect 7066 52742 7078 52794
rect 7130 52742 7142 52794
rect 7194 52742 7206 52794
rect 7258 52742 11950 52794
rect 12002 52742 12014 52794
rect 12066 52742 12078 52794
rect 12130 52742 12142 52794
rect 12194 52742 12206 52794
rect 12258 52742 16950 52794
rect 17002 52742 17014 52794
rect 17066 52742 17078 52794
rect 17130 52742 17142 52794
rect 17194 52742 17206 52794
rect 17258 52742 21950 52794
rect 22002 52742 22014 52794
rect 22066 52742 22078 52794
rect 22130 52742 22142 52794
rect 22194 52742 22206 52794
rect 22258 52742 26950 52794
rect 27002 52742 27014 52794
rect 27066 52742 27078 52794
rect 27130 52742 27142 52794
rect 27194 52742 27206 52794
rect 27258 52742 31950 52794
rect 32002 52742 32014 52794
rect 32066 52742 32078 52794
rect 32130 52742 32142 52794
rect 32194 52742 32206 52794
rect 32258 52742 36950 52794
rect 37002 52742 37014 52794
rect 37066 52742 37078 52794
rect 37130 52742 37142 52794
rect 37194 52742 37206 52794
rect 37258 52742 40848 52794
rect 1104 52720 40848 52742
rect 5994 52640 6000 52692
rect 6052 52680 6058 52692
rect 6546 52680 6552 52692
rect 6052 52652 6552 52680
rect 6052 52640 6058 52652
rect 6546 52640 6552 52652
rect 6604 52640 6610 52692
rect 36814 52640 36820 52692
rect 36872 52680 36878 52692
rect 39301 52683 39359 52689
rect 39301 52680 39313 52683
rect 36872 52652 39313 52680
rect 36872 52640 36878 52652
rect 39301 52649 39313 52652
rect 39347 52649 39359 52683
rect 39301 52643 39359 52649
rect 8202 52612 8208 52624
rect 5552 52584 8208 52612
rect 5552 52485 5580 52584
rect 8202 52572 8208 52584
rect 8260 52572 8266 52624
rect 20990 52612 20996 52624
rect 12406 52584 20996 52612
rect 7377 52547 7435 52553
rect 7377 52513 7389 52547
rect 7423 52544 7435 52547
rect 12406 52544 12434 52584
rect 20990 52572 20996 52584
rect 21048 52612 21054 52624
rect 23474 52612 23480 52624
rect 21048 52584 23480 52612
rect 21048 52572 21054 52584
rect 23474 52572 23480 52584
rect 23532 52572 23538 52624
rect 29454 52572 29460 52624
rect 29512 52612 29518 52624
rect 39117 52615 39175 52621
rect 39117 52612 39129 52615
rect 29512 52584 39129 52612
rect 29512 52572 29518 52584
rect 39117 52581 39129 52584
rect 39163 52581 39175 52615
rect 39117 52575 39175 52581
rect 7423 52516 12434 52544
rect 7423 52513 7435 52516
rect 7377 52507 7435 52513
rect 20530 52504 20536 52556
rect 20588 52544 20594 52556
rect 35253 52547 35311 52553
rect 35253 52544 35265 52547
rect 20588 52516 35265 52544
rect 20588 52504 20594 52516
rect 35253 52513 35265 52516
rect 35299 52513 35311 52547
rect 35253 52507 35311 52513
rect 5537 52479 5595 52485
rect 5537 52445 5549 52479
rect 5583 52445 5595 52479
rect 5537 52439 5595 52445
rect 6457 52479 6515 52485
rect 6457 52445 6469 52479
rect 6503 52476 6515 52479
rect 13906 52476 13912 52488
rect 6503 52448 13912 52476
rect 6503 52445 6515 52448
rect 6457 52439 6515 52445
rect 13906 52436 13912 52448
rect 13964 52436 13970 52488
rect 21726 52436 21732 52488
rect 21784 52476 21790 52488
rect 35069 52479 35127 52485
rect 35069 52476 35081 52479
rect 21784 52448 35081 52476
rect 21784 52436 21790 52448
rect 35069 52445 35081 52448
rect 35115 52476 35127 52479
rect 35529 52479 35587 52485
rect 35529 52476 35541 52479
rect 35115 52448 35541 52476
rect 35115 52445 35127 52448
rect 35069 52439 35127 52445
rect 35529 52445 35541 52448
rect 35575 52445 35587 52479
rect 35529 52439 35587 52445
rect 35802 52436 35808 52488
rect 35860 52436 35866 52488
rect 36538 52436 36544 52488
rect 36596 52436 36602 52488
rect 38194 52436 38200 52488
rect 38252 52476 38258 52488
rect 38841 52479 38899 52485
rect 38841 52476 38853 52479
rect 38252 52448 38853 52476
rect 38252 52436 38258 52448
rect 38841 52445 38853 52448
rect 38887 52445 38899 52479
rect 38841 52439 38899 52445
rect 34698 52368 34704 52420
rect 34756 52368 34762 52420
rect 34882 52300 34888 52352
rect 34940 52300 34946 52352
rect 34974 52300 34980 52352
rect 35032 52300 35038 52352
rect 1104 52250 40848 52272
rect 1104 52198 2610 52250
rect 2662 52198 2674 52250
rect 2726 52198 2738 52250
rect 2790 52198 2802 52250
rect 2854 52198 2866 52250
rect 2918 52198 7610 52250
rect 7662 52198 7674 52250
rect 7726 52198 7738 52250
rect 7790 52198 7802 52250
rect 7854 52198 7866 52250
rect 7918 52198 12610 52250
rect 12662 52198 12674 52250
rect 12726 52198 12738 52250
rect 12790 52198 12802 52250
rect 12854 52198 12866 52250
rect 12918 52198 17610 52250
rect 17662 52198 17674 52250
rect 17726 52198 17738 52250
rect 17790 52198 17802 52250
rect 17854 52198 17866 52250
rect 17918 52198 22610 52250
rect 22662 52198 22674 52250
rect 22726 52198 22738 52250
rect 22790 52198 22802 52250
rect 22854 52198 22866 52250
rect 22918 52198 27610 52250
rect 27662 52198 27674 52250
rect 27726 52198 27738 52250
rect 27790 52198 27802 52250
rect 27854 52198 27866 52250
rect 27918 52198 32610 52250
rect 32662 52198 32674 52250
rect 32726 52198 32738 52250
rect 32790 52198 32802 52250
rect 32854 52198 32866 52250
rect 32918 52198 37610 52250
rect 37662 52198 37674 52250
rect 37726 52198 37738 52250
rect 37790 52198 37802 52250
rect 37854 52198 37866 52250
rect 37918 52198 40848 52250
rect 1104 52176 40848 52198
rect 16850 52096 16856 52148
rect 16908 52136 16914 52148
rect 21634 52136 21640 52148
rect 16908 52108 21640 52136
rect 16908 52096 16914 52108
rect 21634 52096 21640 52108
rect 21692 52096 21698 52148
rect 35802 52096 35808 52148
rect 35860 52096 35866 52148
rect 10870 52028 10876 52080
rect 10928 52068 10934 52080
rect 20530 52068 20536 52080
rect 10928 52040 20536 52068
rect 10928 52028 10934 52040
rect 20530 52028 20536 52040
rect 20588 52028 20594 52080
rect 21361 52071 21419 52077
rect 21008 52040 21168 52068
rect 4709 52003 4767 52009
rect 4709 51969 4721 52003
rect 4755 51969 4767 52003
rect 4709 51963 4767 51969
rect 4724 51864 4752 51963
rect 4890 51960 4896 52012
rect 4948 51960 4954 52012
rect 5445 52003 5503 52009
rect 5445 51969 5457 52003
rect 5491 52000 5503 52003
rect 11238 52000 11244 52012
rect 5491 51972 11244 52000
rect 5491 51969 5503 51972
rect 5445 51963 5503 51969
rect 11238 51960 11244 51972
rect 11296 51960 11302 52012
rect 15378 51960 15384 52012
rect 15436 52000 15442 52012
rect 15436 51972 20760 52000
rect 15436 51960 15442 51972
rect 5353 51935 5411 51941
rect 5353 51901 5365 51935
rect 5399 51932 5411 51935
rect 18138 51932 18144 51944
rect 5399 51904 18144 51932
rect 5399 51901 5411 51904
rect 5353 51895 5411 51901
rect 18138 51892 18144 51904
rect 18196 51892 18202 51944
rect 20622 51892 20628 51944
rect 20680 51892 20686 51944
rect 20732 51932 20760 51972
rect 21008 51932 21036 52040
rect 21140 52009 21168 52040
rect 21361 52037 21373 52071
rect 21407 52068 21419 52071
rect 21450 52068 21456 52080
rect 21407 52040 21456 52068
rect 21407 52037 21419 52040
rect 21361 52031 21419 52037
rect 21450 52028 21456 52040
rect 21508 52068 21514 52080
rect 25682 52068 25688 52080
rect 21508 52040 25688 52068
rect 21508 52028 21514 52040
rect 25682 52028 25688 52040
rect 25740 52028 25746 52080
rect 21140 52003 21206 52009
rect 21140 51972 21160 52003
rect 21148 51969 21160 51972
rect 21194 51969 21206 52003
rect 21148 51963 21206 51969
rect 21269 52003 21327 52009
rect 21269 51969 21281 52003
rect 21315 51969 21327 52003
rect 21269 51963 21327 51969
rect 20732 51904 21036 51932
rect 21284 51932 21312 51963
rect 21542 51960 21548 52012
rect 21600 51960 21606 52012
rect 38286 52000 38292 52012
rect 22066 51972 38292 52000
rect 21634 51932 21640 51944
rect 21284 51904 21640 51932
rect 10778 51864 10784 51876
rect 4724 51836 10784 51864
rect 10778 51824 10784 51836
rect 10836 51824 10842 51876
rect 4982 51756 4988 51808
rect 5040 51796 5046 51808
rect 20640 51796 20668 51892
rect 20732 51864 20760 51904
rect 21634 51892 21640 51904
rect 21692 51932 21698 51944
rect 22066 51932 22094 51972
rect 38286 51960 38292 51972
rect 38344 51960 38350 52012
rect 36262 51932 36268 51944
rect 21692 51904 22094 51932
rect 28966 51904 36268 51932
rect 21692 51892 21698 51904
rect 28966 51864 28994 51904
rect 36262 51892 36268 51904
rect 36320 51892 36326 51944
rect 20732 51836 28994 51864
rect 5040 51768 20668 51796
rect 20993 51799 21051 51805
rect 5040 51756 5046 51768
rect 20993 51765 21005 51799
rect 21039 51796 21051 51799
rect 21726 51796 21732 51808
rect 21039 51768 21732 51796
rect 21039 51765 21051 51768
rect 20993 51759 21051 51765
rect 21726 51756 21732 51768
rect 21784 51756 21790 51808
rect 1104 51706 40848 51728
rect 1104 51654 1950 51706
rect 2002 51654 2014 51706
rect 2066 51654 2078 51706
rect 2130 51654 2142 51706
rect 2194 51654 2206 51706
rect 2258 51654 6950 51706
rect 7002 51654 7014 51706
rect 7066 51654 7078 51706
rect 7130 51654 7142 51706
rect 7194 51654 7206 51706
rect 7258 51654 11950 51706
rect 12002 51654 12014 51706
rect 12066 51654 12078 51706
rect 12130 51654 12142 51706
rect 12194 51654 12206 51706
rect 12258 51654 16950 51706
rect 17002 51654 17014 51706
rect 17066 51654 17078 51706
rect 17130 51654 17142 51706
rect 17194 51654 17206 51706
rect 17258 51654 21950 51706
rect 22002 51654 22014 51706
rect 22066 51654 22078 51706
rect 22130 51654 22142 51706
rect 22194 51654 22206 51706
rect 22258 51654 26950 51706
rect 27002 51654 27014 51706
rect 27066 51654 27078 51706
rect 27130 51654 27142 51706
rect 27194 51654 27206 51706
rect 27258 51654 31950 51706
rect 32002 51654 32014 51706
rect 32066 51654 32078 51706
rect 32130 51654 32142 51706
rect 32194 51654 32206 51706
rect 32258 51654 36950 51706
rect 37002 51654 37014 51706
rect 37066 51654 37078 51706
rect 37130 51654 37142 51706
rect 37194 51654 37206 51706
rect 37258 51654 40848 51706
rect 1104 51632 40848 51654
rect 31754 51348 31760 51400
rect 31812 51348 31818 51400
rect 32677 51391 32735 51397
rect 32677 51357 32689 51391
rect 32723 51388 32735 51391
rect 36814 51388 36820 51400
rect 32723 51360 36820 51388
rect 32723 51357 32735 51360
rect 32677 51351 32735 51357
rect 36814 51348 36820 51360
rect 36872 51348 36878 51400
rect 6822 51280 6828 51332
rect 6880 51320 6886 51332
rect 30837 51323 30895 51329
rect 30837 51320 30849 51323
rect 6880 51292 30849 51320
rect 6880 51280 6886 51292
rect 30837 51289 30849 51292
rect 30883 51289 30895 51323
rect 30837 51283 30895 51289
rect 1104 51162 40848 51184
rect 1104 51110 2610 51162
rect 2662 51110 2674 51162
rect 2726 51110 2738 51162
rect 2790 51110 2802 51162
rect 2854 51110 2866 51162
rect 2918 51110 7610 51162
rect 7662 51110 7674 51162
rect 7726 51110 7738 51162
rect 7790 51110 7802 51162
rect 7854 51110 7866 51162
rect 7918 51110 12610 51162
rect 12662 51110 12674 51162
rect 12726 51110 12738 51162
rect 12790 51110 12802 51162
rect 12854 51110 12866 51162
rect 12918 51110 17610 51162
rect 17662 51110 17674 51162
rect 17726 51110 17738 51162
rect 17790 51110 17802 51162
rect 17854 51110 17866 51162
rect 17918 51110 22610 51162
rect 22662 51110 22674 51162
rect 22726 51110 22738 51162
rect 22790 51110 22802 51162
rect 22854 51110 22866 51162
rect 22918 51110 27610 51162
rect 27662 51110 27674 51162
rect 27726 51110 27738 51162
rect 27790 51110 27802 51162
rect 27854 51110 27866 51162
rect 27918 51110 32610 51162
rect 32662 51110 32674 51162
rect 32726 51110 32738 51162
rect 32790 51110 32802 51162
rect 32854 51110 32866 51162
rect 32918 51110 37610 51162
rect 37662 51110 37674 51162
rect 37726 51110 37738 51162
rect 37790 51110 37802 51162
rect 37854 51110 37866 51162
rect 37918 51110 40848 51162
rect 1104 51088 40848 51110
rect 8202 51008 8208 51060
rect 8260 51048 8266 51060
rect 10137 51051 10195 51057
rect 10137 51048 10149 51051
rect 8260 51020 10149 51048
rect 8260 51008 8266 51020
rect 10137 51017 10149 51020
rect 10183 51017 10195 51051
rect 10137 51011 10195 51017
rect 12463 51051 12521 51057
rect 12463 51017 12475 51051
rect 12509 51048 12521 51051
rect 13446 51048 13452 51060
rect 12509 51020 13452 51048
rect 12509 51017 12521 51020
rect 12463 51011 12521 51017
rect 13446 51008 13452 51020
rect 13504 51008 13510 51060
rect 22278 51008 22284 51060
rect 22336 51048 22342 51060
rect 23106 51048 23112 51060
rect 22336 51020 23112 51048
rect 22336 51008 22342 51020
rect 23106 51008 23112 51020
rect 23164 51008 23170 51060
rect 32398 51008 32404 51060
rect 32456 51048 32462 51060
rect 37458 51048 37464 51060
rect 32456 51020 37464 51048
rect 32456 51008 32462 51020
rect 37458 51008 37464 51020
rect 37516 51008 37522 51060
rect 11606 50940 11612 50992
rect 11664 50980 11670 50992
rect 12253 50983 12311 50989
rect 12253 50980 12265 50983
rect 11664 50952 12265 50980
rect 11664 50940 11670 50952
rect 12253 50949 12265 50952
rect 12299 50949 12311 50983
rect 12253 50943 12311 50949
rect 22097 50983 22155 50989
rect 22097 50949 22109 50983
rect 22143 50980 22155 50983
rect 22370 50980 22376 50992
rect 22143 50952 22376 50980
rect 22143 50949 22155 50952
rect 22097 50943 22155 50949
rect 22370 50940 22376 50952
rect 22428 50940 22434 50992
rect 7926 50872 7932 50924
rect 7984 50912 7990 50924
rect 8202 50912 8208 50924
rect 7984 50884 8208 50912
rect 7984 50872 7990 50884
rect 8202 50872 8208 50884
rect 8260 50872 8266 50924
rect 10686 50872 10692 50924
rect 10744 50872 10750 50924
rect 10870 50872 10876 50924
rect 10928 50872 10934 50924
rect 12986 50921 12992 50924
rect 12955 50915 12992 50921
rect 12955 50881 12967 50915
rect 12955 50875 12992 50881
rect 12986 50872 12992 50875
rect 13044 50872 13050 50924
rect 21818 50872 21824 50924
rect 21876 50872 21882 50924
rect 22005 50915 22063 50921
rect 22005 50881 22017 50915
rect 22051 50881 22063 50915
rect 22005 50875 22063 50881
rect 22189 50915 22247 50921
rect 22189 50881 22201 50915
rect 22235 50881 22247 50915
rect 22189 50875 22247 50881
rect 11422 50804 11428 50856
rect 11480 50844 11486 50856
rect 13265 50847 13323 50853
rect 13265 50844 13277 50847
rect 11480 50816 13277 50844
rect 11480 50804 11486 50816
rect 13265 50813 13277 50816
rect 13311 50813 13323 50847
rect 13265 50807 13323 50813
rect 13357 50847 13415 50853
rect 13357 50813 13369 50847
rect 13403 50844 13415 50847
rect 17494 50844 17500 50856
rect 13403 50816 17500 50844
rect 13403 50813 13415 50816
rect 13357 50807 13415 50813
rect 17494 50804 17500 50816
rect 17552 50804 17558 50856
rect 21726 50804 21732 50856
rect 21784 50844 21790 50856
rect 22020 50844 22048 50875
rect 21784 50816 22048 50844
rect 22204 50844 22232 50875
rect 22278 50872 22284 50924
rect 22336 50872 22342 50924
rect 26142 50844 26148 50856
rect 22204 50816 26148 50844
rect 21784 50804 21790 50816
rect 26142 50804 26148 50816
rect 26200 50804 26206 50856
rect 12621 50779 12679 50785
rect 12621 50745 12633 50779
rect 12667 50776 12679 50779
rect 12667 50748 13308 50776
rect 12667 50745 12679 50748
rect 12621 50739 12679 50745
rect 13280 50720 13308 50748
rect 12434 50668 12440 50720
rect 12492 50668 12498 50720
rect 12802 50668 12808 50720
rect 12860 50668 12866 50720
rect 13262 50668 13268 50720
rect 13320 50668 13326 50720
rect 22465 50711 22523 50717
rect 22465 50677 22477 50711
rect 22511 50708 22523 50711
rect 23198 50708 23204 50720
rect 22511 50680 23204 50708
rect 22511 50677 22523 50680
rect 22465 50671 22523 50677
rect 23198 50668 23204 50680
rect 23256 50668 23262 50720
rect 1104 50618 40848 50640
rect 1104 50566 1950 50618
rect 2002 50566 2014 50618
rect 2066 50566 2078 50618
rect 2130 50566 2142 50618
rect 2194 50566 2206 50618
rect 2258 50566 6950 50618
rect 7002 50566 7014 50618
rect 7066 50566 7078 50618
rect 7130 50566 7142 50618
rect 7194 50566 7206 50618
rect 7258 50566 11950 50618
rect 12002 50566 12014 50618
rect 12066 50566 12078 50618
rect 12130 50566 12142 50618
rect 12194 50566 12206 50618
rect 12258 50566 16950 50618
rect 17002 50566 17014 50618
rect 17066 50566 17078 50618
rect 17130 50566 17142 50618
rect 17194 50566 17206 50618
rect 17258 50566 21950 50618
rect 22002 50566 22014 50618
rect 22066 50566 22078 50618
rect 22130 50566 22142 50618
rect 22194 50566 22206 50618
rect 22258 50566 26950 50618
rect 27002 50566 27014 50618
rect 27066 50566 27078 50618
rect 27130 50566 27142 50618
rect 27194 50566 27206 50618
rect 27258 50566 31950 50618
rect 32002 50566 32014 50618
rect 32066 50566 32078 50618
rect 32130 50566 32142 50618
rect 32194 50566 32206 50618
rect 32258 50566 36950 50618
rect 37002 50566 37014 50618
rect 37066 50566 37078 50618
rect 37130 50566 37142 50618
rect 37194 50566 37206 50618
rect 37258 50566 40848 50618
rect 1104 50544 40848 50566
rect 19886 50464 19892 50516
rect 19944 50504 19950 50516
rect 29822 50504 29828 50516
rect 19944 50476 29828 50504
rect 19944 50464 19950 50476
rect 29822 50464 29828 50476
rect 29880 50464 29886 50516
rect 2961 50439 3019 50445
rect 2961 50405 2973 50439
rect 3007 50436 3019 50439
rect 3050 50436 3056 50448
rect 3007 50408 3056 50436
rect 3007 50405 3019 50408
rect 2961 50399 3019 50405
rect 3050 50396 3056 50408
rect 3108 50396 3114 50448
rect 9214 50436 9220 50448
rect 3160 50408 9220 50436
rect 2225 50371 2283 50377
rect 2225 50337 2237 50371
rect 2271 50368 2283 50371
rect 3160 50368 3188 50408
rect 9214 50396 9220 50408
rect 9272 50436 9278 50448
rect 10594 50436 10600 50448
rect 9272 50408 10600 50436
rect 9272 50396 9278 50408
rect 10594 50396 10600 50408
rect 10652 50396 10658 50448
rect 14182 50396 14188 50448
rect 14240 50436 14246 50448
rect 20622 50436 20628 50448
rect 14240 50408 20628 50436
rect 14240 50396 14246 50408
rect 20622 50396 20628 50408
rect 20680 50396 20686 50448
rect 23474 50396 23480 50448
rect 23532 50436 23538 50448
rect 35250 50436 35256 50448
rect 23532 50408 35256 50436
rect 23532 50396 23538 50408
rect 35250 50396 35256 50408
rect 35308 50396 35314 50448
rect 2271 50340 3188 50368
rect 3237 50371 3295 50377
rect 2271 50337 2283 50340
rect 2225 50331 2283 50337
rect 3237 50337 3249 50371
rect 3283 50368 3295 50371
rect 8018 50368 8024 50380
rect 3283 50340 8024 50368
rect 3283 50337 3295 50340
rect 3237 50331 3295 50337
rect 8018 50328 8024 50340
rect 8076 50368 8082 50380
rect 8202 50368 8208 50380
rect 8076 50340 8208 50368
rect 8076 50328 8082 50340
rect 8202 50328 8208 50340
rect 8260 50328 8266 50380
rect 39666 50368 39672 50380
rect 22066 50340 39672 50368
rect 2501 50303 2559 50309
rect 2501 50269 2513 50303
rect 2547 50269 2559 50303
rect 8938 50300 8944 50312
rect 2501 50263 2559 50269
rect 3344 50272 8944 50300
rect 2516 50232 2544 50263
rect 3344 50232 3372 50272
rect 8938 50260 8944 50272
rect 8996 50260 9002 50312
rect 12802 50300 12808 50312
rect 9876 50272 12808 50300
rect 2516 50204 3372 50232
rect 6730 50192 6736 50244
rect 6788 50232 6794 50244
rect 9876 50232 9904 50272
rect 12802 50260 12808 50272
rect 12860 50260 12866 50312
rect 20530 50260 20536 50312
rect 20588 50300 20594 50312
rect 22066 50300 22094 50340
rect 39666 50328 39672 50340
rect 39724 50328 39730 50380
rect 20588 50272 22094 50300
rect 20588 50260 20594 50272
rect 6788 50204 9904 50232
rect 6788 50192 6794 50204
rect 11606 50192 11612 50244
rect 11664 50232 11670 50244
rect 12529 50235 12587 50241
rect 12529 50232 12541 50235
rect 11664 50204 12541 50232
rect 11664 50192 11670 50204
rect 12529 50201 12541 50204
rect 12575 50201 12587 50235
rect 12529 50195 12587 50201
rect 12621 50167 12679 50173
rect 12621 50133 12633 50167
rect 12667 50164 12679 50167
rect 25590 50164 25596 50176
rect 12667 50136 25596 50164
rect 12667 50133 12679 50136
rect 12621 50127 12679 50133
rect 25590 50124 25596 50136
rect 25648 50124 25654 50176
rect 1104 50074 40848 50096
rect 1104 50022 2610 50074
rect 2662 50022 2674 50074
rect 2726 50022 2738 50074
rect 2790 50022 2802 50074
rect 2854 50022 2866 50074
rect 2918 50022 7610 50074
rect 7662 50022 7674 50074
rect 7726 50022 7738 50074
rect 7790 50022 7802 50074
rect 7854 50022 7866 50074
rect 7918 50022 12610 50074
rect 12662 50022 12674 50074
rect 12726 50022 12738 50074
rect 12790 50022 12802 50074
rect 12854 50022 12866 50074
rect 12918 50022 17610 50074
rect 17662 50022 17674 50074
rect 17726 50022 17738 50074
rect 17790 50022 17802 50074
rect 17854 50022 17866 50074
rect 17918 50022 22610 50074
rect 22662 50022 22674 50074
rect 22726 50022 22738 50074
rect 22790 50022 22802 50074
rect 22854 50022 22866 50074
rect 22918 50022 27610 50074
rect 27662 50022 27674 50074
rect 27726 50022 27738 50074
rect 27790 50022 27802 50074
rect 27854 50022 27866 50074
rect 27918 50022 32610 50074
rect 32662 50022 32674 50074
rect 32726 50022 32738 50074
rect 32790 50022 32802 50074
rect 32854 50022 32866 50074
rect 32918 50022 37610 50074
rect 37662 50022 37674 50074
rect 37726 50022 37738 50074
rect 37790 50022 37802 50074
rect 37854 50022 37866 50074
rect 37918 50022 40848 50074
rect 1104 50000 40848 50022
rect 3878 49920 3884 49972
rect 3936 49960 3942 49972
rect 3936 49932 16574 49960
rect 3936 49920 3942 49932
rect 2593 49895 2651 49901
rect 2593 49861 2605 49895
rect 2639 49892 2651 49895
rect 7282 49892 7288 49904
rect 2639 49864 7288 49892
rect 2639 49861 2651 49864
rect 2593 49855 2651 49861
rect 7282 49852 7288 49864
rect 7340 49852 7346 49904
rect 16546 49892 16574 49932
rect 23106 49920 23112 49972
rect 23164 49960 23170 49972
rect 23164 49932 23704 49960
rect 23164 49920 23170 49932
rect 23676 49892 23704 49932
rect 39669 49895 39727 49901
rect 39669 49892 39681 49895
rect 16546 49864 23612 49892
rect 23676 49864 39681 49892
rect 1394 49784 1400 49836
rect 1452 49784 1458 49836
rect 13906 49784 13912 49836
rect 13964 49784 13970 49836
rect 14182 49784 14188 49836
rect 14240 49784 14246 49836
rect 23584 49768 23612 49864
rect 23768 49836 23796 49864
rect 39669 49861 39681 49864
rect 39715 49861 39727 49895
rect 39669 49855 39727 49861
rect 23658 49784 23664 49836
rect 23716 49784 23722 49836
rect 23750 49784 23756 49836
rect 23808 49784 23814 49836
rect 23937 49827 23995 49833
rect 23937 49793 23949 49827
rect 23983 49793 23995 49827
rect 23937 49787 23995 49793
rect 8938 49716 8944 49768
rect 8996 49756 9002 49768
rect 11146 49756 11152 49768
rect 8996 49728 11152 49756
rect 8996 49716 9002 49728
rect 11146 49716 11152 49728
rect 11204 49756 11210 49768
rect 14277 49759 14335 49765
rect 14277 49756 14289 49759
rect 11204 49728 14289 49756
rect 11204 49716 11210 49728
rect 14277 49725 14289 49728
rect 14323 49725 14335 49759
rect 14277 49719 14335 49725
rect 22370 49716 22376 49768
rect 22428 49756 22434 49768
rect 23106 49756 23112 49768
rect 22428 49728 23112 49756
rect 22428 49716 22434 49728
rect 23106 49716 23112 49728
rect 23164 49716 23170 49768
rect 23566 49716 23572 49768
rect 23624 49756 23630 49768
rect 23952 49756 23980 49787
rect 24302 49784 24308 49836
rect 24360 49784 24366 49836
rect 24670 49784 24676 49836
rect 24728 49784 24734 49836
rect 33778 49784 33784 49836
rect 33836 49784 33842 49836
rect 35802 49784 35808 49836
rect 35860 49784 35866 49836
rect 36357 49827 36415 49833
rect 36357 49793 36369 49827
rect 36403 49793 36415 49827
rect 36357 49787 36415 49793
rect 23624 49728 23980 49756
rect 23624 49716 23630 49728
rect 25038 49716 25044 49768
rect 25096 49716 25102 49768
rect 31570 49716 31576 49768
rect 31628 49756 31634 49768
rect 33796 49756 33824 49784
rect 36372 49756 36400 49787
rect 36630 49784 36636 49836
rect 36688 49784 36694 49836
rect 40494 49784 40500 49836
rect 40552 49784 40558 49836
rect 31628 49728 36400 49756
rect 31628 49716 31634 49728
rect 13078 49648 13084 49700
rect 13136 49688 13142 49700
rect 13354 49688 13360 49700
rect 13136 49660 13360 49688
rect 13136 49648 13142 49660
rect 13354 49648 13360 49660
rect 13412 49688 13418 49700
rect 29546 49688 29552 49700
rect 13412 49660 29552 49688
rect 13412 49648 13418 49660
rect 29546 49648 29552 49660
rect 29604 49648 29610 49700
rect 33778 49648 33784 49700
rect 33836 49688 33842 49700
rect 34146 49688 34152 49700
rect 33836 49660 34152 49688
rect 33836 49648 33842 49660
rect 34146 49648 34152 49660
rect 34204 49688 34210 49700
rect 35989 49691 36047 49697
rect 35989 49688 36001 49691
rect 34204 49660 36001 49688
rect 34204 49648 34210 49660
rect 35989 49657 36001 49660
rect 36035 49657 36047 49691
rect 35989 49651 36047 49657
rect 1104 49530 40848 49552
rect 1104 49478 1950 49530
rect 2002 49478 2014 49530
rect 2066 49478 2078 49530
rect 2130 49478 2142 49530
rect 2194 49478 2206 49530
rect 2258 49478 6950 49530
rect 7002 49478 7014 49530
rect 7066 49478 7078 49530
rect 7130 49478 7142 49530
rect 7194 49478 7206 49530
rect 7258 49478 11950 49530
rect 12002 49478 12014 49530
rect 12066 49478 12078 49530
rect 12130 49478 12142 49530
rect 12194 49478 12206 49530
rect 12258 49478 16950 49530
rect 17002 49478 17014 49530
rect 17066 49478 17078 49530
rect 17130 49478 17142 49530
rect 17194 49478 17206 49530
rect 17258 49478 21950 49530
rect 22002 49478 22014 49530
rect 22066 49478 22078 49530
rect 22130 49478 22142 49530
rect 22194 49478 22206 49530
rect 22258 49478 26950 49530
rect 27002 49478 27014 49530
rect 27066 49478 27078 49530
rect 27130 49478 27142 49530
rect 27194 49478 27206 49530
rect 27258 49478 31950 49530
rect 32002 49478 32014 49530
rect 32066 49478 32078 49530
rect 32130 49478 32142 49530
rect 32194 49478 32206 49530
rect 32258 49478 36950 49530
rect 37002 49478 37014 49530
rect 37066 49478 37078 49530
rect 37130 49478 37142 49530
rect 37194 49478 37206 49530
rect 37258 49478 40848 49530
rect 1104 49456 40848 49478
rect 22278 49308 22284 49360
rect 22336 49348 22342 49360
rect 23474 49348 23480 49360
rect 22336 49320 23480 49348
rect 22336 49308 22342 49320
rect 23474 49308 23480 49320
rect 23532 49348 23538 49360
rect 23532 49320 24808 49348
rect 23532 49308 23538 49320
rect 20162 49240 20168 49292
rect 20220 49280 20226 49292
rect 20220 49252 24532 49280
rect 20220 49240 20226 49252
rect 24394 49172 24400 49224
rect 24452 49172 24458 49224
rect 24504 49212 24532 49252
rect 24504 49184 24716 49212
rect 19242 49036 19248 49088
rect 19300 49076 19306 49088
rect 24688 49085 24716 49184
rect 24780 49153 24808 49320
rect 24765 49147 24823 49153
rect 24765 49113 24777 49147
rect 24811 49144 24823 49147
rect 37366 49144 37372 49156
rect 24811 49116 37372 49144
rect 24811 49113 24823 49116
rect 24765 49107 24823 49113
rect 37366 49104 37372 49116
rect 37424 49104 37430 49156
rect 24581 49079 24639 49085
rect 24581 49076 24593 49079
rect 19300 49048 24593 49076
rect 19300 49036 19306 49048
rect 24581 49045 24593 49048
rect 24627 49045 24639 49079
rect 24581 49039 24639 49045
rect 24673 49079 24731 49085
rect 24673 49045 24685 49079
rect 24719 49045 24731 49079
rect 24673 49039 24731 49045
rect 24854 49036 24860 49088
rect 24912 49036 24918 49088
rect 1104 48986 40848 49008
rect 1104 48934 2610 48986
rect 2662 48934 2674 48986
rect 2726 48934 2738 48986
rect 2790 48934 2802 48986
rect 2854 48934 2866 48986
rect 2918 48934 7610 48986
rect 7662 48934 7674 48986
rect 7726 48934 7738 48986
rect 7790 48934 7802 48986
rect 7854 48934 7866 48986
rect 7918 48934 12610 48986
rect 12662 48934 12674 48986
rect 12726 48934 12738 48986
rect 12790 48934 12802 48986
rect 12854 48934 12866 48986
rect 12918 48934 17610 48986
rect 17662 48934 17674 48986
rect 17726 48934 17738 48986
rect 17790 48934 17802 48986
rect 17854 48934 17866 48986
rect 17918 48934 22610 48986
rect 22662 48934 22674 48986
rect 22726 48934 22738 48986
rect 22790 48934 22802 48986
rect 22854 48934 22866 48986
rect 22918 48934 27610 48986
rect 27662 48934 27674 48986
rect 27726 48934 27738 48986
rect 27790 48934 27802 48986
rect 27854 48934 27866 48986
rect 27918 48934 32610 48986
rect 32662 48934 32674 48986
rect 32726 48934 32738 48986
rect 32790 48934 32802 48986
rect 32854 48934 32866 48986
rect 32918 48934 37610 48986
rect 37662 48934 37674 48986
rect 37726 48934 37738 48986
rect 37790 48934 37802 48986
rect 37854 48934 37866 48986
rect 37918 48934 40848 48986
rect 1104 48912 40848 48934
rect 16574 48832 16580 48884
rect 16632 48872 16638 48884
rect 17313 48875 17371 48881
rect 17313 48872 17325 48875
rect 16632 48844 17325 48872
rect 16632 48832 16638 48844
rect 17313 48841 17325 48844
rect 17359 48841 17371 48875
rect 17313 48835 17371 48841
rect 37366 48832 37372 48884
rect 37424 48832 37430 48884
rect 13354 48804 13360 48816
rect 10244 48776 13360 48804
rect 10244 48745 10272 48776
rect 13354 48764 13360 48776
rect 13412 48764 13418 48816
rect 19978 48804 19984 48816
rect 16776 48776 19984 48804
rect 10229 48739 10287 48745
rect 10229 48705 10241 48739
rect 10275 48705 10287 48739
rect 10229 48699 10287 48705
rect 10413 48739 10471 48745
rect 10413 48705 10425 48739
rect 10459 48736 10471 48739
rect 11422 48736 11428 48748
rect 10459 48708 11428 48736
rect 10459 48705 10471 48708
rect 10413 48699 10471 48705
rect 11422 48696 11428 48708
rect 11480 48696 11486 48748
rect 16776 48745 16804 48776
rect 19978 48764 19984 48776
rect 20036 48764 20042 48816
rect 16761 48739 16819 48745
rect 16761 48705 16773 48739
rect 16807 48705 16819 48739
rect 16761 48699 16819 48705
rect 17037 48739 17095 48745
rect 17037 48705 17049 48739
rect 17083 48705 17095 48739
rect 17037 48699 17095 48705
rect 17129 48739 17187 48745
rect 17129 48705 17141 48739
rect 17175 48736 17187 48739
rect 17310 48736 17316 48748
rect 17175 48708 17316 48736
rect 17175 48705 17187 48708
rect 17129 48699 17187 48705
rect 8938 48628 8944 48680
rect 8996 48668 9002 48680
rect 10781 48671 10839 48677
rect 10781 48668 10793 48671
rect 8996 48640 10793 48668
rect 8996 48628 9002 48640
rect 10781 48637 10793 48640
rect 10827 48668 10839 48671
rect 11514 48668 11520 48680
rect 10827 48640 11520 48668
rect 10827 48637 10839 48640
rect 10781 48631 10839 48637
rect 11514 48628 11520 48640
rect 11572 48668 11578 48680
rect 16942 48668 16948 48680
rect 11572 48640 16948 48668
rect 11572 48628 11578 48640
rect 16942 48628 16948 48640
rect 17000 48628 17006 48680
rect 17052 48668 17080 48699
rect 17310 48696 17316 48708
rect 17368 48696 17374 48748
rect 22370 48696 22376 48748
rect 22428 48696 22434 48748
rect 22557 48739 22615 48745
rect 22557 48705 22569 48739
rect 22603 48736 22615 48739
rect 24118 48736 24124 48748
rect 22603 48708 24124 48736
rect 22603 48705 22615 48708
rect 22557 48699 22615 48705
rect 24118 48696 24124 48708
rect 24176 48696 24182 48748
rect 32950 48696 32956 48748
rect 33008 48736 33014 48748
rect 37277 48739 37335 48745
rect 37277 48736 37289 48739
rect 33008 48708 37289 48736
rect 33008 48696 33014 48708
rect 37277 48705 37289 48708
rect 37323 48705 37335 48739
rect 37829 48739 37887 48745
rect 37829 48736 37841 48739
rect 37277 48699 37335 48705
rect 37476 48708 37841 48736
rect 37476 48680 37504 48708
rect 37829 48705 37841 48708
rect 37875 48736 37887 48739
rect 38378 48736 38384 48748
rect 37875 48708 38384 48736
rect 37875 48705 37887 48708
rect 37829 48699 37887 48705
rect 38378 48696 38384 48708
rect 38436 48696 38442 48748
rect 17402 48668 17408 48680
rect 17052 48640 17408 48668
rect 17402 48628 17408 48640
rect 17460 48628 17466 48680
rect 37458 48628 37464 48680
rect 37516 48628 37522 48680
rect 10686 48560 10692 48612
rect 10744 48560 10750 48612
rect 13722 48560 13728 48612
rect 13780 48600 13786 48612
rect 22465 48603 22523 48609
rect 22465 48600 22477 48603
rect 13780 48572 22477 48600
rect 13780 48560 13786 48572
rect 22465 48569 22477 48572
rect 22511 48569 22523 48603
rect 22465 48563 22523 48569
rect 11422 48492 11428 48544
rect 11480 48532 11486 48544
rect 16758 48532 16764 48544
rect 11480 48504 16764 48532
rect 11480 48492 11486 48504
rect 16758 48492 16764 48504
rect 16816 48492 16822 48544
rect 16853 48535 16911 48541
rect 16853 48501 16865 48535
rect 16899 48532 16911 48535
rect 16942 48532 16948 48544
rect 16899 48504 16948 48532
rect 16899 48501 16911 48504
rect 16853 48495 16911 48501
rect 16942 48492 16948 48504
rect 17000 48532 17006 48544
rect 22278 48532 22284 48544
rect 17000 48504 22284 48532
rect 17000 48492 17006 48504
rect 22278 48492 22284 48504
rect 22336 48492 22342 48544
rect 1104 48442 40848 48464
rect 1104 48390 1950 48442
rect 2002 48390 2014 48442
rect 2066 48390 2078 48442
rect 2130 48390 2142 48442
rect 2194 48390 2206 48442
rect 2258 48390 6950 48442
rect 7002 48390 7014 48442
rect 7066 48390 7078 48442
rect 7130 48390 7142 48442
rect 7194 48390 7206 48442
rect 7258 48390 11950 48442
rect 12002 48390 12014 48442
rect 12066 48390 12078 48442
rect 12130 48390 12142 48442
rect 12194 48390 12206 48442
rect 12258 48390 16950 48442
rect 17002 48390 17014 48442
rect 17066 48390 17078 48442
rect 17130 48390 17142 48442
rect 17194 48390 17206 48442
rect 17258 48390 21950 48442
rect 22002 48390 22014 48442
rect 22066 48390 22078 48442
rect 22130 48390 22142 48442
rect 22194 48390 22206 48442
rect 22258 48390 26950 48442
rect 27002 48390 27014 48442
rect 27066 48390 27078 48442
rect 27130 48390 27142 48442
rect 27194 48390 27206 48442
rect 27258 48390 31950 48442
rect 32002 48390 32014 48442
rect 32066 48390 32078 48442
rect 32130 48390 32142 48442
rect 32194 48390 32206 48442
rect 32258 48390 36950 48442
rect 37002 48390 37014 48442
rect 37066 48390 37078 48442
rect 37130 48390 37142 48442
rect 37194 48390 37206 48442
rect 37258 48390 40848 48442
rect 1104 48368 40848 48390
rect 13538 48288 13544 48340
rect 13596 48328 13602 48340
rect 24854 48328 24860 48340
rect 13596 48300 24860 48328
rect 13596 48288 13602 48300
rect 24854 48288 24860 48300
rect 24912 48288 24918 48340
rect 10502 48220 10508 48272
rect 10560 48260 10566 48272
rect 11330 48260 11336 48272
rect 10560 48232 11336 48260
rect 10560 48220 10566 48232
rect 11330 48220 11336 48232
rect 11388 48220 11394 48272
rect 14090 48084 14096 48136
rect 14148 48124 14154 48136
rect 19150 48124 19156 48136
rect 14148 48096 19156 48124
rect 14148 48084 14154 48096
rect 19150 48084 19156 48096
rect 19208 48084 19214 48136
rect 6454 47948 6460 48000
rect 6512 47988 6518 48000
rect 14734 47988 14740 48000
rect 6512 47960 14740 47988
rect 6512 47948 6518 47960
rect 14734 47948 14740 47960
rect 14792 47948 14798 48000
rect 19150 47948 19156 48000
rect 19208 47988 19214 48000
rect 38838 47988 38844 48000
rect 19208 47960 38844 47988
rect 19208 47948 19214 47960
rect 38838 47948 38844 47960
rect 38896 47948 38902 48000
rect 1104 47898 40848 47920
rect 1104 47846 2610 47898
rect 2662 47846 2674 47898
rect 2726 47846 2738 47898
rect 2790 47846 2802 47898
rect 2854 47846 2866 47898
rect 2918 47846 7610 47898
rect 7662 47846 7674 47898
rect 7726 47846 7738 47898
rect 7790 47846 7802 47898
rect 7854 47846 7866 47898
rect 7918 47846 12610 47898
rect 12662 47846 12674 47898
rect 12726 47846 12738 47898
rect 12790 47846 12802 47898
rect 12854 47846 12866 47898
rect 12918 47846 17610 47898
rect 17662 47846 17674 47898
rect 17726 47846 17738 47898
rect 17790 47846 17802 47898
rect 17854 47846 17866 47898
rect 17918 47846 22610 47898
rect 22662 47846 22674 47898
rect 22726 47846 22738 47898
rect 22790 47846 22802 47898
rect 22854 47846 22866 47898
rect 22918 47846 27610 47898
rect 27662 47846 27674 47898
rect 27726 47846 27738 47898
rect 27790 47846 27802 47898
rect 27854 47846 27866 47898
rect 27918 47846 32610 47898
rect 32662 47846 32674 47898
rect 32726 47846 32738 47898
rect 32790 47846 32802 47898
rect 32854 47846 32866 47898
rect 32918 47846 37610 47898
rect 37662 47846 37674 47898
rect 37726 47846 37738 47898
rect 37790 47846 37802 47898
rect 37854 47846 37866 47898
rect 37918 47846 40848 47898
rect 1104 47824 40848 47846
rect 14458 47744 14464 47796
rect 14516 47784 14522 47796
rect 38838 47784 38844 47796
rect 14516 47756 38844 47784
rect 14516 47744 14522 47756
rect 38838 47744 38844 47756
rect 38896 47744 38902 47796
rect 9674 47676 9680 47728
rect 9732 47716 9738 47728
rect 35802 47716 35808 47728
rect 9732 47688 35808 47716
rect 9732 47676 9738 47688
rect 35802 47676 35808 47688
rect 35860 47676 35866 47728
rect 3970 47608 3976 47660
rect 4028 47648 4034 47660
rect 21818 47648 21824 47660
rect 4028 47620 21824 47648
rect 4028 47608 4034 47620
rect 21818 47608 21824 47620
rect 21876 47608 21882 47660
rect 27982 47608 27988 47660
rect 28040 47648 28046 47660
rect 31021 47651 31079 47657
rect 31021 47648 31033 47651
rect 28040 47620 31033 47648
rect 28040 47608 28046 47620
rect 31021 47617 31033 47620
rect 31067 47617 31079 47651
rect 31021 47611 31079 47617
rect 2314 47540 2320 47592
rect 2372 47580 2378 47592
rect 28166 47580 28172 47592
rect 2372 47552 28172 47580
rect 2372 47540 2378 47552
rect 28166 47540 28172 47552
rect 28224 47540 28230 47592
rect 29914 47540 29920 47592
rect 29972 47580 29978 47592
rect 31757 47583 31815 47589
rect 31757 47580 31769 47583
rect 29972 47552 31769 47580
rect 29972 47540 29978 47552
rect 31757 47549 31769 47552
rect 31803 47549 31815 47583
rect 31757 47543 31815 47549
rect 1104 47354 40848 47376
rect 1104 47302 1950 47354
rect 2002 47302 2014 47354
rect 2066 47302 2078 47354
rect 2130 47302 2142 47354
rect 2194 47302 2206 47354
rect 2258 47302 6950 47354
rect 7002 47302 7014 47354
rect 7066 47302 7078 47354
rect 7130 47302 7142 47354
rect 7194 47302 7206 47354
rect 7258 47302 11950 47354
rect 12002 47302 12014 47354
rect 12066 47302 12078 47354
rect 12130 47302 12142 47354
rect 12194 47302 12206 47354
rect 12258 47302 16950 47354
rect 17002 47302 17014 47354
rect 17066 47302 17078 47354
rect 17130 47302 17142 47354
rect 17194 47302 17206 47354
rect 17258 47302 21950 47354
rect 22002 47302 22014 47354
rect 22066 47302 22078 47354
rect 22130 47302 22142 47354
rect 22194 47302 22206 47354
rect 22258 47302 26950 47354
rect 27002 47302 27014 47354
rect 27066 47302 27078 47354
rect 27130 47302 27142 47354
rect 27194 47302 27206 47354
rect 27258 47302 31950 47354
rect 32002 47302 32014 47354
rect 32066 47302 32078 47354
rect 32130 47302 32142 47354
rect 32194 47302 32206 47354
rect 32258 47302 36950 47354
rect 37002 47302 37014 47354
rect 37066 47302 37078 47354
rect 37130 47302 37142 47354
rect 37194 47302 37206 47354
rect 37258 47302 40848 47354
rect 1104 47280 40848 47302
rect 25866 46928 25872 46980
rect 25924 46968 25930 46980
rect 31294 46968 31300 46980
rect 25924 46940 31300 46968
rect 25924 46928 25930 46940
rect 31294 46928 31300 46940
rect 31352 46928 31358 46980
rect 1104 46810 40848 46832
rect 1104 46758 2610 46810
rect 2662 46758 2674 46810
rect 2726 46758 2738 46810
rect 2790 46758 2802 46810
rect 2854 46758 2866 46810
rect 2918 46758 7610 46810
rect 7662 46758 7674 46810
rect 7726 46758 7738 46810
rect 7790 46758 7802 46810
rect 7854 46758 7866 46810
rect 7918 46758 12610 46810
rect 12662 46758 12674 46810
rect 12726 46758 12738 46810
rect 12790 46758 12802 46810
rect 12854 46758 12866 46810
rect 12918 46758 17610 46810
rect 17662 46758 17674 46810
rect 17726 46758 17738 46810
rect 17790 46758 17802 46810
rect 17854 46758 17866 46810
rect 17918 46758 22610 46810
rect 22662 46758 22674 46810
rect 22726 46758 22738 46810
rect 22790 46758 22802 46810
rect 22854 46758 22866 46810
rect 22918 46758 27610 46810
rect 27662 46758 27674 46810
rect 27726 46758 27738 46810
rect 27790 46758 27802 46810
rect 27854 46758 27866 46810
rect 27918 46758 32610 46810
rect 32662 46758 32674 46810
rect 32726 46758 32738 46810
rect 32790 46758 32802 46810
rect 32854 46758 32866 46810
rect 32918 46758 37610 46810
rect 37662 46758 37674 46810
rect 37726 46758 37738 46810
rect 37790 46758 37802 46810
rect 37854 46758 37866 46810
rect 37918 46758 40848 46810
rect 1104 46736 40848 46758
rect 14458 46520 14464 46572
rect 14516 46560 14522 46572
rect 22370 46560 22376 46572
rect 14516 46532 22376 46560
rect 14516 46520 14522 46532
rect 22370 46520 22376 46532
rect 22428 46520 22434 46572
rect 20622 46452 20628 46504
rect 20680 46492 20686 46504
rect 30374 46492 30380 46504
rect 20680 46464 30380 46492
rect 20680 46452 20686 46464
rect 30374 46452 30380 46464
rect 30432 46452 30438 46504
rect 10318 46384 10324 46436
rect 10376 46424 10382 46436
rect 20346 46424 20352 46436
rect 10376 46396 20352 46424
rect 10376 46384 10382 46396
rect 20346 46384 20352 46396
rect 20404 46384 20410 46436
rect 22370 46384 22376 46436
rect 22428 46424 22434 46436
rect 23014 46424 23020 46436
rect 22428 46396 23020 46424
rect 22428 46384 22434 46396
rect 23014 46384 23020 46396
rect 23072 46384 23078 46436
rect 23198 46384 23204 46436
rect 23256 46424 23262 46436
rect 39482 46424 39488 46436
rect 23256 46396 39488 46424
rect 23256 46384 23262 46396
rect 39482 46384 39488 46396
rect 39540 46384 39546 46436
rect 10778 46316 10784 46368
rect 10836 46356 10842 46368
rect 36722 46356 36728 46368
rect 10836 46328 36728 46356
rect 10836 46316 10842 46328
rect 36722 46316 36728 46328
rect 36780 46316 36786 46368
rect 1104 46266 40848 46288
rect 1104 46214 1950 46266
rect 2002 46214 2014 46266
rect 2066 46214 2078 46266
rect 2130 46214 2142 46266
rect 2194 46214 2206 46266
rect 2258 46214 6950 46266
rect 7002 46214 7014 46266
rect 7066 46214 7078 46266
rect 7130 46214 7142 46266
rect 7194 46214 7206 46266
rect 7258 46214 11950 46266
rect 12002 46214 12014 46266
rect 12066 46214 12078 46266
rect 12130 46214 12142 46266
rect 12194 46214 12206 46266
rect 12258 46214 16950 46266
rect 17002 46214 17014 46266
rect 17066 46214 17078 46266
rect 17130 46214 17142 46266
rect 17194 46214 17206 46266
rect 17258 46214 21950 46266
rect 22002 46214 22014 46266
rect 22066 46214 22078 46266
rect 22130 46214 22142 46266
rect 22194 46214 22206 46266
rect 22258 46214 26950 46266
rect 27002 46214 27014 46266
rect 27066 46214 27078 46266
rect 27130 46214 27142 46266
rect 27194 46214 27206 46266
rect 27258 46214 31950 46266
rect 32002 46214 32014 46266
rect 32066 46214 32078 46266
rect 32130 46214 32142 46266
rect 32194 46214 32206 46266
rect 32258 46214 36950 46266
rect 37002 46214 37014 46266
rect 37066 46214 37078 46266
rect 37130 46214 37142 46266
rect 37194 46214 37206 46266
rect 37258 46214 40848 46266
rect 1104 46192 40848 46214
rect 23014 46112 23020 46164
rect 23072 46152 23078 46164
rect 23382 46152 23388 46164
rect 23072 46124 23388 46152
rect 23072 46112 23078 46124
rect 23382 46112 23388 46124
rect 23440 46112 23446 46164
rect 30374 45976 30380 46028
rect 30432 46016 30438 46028
rect 31294 46016 31300 46028
rect 30432 45988 31300 46016
rect 30432 45976 30438 45988
rect 31294 45976 31300 45988
rect 31352 46016 31358 46028
rect 32493 46019 32551 46025
rect 32493 46016 32505 46019
rect 31352 45988 32505 46016
rect 31352 45976 31358 45988
rect 32493 45985 32505 45988
rect 32539 45985 32551 46019
rect 32493 45979 32551 45985
rect 32125 45951 32183 45957
rect 32125 45948 32137 45951
rect 22066 45920 32137 45948
rect 18138 45840 18144 45892
rect 18196 45880 18202 45892
rect 22066 45880 22094 45920
rect 32125 45917 32137 45920
rect 32171 45917 32183 45951
rect 32125 45911 32183 45917
rect 32585 45951 32643 45957
rect 32585 45917 32597 45951
rect 32631 45917 32643 45951
rect 32585 45911 32643 45917
rect 18196 45852 22094 45880
rect 18196 45840 18202 45852
rect 31018 45840 31024 45892
rect 31076 45880 31082 45892
rect 32600 45880 32628 45911
rect 31076 45852 32628 45880
rect 31076 45840 31082 45852
rect 1104 45722 40848 45744
rect 1104 45670 2610 45722
rect 2662 45670 2674 45722
rect 2726 45670 2738 45722
rect 2790 45670 2802 45722
rect 2854 45670 2866 45722
rect 2918 45670 7610 45722
rect 7662 45670 7674 45722
rect 7726 45670 7738 45722
rect 7790 45670 7802 45722
rect 7854 45670 7866 45722
rect 7918 45670 12610 45722
rect 12662 45670 12674 45722
rect 12726 45670 12738 45722
rect 12790 45670 12802 45722
rect 12854 45670 12866 45722
rect 12918 45670 17610 45722
rect 17662 45670 17674 45722
rect 17726 45670 17738 45722
rect 17790 45670 17802 45722
rect 17854 45670 17866 45722
rect 17918 45670 22610 45722
rect 22662 45670 22674 45722
rect 22726 45670 22738 45722
rect 22790 45670 22802 45722
rect 22854 45670 22866 45722
rect 22918 45670 27610 45722
rect 27662 45670 27674 45722
rect 27726 45670 27738 45722
rect 27790 45670 27802 45722
rect 27854 45670 27866 45722
rect 27918 45670 32610 45722
rect 32662 45670 32674 45722
rect 32726 45670 32738 45722
rect 32790 45670 32802 45722
rect 32854 45670 32866 45722
rect 32918 45670 37610 45722
rect 37662 45670 37674 45722
rect 37726 45670 37738 45722
rect 37790 45670 37802 45722
rect 37854 45670 37866 45722
rect 37918 45670 40848 45722
rect 1104 45648 40848 45670
rect 20162 45540 20168 45552
rect 6748 45512 20168 45540
rect 3418 45432 3424 45484
rect 3476 45472 3482 45484
rect 6748 45481 6776 45512
rect 20162 45500 20168 45512
rect 20220 45500 20226 45552
rect 23198 45500 23204 45552
rect 23256 45540 23262 45552
rect 23750 45540 23756 45552
rect 23256 45512 23756 45540
rect 23256 45500 23262 45512
rect 23750 45500 23756 45512
rect 23808 45500 23814 45552
rect 6457 45475 6515 45481
rect 6457 45472 6469 45475
rect 3476 45444 6469 45472
rect 3476 45432 3482 45444
rect 6457 45441 6469 45444
rect 6503 45441 6515 45475
rect 6457 45435 6515 45441
rect 6733 45475 6791 45481
rect 6733 45441 6745 45475
rect 6779 45441 6791 45475
rect 6733 45435 6791 45441
rect 7469 45475 7527 45481
rect 7469 45441 7481 45475
rect 7515 45441 7527 45475
rect 7469 45435 7527 45441
rect 8205 45475 8263 45481
rect 8205 45441 8217 45475
rect 8251 45472 8263 45475
rect 8938 45472 8944 45484
rect 8251 45444 8944 45472
rect 8251 45441 8263 45444
rect 8205 45435 8263 45441
rect 7484 45404 7512 45435
rect 8938 45432 8944 45444
rect 8996 45432 9002 45484
rect 9030 45404 9036 45416
rect 7484 45376 9036 45404
rect 9030 45364 9036 45376
rect 9088 45364 9094 45416
rect 6454 45228 6460 45280
rect 6512 45268 6518 45280
rect 6641 45271 6699 45277
rect 6641 45268 6653 45271
rect 6512 45240 6653 45268
rect 6512 45228 6518 45240
rect 6641 45237 6653 45240
rect 6687 45237 6699 45271
rect 6641 45231 6699 45237
rect 20162 45228 20168 45280
rect 20220 45268 20226 45280
rect 24486 45268 24492 45280
rect 20220 45240 24492 45268
rect 20220 45228 20226 45240
rect 24486 45228 24492 45240
rect 24544 45228 24550 45280
rect 1104 45178 40848 45200
rect 1104 45126 1950 45178
rect 2002 45126 2014 45178
rect 2066 45126 2078 45178
rect 2130 45126 2142 45178
rect 2194 45126 2206 45178
rect 2258 45126 6950 45178
rect 7002 45126 7014 45178
rect 7066 45126 7078 45178
rect 7130 45126 7142 45178
rect 7194 45126 7206 45178
rect 7258 45126 11950 45178
rect 12002 45126 12014 45178
rect 12066 45126 12078 45178
rect 12130 45126 12142 45178
rect 12194 45126 12206 45178
rect 12258 45126 16950 45178
rect 17002 45126 17014 45178
rect 17066 45126 17078 45178
rect 17130 45126 17142 45178
rect 17194 45126 17206 45178
rect 17258 45126 21950 45178
rect 22002 45126 22014 45178
rect 22066 45126 22078 45178
rect 22130 45126 22142 45178
rect 22194 45126 22206 45178
rect 22258 45126 26950 45178
rect 27002 45126 27014 45178
rect 27066 45126 27078 45178
rect 27130 45126 27142 45178
rect 27194 45126 27206 45178
rect 27258 45126 31950 45178
rect 32002 45126 32014 45178
rect 32066 45126 32078 45178
rect 32130 45126 32142 45178
rect 32194 45126 32206 45178
rect 32258 45126 36950 45178
rect 37002 45126 37014 45178
rect 37066 45126 37078 45178
rect 37130 45126 37142 45178
rect 37194 45126 37206 45178
rect 37258 45126 40848 45178
rect 1104 45104 40848 45126
rect 10410 44956 10416 45008
rect 10468 44996 10474 45008
rect 19518 44996 19524 45008
rect 10468 44968 19524 44996
rect 10468 44956 10474 44968
rect 19518 44956 19524 44968
rect 19576 44956 19582 45008
rect 19628 44968 19932 44996
rect 12342 44888 12348 44940
rect 12400 44928 12406 44940
rect 19628 44928 19656 44968
rect 12400 44900 19656 44928
rect 12400 44888 12406 44900
rect 19794 44888 19800 44940
rect 19852 44888 19858 44940
rect 19904 44928 19932 44968
rect 21358 44956 21364 45008
rect 21416 44996 21422 45008
rect 38746 44996 38752 45008
rect 21416 44968 38752 44996
rect 21416 44956 21422 44968
rect 38746 44956 38752 44968
rect 38804 44956 38810 45008
rect 26878 44928 26884 44940
rect 19904 44900 26884 44928
rect 26878 44888 26884 44900
rect 26936 44888 26942 44940
rect 30098 44888 30104 44940
rect 30156 44928 30162 44940
rect 32398 44928 32404 44940
rect 30156 44900 32404 44928
rect 30156 44888 30162 44900
rect 32398 44888 32404 44900
rect 32456 44888 32462 44940
rect 6365 44863 6423 44869
rect 6365 44829 6377 44863
rect 6411 44860 6423 44863
rect 6454 44860 6460 44872
rect 6411 44832 6460 44860
rect 6411 44829 6423 44832
rect 6365 44823 6423 44829
rect 6454 44820 6460 44832
rect 6512 44820 6518 44872
rect 6730 44820 6736 44872
rect 6788 44820 6794 44872
rect 19613 44863 19671 44869
rect 19613 44829 19625 44863
rect 19659 44862 19671 44863
rect 19659 44860 19748 44862
rect 22370 44860 22376 44872
rect 19659 44834 22376 44860
rect 19659 44829 19671 44834
rect 19720 44832 22376 44834
rect 19613 44823 19671 44829
rect 22370 44820 22376 44832
rect 22428 44820 22434 44872
rect 32493 44863 32551 44869
rect 32493 44829 32505 44863
rect 32539 44829 32551 44863
rect 32493 44823 32551 44829
rect 31846 44792 31852 44804
rect 7498 44764 31852 44792
rect 31846 44752 31852 44764
rect 31904 44792 31910 44804
rect 32508 44792 32536 44823
rect 32582 44820 32588 44872
rect 32640 44860 32646 44872
rect 32861 44863 32919 44869
rect 32861 44860 32873 44863
rect 32640 44832 32873 44860
rect 32640 44820 32646 44832
rect 32861 44829 32873 44832
rect 32907 44829 32919 44863
rect 32861 44823 32919 44829
rect 31904 44764 32536 44792
rect 32769 44795 32827 44801
rect 31904 44752 31910 44764
rect 32769 44761 32781 44795
rect 32815 44761 32827 44795
rect 32769 44755 32827 44761
rect 19426 44684 19432 44736
rect 19484 44684 19490 44736
rect 32306 44684 32312 44736
rect 32364 44724 32370 44736
rect 32784 44724 32812 44755
rect 32364 44696 32812 44724
rect 32364 44684 32370 44696
rect 1104 44634 40848 44656
rect 1104 44582 2610 44634
rect 2662 44582 2674 44634
rect 2726 44582 2738 44634
rect 2790 44582 2802 44634
rect 2854 44582 2866 44634
rect 2918 44582 7610 44634
rect 7662 44582 7674 44634
rect 7726 44582 7738 44634
rect 7790 44582 7802 44634
rect 7854 44582 7866 44634
rect 7918 44582 12610 44634
rect 12662 44582 12674 44634
rect 12726 44582 12738 44634
rect 12790 44582 12802 44634
rect 12854 44582 12866 44634
rect 12918 44582 17610 44634
rect 17662 44582 17674 44634
rect 17726 44582 17738 44634
rect 17790 44582 17802 44634
rect 17854 44582 17866 44634
rect 17918 44582 22610 44634
rect 22662 44582 22674 44634
rect 22726 44582 22738 44634
rect 22790 44582 22802 44634
rect 22854 44582 22866 44634
rect 22918 44582 27610 44634
rect 27662 44582 27674 44634
rect 27726 44582 27738 44634
rect 27790 44582 27802 44634
rect 27854 44582 27866 44634
rect 27918 44582 32610 44634
rect 32662 44582 32674 44634
rect 32726 44582 32738 44634
rect 32790 44582 32802 44634
rect 32854 44582 32866 44634
rect 32918 44582 37610 44634
rect 37662 44582 37674 44634
rect 37726 44582 37738 44634
rect 37790 44582 37802 44634
rect 37854 44582 37866 44634
rect 37918 44582 40848 44634
rect 1104 44560 40848 44582
rect 18690 44480 18696 44532
rect 18748 44520 18754 44532
rect 19058 44520 19064 44532
rect 18748 44492 19064 44520
rect 18748 44480 18754 44492
rect 19058 44480 19064 44492
rect 19116 44480 19122 44532
rect 10413 44455 10471 44461
rect 10413 44421 10425 44455
rect 10459 44452 10471 44455
rect 12434 44452 12440 44464
rect 10459 44424 12440 44452
rect 10459 44421 10471 44424
rect 10413 44415 10471 44421
rect 12434 44412 12440 44424
rect 12492 44412 12498 44464
rect 18892 44424 22094 44452
rect 4709 44387 4767 44393
rect 4709 44353 4721 44387
rect 4755 44353 4767 44387
rect 4709 44347 4767 44353
rect 4985 44387 5043 44393
rect 4985 44353 4997 44387
rect 5031 44353 5043 44387
rect 4985 44347 5043 44353
rect 5169 44387 5227 44393
rect 5169 44353 5181 44387
rect 5215 44384 5227 44387
rect 9214 44384 9220 44396
rect 5215 44356 9220 44384
rect 5215 44353 5227 44356
rect 5169 44347 5227 44353
rect 4724 44248 4752 44347
rect 5000 44316 5028 44347
rect 9214 44344 9220 44356
rect 9272 44344 9278 44396
rect 18892 44393 18920 44424
rect 18877 44387 18935 44393
rect 18877 44353 18889 44387
rect 18923 44353 18935 44387
rect 18877 44347 18935 44353
rect 18969 44387 19027 44393
rect 18969 44353 18981 44387
rect 19015 44384 19027 44387
rect 19058 44384 19064 44396
rect 19015 44356 19064 44384
rect 19015 44353 19027 44356
rect 18969 44347 19027 44353
rect 19058 44344 19064 44356
rect 19116 44344 19122 44396
rect 19245 44387 19303 44393
rect 19245 44384 19257 44387
rect 19168 44356 19257 44384
rect 19168 44328 19196 44356
rect 19245 44353 19257 44356
rect 19291 44353 19303 44387
rect 19245 44347 19303 44353
rect 9950 44316 9956 44328
rect 5000 44288 9956 44316
rect 9950 44276 9956 44288
rect 10008 44276 10014 44328
rect 19150 44276 19156 44328
rect 19208 44276 19214 44328
rect 9490 44248 9496 44260
rect 4724 44220 9496 44248
rect 9490 44208 9496 44220
rect 9548 44208 9554 44260
rect 10226 44208 10232 44260
rect 10284 44208 10290 44260
rect 22066 44248 22094 44424
rect 26878 44412 26884 44464
rect 26936 44452 26942 44464
rect 33594 44452 33600 44464
rect 26936 44424 33600 44452
rect 26936 44412 26942 44424
rect 33594 44412 33600 44424
rect 33652 44452 33658 44464
rect 33652 44424 38148 44452
rect 33652 44412 33658 44424
rect 38120 44393 38148 44424
rect 37461 44387 37519 44393
rect 37461 44353 37473 44387
rect 37507 44353 37519 44387
rect 37461 44347 37519 44353
rect 38105 44387 38163 44393
rect 38105 44353 38117 44387
rect 38151 44353 38163 44387
rect 38105 44347 38163 44353
rect 34974 44276 34980 44328
rect 35032 44316 35038 44328
rect 35434 44316 35440 44328
rect 35032 44288 35440 44316
rect 35032 44276 35038 44288
rect 35434 44276 35440 44288
rect 35492 44316 35498 44328
rect 37476 44316 37504 44347
rect 35492 44288 37504 44316
rect 35492 44276 35498 44288
rect 35894 44248 35900 44260
rect 22066 44220 35900 44248
rect 35894 44208 35900 44220
rect 35952 44248 35958 44260
rect 36446 44248 36452 44260
rect 35952 44220 36452 44248
rect 35952 44208 35958 44220
rect 36446 44208 36452 44220
rect 36504 44208 36510 44260
rect 4890 44140 4896 44192
rect 4948 44180 4954 44192
rect 5074 44180 5080 44192
rect 4948 44152 5080 44180
rect 4948 44140 4954 44152
rect 5074 44140 5080 44152
rect 5132 44140 5138 44192
rect 9030 44140 9036 44192
rect 9088 44180 9094 44192
rect 9306 44180 9312 44192
rect 9088 44152 9312 44180
rect 9088 44140 9094 44152
rect 9306 44140 9312 44152
rect 9364 44140 9370 44192
rect 9950 44140 9956 44192
rect 10008 44180 10014 44192
rect 14274 44180 14280 44192
rect 10008 44152 14280 44180
rect 10008 44140 10014 44152
rect 14274 44140 14280 44152
rect 14332 44140 14338 44192
rect 33686 44140 33692 44192
rect 33744 44180 33750 44192
rect 37553 44183 37611 44189
rect 37553 44180 37565 44183
rect 33744 44152 37565 44180
rect 33744 44140 33750 44152
rect 37553 44149 37565 44152
rect 37599 44149 37611 44183
rect 37553 44143 37611 44149
rect 1104 44090 40848 44112
rect 1104 44038 1950 44090
rect 2002 44038 2014 44090
rect 2066 44038 2078 44090
rect 2130 44038 2142 44090
rect 2194 44038 2206 44090
rect 2258 44038 6950 44090
rect 7002 44038 7014 44090
rect 7066 44038 7078 44090
rect 7130 44038 7142 44090
rect 7194 44038 7206 44090
rect 7258 44038 11950 44090
rect 12002 44038 12014 44090
rect 12066 44038 12078 44090
rect 12130 44038 12142 44090
rect 12194 44038 12206 44090
rect 12258 44038 16950 44090
rect 17002 44038 17014 44090
rect 17066 44038 17078 44090
rect 17130 44038 17142 44090
rect 17194 44038 17206 44090
rect 17258 44038 21950 44090
rect 22002 44038 22014 44090
rect 22066 44038 22078 44090
rect 22130 44038 22142 44090
rect 22194 44038 22206 44090
rect 22258 44038 26950 44090
rect 27002 44038 27014 44090
rect 27066 44038 27078 44090
rect 27130 44038 27142 44090
rect 27194 44038 27206 44090
rect 27258 44038 31950 44090
rect 32002 44038 32014 44090
rect 32066 44038 32078 44090
rect 32130 44038 32142 44090
rect 32194 44038 32206 44090
rect 32258 44038 36950 44090
rect 37002 44038 37014 44090
rect 37066 44038 37078 44090
rect 37130 44038 37142 44090
rect 37194 44038 37206 44090
rect 37258 44038 40848 44090
rect 1104 44016 40848 44038
rect 19610 43936 19616 43988
rect 19668 43976 19674 43988
rect 32490 43976 32496 43988
rect 19668 43948 32496 43976
rect 19668 43936 19674 43948
rect 32490 43936 32496 43948
rect 32548 43936 32554 43988
rect 25958 43596 25964 43648
rect 26016 43636 26022 43648
rect 36630 43636 36636 43648
rect 26016 43608 36636 43636
rect 26016 43596 26022 43608
rect 36630 43596 36636 43608
rect 36688 43596 36694 43648
rect 1104 43546 40848 43568
rect 1104 43494 2610 43546
rect 2662 43494 2674 43546
rect 2726 43494 2738 43546
rect 2790 43494 2802 43546
rect 2854 43494 2866 43546
rect 2918 43494 7610 43546
rect 7662 43494 7674 43546
rect 7726 43494 7738 43546
rect 7790 43494 7802 43546
rect 7854 43494 7866 43546
rect 7918 43494 12610 43546
rect 12662 43494 12674 43546
rect 12726 43494 12738 43546
rect 12790 43494 12802 43546
rect 12854 43494 12866 43546
rect 12918 43494 17610 43546
rect 17662 43494 17674 43546
rect 17726 43494 17738 43546
rect 17790 43494 17802 43546
rect 17854 43494 17866 43546
rect 17918 43494 22610 43546
rect 22662 43494 22674 43546
rect 22726 43494 22738 43546
rect 22790 43494 22802 43546
rect 22854 43494 22866 43546
rect 22918 43494 27610 43546
rect 27662 43494 27674 43546
rect 27726 43494 27738 43546
rect 27790 43494 27802 43546
rect 27854 43494 27866 43546
rect 27918 43494 32610 43546
rect 32662 43494 32674 43546
rect 32726 43494 32738 43546
rect 32790 43494 32802 43546
rect 32854 43494 32866 43546
rect 32918 43494 37610 43546
rect 37662 43494 37674 43546
rect 37726 43494 37738 43546
rect 37790 43494 37802 43546
rect 37854 43494 37866 43546
rect 37918 43494 40848 43546
rect 1104 43472 40848 43494
rect 10870 43392 10876 43444
rect 10928 43432 10934 43444
rect 10928 43404 11744 43432
rect 10928 43392 10934 43404
rect 5074 43324 5080 43376
rect 5132 43364 5138 43376
rect 11716 43364 11744 43404
rect 14182 43392 14188 43444
rect 14240 43432 14246 43444
rect 33042 43432 33048 43444
rect 14240 43404 33048 43432
rect 14240 43392 14246 43404
rect 33042 43392 33048 43404
rect 33100 43392 33106 43444
rect 5132 43336 11652 43364
rect 5132 43324 5138 43336
rect 9582 43256 9588 43308
rect 9640 43256 9646 43308
rect 9674 43256 9680 43308
rect 9732 43296 9738 43308
rect 10042 43296 10048 43308
rect 9732 43268 10048 43296
rect 9732 43256 9738 43268
rect 10042 43256 10048 43268
rect 10100 43256 10106 43308
rect 11624 43305 11652 43336
rect 11716 43336 16574 43364
rect 11716 43305 11744 43336
rect 11609 43299 11667 43305
rect 11609 43265 11621 43299
rect 11655 43265 11667 43299
rect 11609 43259 11667 43265
rect 11701 43299 11759 43305
rect 11701 43265 11713 43299
rect 11747 43265 11759 43299
rect 11701 43259 11759 43265
rect 12069 43299 12127 43305
rect 12069 43265 12081 43299
rect 12115 43265 12127 43299
rect 16546 43296 16574 43336
rect 27982 43296 27988 43308
rect 16546 43268 27988 43296
rect 12069 43259 12127 43265
rect 9769 43231 9827 43237
rect 9769 43197 9781 43231
rect 9815 43197 9827 43231
rect 9769 43191 9827 43197
rect 9861 43231 9919 43237
rect 9861 43197 9873 43231
rect 9907 43228 9919 43231
rect 10502 43228 10508 43240
rect 9907 43200 10508 43228
rect 9907 43197 9919 43200
rect 9861 43191 9919 43197
rect 9398 43052 9404 43104
rect 9456 43052 9462 43104
rect 9784 43092 9812 43191
rect 10502 43188 10508 43200
rect 10560 43188 10566 43240
rect 11238 43188 11244 43240
rect 11296 43228 11302 43240
rect 11422 43228 11428 43240
rect 11296 43200 11428 43228
rect 11296 43188 11302 43200
rect 11422 43188 11428 43200
rect 11480 43228 11486 43240
rect 12084 43228 12112 43259
rect 27982 43256 27988 43268
rect 28040 43256 28046 43308
rect 11480 43200 12112 43228
rect 11480 43188 11486 43200
rect 16574 43188 16580 43240
rect 16632 43228 16638 43240
rect 16758 43228 16764 43240
rect 16632 43200 16764 43228
rect 16632 43188 16638 43200
rect 16758 43188 16764 43200
rect 16816 43188 16822 43240
rect 12253 43163 12311 43169
rect 12253 43129 12265 43163
rect 12299 43160 12311 43163
rect 12342 43160 12348 43172
rect 12299 43132 12348 43160
rect 12299 43129 12311 43132
rect 12253 43123 12311 43129
rect 12342 43120 12348 43132
rect 12400 43120 12406 43172
rect 16758 43092 16764 43104
rect 9784 43064 16764 43092
rect 16758 43052 16764 43064
rect 16816 43092 16822 43104
rect 19610 43092 19616 43104
rect 16816 43064 19616 43092
rect 16816 43052 16822 43064
rect 19610 43052 19616 43064
rect 19668 43052 19674 43104
rect 1104 43002 40848 43024
rect 1104 42950 1950 43002
rect 2002 42950 2014 43002
rect 2066 42950 2078 43002
rect 2130 42950 2142 43002
rect 2194 42950 2206 43002
rect 2258 42950 6950 43002
rect 7002 42950 7014 43002
rect 7066 42950 7078 43002
rect 7130 42950 7142 43002
rect 7194 42950 7206 43002
rect 7258 42950 11950 43002
rect 12002 42950 12014 43002
rect 12066 42950 12078 43002
rect 12130 42950 12142 43002
rect 12194 42950 12206 43002
rect 12258 42950 16950 43002
rect 17002 42950 17014 43002
rect 17066 42950 17078 43002
rect 17130 42950 17142 43002
rect 17194 42950 17206 43002
rect 17258 42950 21950 43002
rect 22002 42950 22014 43002
rect 22066 42950 22078 43002
rect 22130 42950 22142 43002
rect 22194 42950 22206 43002
rect 22258 42950 26950 43002
rect 27002 42950 27014 43002
rect 27066 42950 27078 43002
rect 27130 42950 27142 43002
rect 27194 42950 27206 43002
rect 27258 42950 31950 43002
rect 32002 42950 32014 43002
rect 32066 42950 32078 43002
rect 32130 42950 32142 43002
rect 32194 42950 32206 43002
rect 32258 42950 36950 43002
rect 37002 42950 37014 43002
rect 37066 42950 37078 43002
rect 37130 42950 37142 43002
rect 37194 42950 37206 43002
rect 37258 42950 40848 43002
rect 1104 42928 40848 42950
rect 22186 42848 22192 42900
rect 22244 42888 22250 42900
rect 23198 42888 23204 42900
rect 22244 42860 23204 42888
rect 22244 42848 22250 42860
rect 23198 42848 23204 42860
rect 23256 42848 23262 42900
rect 21542 42780 21548 42832
rect 21600 42780 21606 42832
rect 22204 42792 22876 42820
rect 3050 42712 3056 42764
rect 3108 42752 3114 42764
rect 8386 42752 8392 42764
rect 3108 42724 8392 42752
rect 3108 42712 3114 42724
rect 8386 42712 8392 42724
rect 8444 42712 8450 42764
rect 19518 42712 19524 42764
rect 19576 42752 19582 42764
rect 22204 42752 22232 42792
rect 19576 42724 22232 42752
rect 19576 42712 19582 42724
rect 12986 42644 12992 42696
rect 13044 42684 13050 42696
rect 20732 42693 20760 42724
rect 22278 42712 22284 42764
rect 22336 42752 22342 42764
rect 22738 42752 22744 42764
rect 22336 42724 22744 42752
rect 22336 42712 22342 42724
rect 22738 42712 22744 42724
rect 22796 42712 22802 42764
rect 22848 42752 22876 42792
rect 23934 42752 23940 42764
rect 22848 42724 23940 42752
rect 23934 42712 23940 42724
rect 23992 42712 23998 42764
rect 20349 42687 20407 42693
rect 20349 42684 20361 42687
rect 13044 42656 20361 42684
rect 13044 42644 13050 42656
rect 20349 42653 20361 42656
rect 20395 42653 20407 42687
rect 20349 42647 20407 42653
rect 20625 42687 20683 42693
rect 20625 42653 20637 42687
rect 20671 42653 20683 42687
rect 20625 42647 20683 42653
rect 20717 42687 20775 42693
rect 20717 42653 20729 42687
rect 20763 42653 20775 42687
rect 20717 42647 20775 42653
rect 18598 42576 18604 42628
rect 18656 42616 18662 42628
rect 19150 42616 19156 42628
rect 18656 42588 19156 42616
rect 18656 42576 18662 42588
rect 19150 42576 19156 42588
rect 19208 42616 19214 42628
rect 20640 42616 20668 42647
rect 22094 42644 22100 42696
rect 22152 42684 22158 42696
rect 22465 42687 22523 42693
rect 22465 42684 22477 42687
rect 22152 42656 22477 42684
rect 22152 42644 22158 42656
rect 22465 42653 22477 42656
rect 22511 42653 22523 42687
rect 23017 42687 23075 42693
rect 23017 42684 23029 42687
rect 22465 42647 22523 42653
rect 22572 42656 23029 42684
rect 19208 42588 20668 42616
rect 21085 42619 21143 42625
rect 19208 42576 19214 42588
rect 21085 42585 21097 42619
rect 21131 42616 21143 42619
rect 21174 42616 21180 42628
rect 21131 42588 21180 42616
rect 21131 42585 21143 42588
rect 21085 42579 21143 42585
rect 21174 42576 21180 42588
rect 21232 42576 21238 42628
rect 22572 42616 22600 42656
rect 23017 42653 23029 42656
rect 23063 42653 23075 42687
rect 23017 42647 23075 42653
rect 23382 42644 23388 42696
rect 23440 42644 23446 42696
rect 21284 42588 22600 42616
rect 22833 42619 22891 42625
rect 5166 42508 5172 42560
rect 5224 42548 5230 42560
rect 21284 42548 21312 42588
rect 22833 42585 22845 42619
rect 22879 42616 22891 42619
rect 23198 42616 23204 42628
rect 22879 42588 23204 42616
rect 22879 42585 22891 42588
rect 22833 42579 22891 42585
rect 23198 42576 23204 42588
rect 23256 42616 23262 42628
rect 23400 42616 23428 42644
rect 23256 42588 23428 42616
rect 23256 42576 23262 42588
rect 5224 42520 21312 42548
rect 5224 42508 5230 42520
rect 22370 42508 22376 42560
rect 22428 42548 22434 42560
rect 22649 42551 22707 42557
rect 22649 42548 22661 42551
rect 22428 42520 22661 42548
rect 22428 42508 22434 42520
rect 22649 42517 22661 42520
rect 22695 42517 22707 42551
rect 22649 42511 22707 42517
rect 22738 42508 22744 42560
rect 22796 42548 22802 42560
rect 23382 42548 23388 42560
rect 22796 42520 23388 42548
rect 22796 42508 22802 42520
rect 23382 42508 23388 42520
rect 23440 42508 23446 42560
rect 1104 42458 40848 42480
rect 1104 42406 2610 42458
rect 2662 42406 2674 42458
rect 2726 42406 2738 42458
rect 2790 42406 2802 42458
rect 2854 42406 2866 42458
rect 2918 42406 7610 42458
rect 7662 42406 7674 42458
rect 7726 42406 7738 42458
rect 7790 42406 7802 42458
rect 7854 42406 7866 42458
rect 7918 42406 12610 42458
rect 12662 42406 12674 42458
rect 12726 42406 12738 42458
rect 12790 42406 12802 42458
rect 12854 42406 12866 42458
rect 12918 42406 17610 42458
rect 17662 42406 17674 42458
rect 17726 42406 17738 42458
rect 17790 42406 17802 42458
rect 17854 42406 17866 42458
rect 17918 42406 22610 42458
rect 22662 42406 22674 42458
rect 22726 42406 22738 42458
rect 22790 42406 22802 42458
rect 22854 42406 22866 42458
rect 22918 42406 27610 42458
rect 27662 42406 27674 42458
rect 27726 42406 27738 42458
rect 27790 42406 27802 42458
rect 27854 42406 27866 42458
rect 27918 42406 32610 42458
rect 32662 42406 32674 42458
rect 32726 42406 32738 42458
rect 32790 42406 32802 42458
rect 32854 42406 32866 42458
rect 32918 42406 37610 42458
rect 37662 42406 37674 42458
rect 37726 42406 37738 42458
rect 37790 42406 37802 42458
rect 37854 42406 37866 42458
rect 37918 42406 40848 42458
rect 1104 42384 40848 42406
rect 13998 42304 14004 42356
rect 14056 42344 14062 42356
rect 25682 42344 25688 42356
rect 14056 42316 25688 42344
rect 14056 42304 14062 42316
rect 25682 42304 25688 42316
rect 25740 42304 25746 42356
rect 18506 42236 18512 42288
rect 18564 42276 18570 42288
rect 24670 42276 24676 42288
rect 18564 42248 23060 42276
rect 18564 42236 18570 42248
rect 19886 42168 19892 42220
rect 19944 42208 19950 42220
rect 22370 42208 22376 42220
rect 19944 42180 22376 42208
rect 19944 42168 19950 42180
rect 22370 42168 22376 42180
rect 22428 42168 22434 42220
rect 5534 42032 5540 42084
rect 5592 42072 5598 42084
rect 6086 42072 6092 42084
rect 5592 42044 6092 42072
rect 5592 42032 5598 42044
rect 6086 42032 6092 42044
rect 6144 42072 6150 42084
rect 18598 42072 18604 42084
rect 6144 42044 18604 42072
rect 6144 42032 6150 42044
rect 18598 42032 18604 42044
rect 18656 42032 18662 42084
rect 23032 42013 23060 42248
rect 23952 42248 24676 42276
rect 23566 42168 23572 42220
rect 23624 42168 23630 42220
rect 23658 42168 23664 42220
rect 23716 42168 23722 42220
rect 23952 42217 23980 42248
rect 24670 42236 24676 42248
rect 24728 42236 24734 42288
rect 27982 42236 27988 42288
rect 28040 42276 28046 42288
rect 28040 42248 35894 42276
rect 28040 42236 28046 42248
rect 23937 42211 23995 42217
rect 23937 42177 23949 42211
rect 23983 42177 23995 42211
rect 23937 42171 23995 42177
rect 24026 42168 24032 42220
rect 24084 42208 24090 42220
rect 24121 42211 24179 42217
rect 24121 42208 24133 42211
rect 24084 42180 24133 42208
rect 24084 42168 24090 42180
rect 24121 42177 24133 42180
rect 24167 42208 24179 42211
rect 24302 42208 24308 42220
rect 24167 42180 24308 42208
rect 24167 42177 24179 42180
rect 24121 42171 24179 42177
rect 24302 42168 24308 42180
rect 24360 42168 24366 42220
rect 26326 42168 26332 42220
rect 26384 42208 26390 42220
rect 26786 42208 26792 42220
rect 26384 42180 26792 42208
rect 26384 42168 26390 42180
rect 26786 42168 26792 42180
rect 26844 42208 26850 42220
rect 26973 42211 27031 42217
rect 26973 42208 26985 42211
rect 26844 42180 26985 42208
rect 26844 42168 26850 42180
rect 26973 42177 26985 42180
rect 27019 42177 27031 42211
rect 26973 42171 27031 42177
rect 27338 42168 27344 42220
rect 27396 42208 27402 42220
rect 32125 42211 32183 42217
rect 32125 42208 32137 42211
rect 27396 42180 32137 42208
rect 27396 42168 27402 42180
rect 32125 42177 32137 42180
rect 32171 42177 32183 42211
rect 32125 42171 32183 42177
rect 32232 42180 33180 42208
rect 26050 42100 26056 42152
rect 26108 42140 26114 42152
rect 27433 42143 27491 42149
rect 27433 42140 27445 42143
rect 26108 42112 27445 42140
rect 26108 42100 26114 42112
rect 27433 42109 27445 42112
rect 27479 42109 27491 42143
rect 27433 42103 27491 42109
rect 29546 42100 29552 42152
rect 29604 42140 29610 42152
rect 32232 42140 32260 42180
rect 29604 42112 32260 42140
rect 29604 42100 29610 42112
rect 32858 42100 32864 42152
rect 32916 42100 32922 42152
rect 33152 42140 33180 42180
rect 33226 42168 33232 42220
rect 33284 42208 33290 42220
rect 33689 42211 33747 42217
rect 33689 42208 33701 42211
rect 33284 42180 33701 42208
rect 33284 42168 33290 42180
rect 33689 42177 33701 42180
rect 33735 42177 33747 42211
rect 33689 42171 33747 42177
rect 33965 42143 34023 42149
rect 33965 42140 33977 42143
rect 33152 42112 33977 42140
rect 33965 42109 33977 42112
rect 34011 42109 34023 42143
rect 35866 42140 35894 42248
rect 36078 42140 36084 42152
rect 35866 42112 36084 42140
rect 33965 42103 34023 42109
rect 36078 42100 36084 42112
rect 36136 42100 36142 42152
rect 23934 42032 23940 42084
rect 23992 42072 23998 42084
rect 35986 42072 35992 42084
rect 23992 42044 35992 42072
rect 23992 42032 23998 42044
rect 35986 42032 35992 42044
rect 36044 42032 36050 42084
rect 23017 42007 23075 42013
rect 23017 41973 23029 42007
rect 23063 42004 23075 42007
rect 26418 42004 26424 42016
rect 23063 41976 26424 42004
rect 23063 41973 23075 41976
rect 23017 41967 23075 41973
rect 26418 41964 26424 41976
rect 26476 41964 26482 42016
rect 1104 41914 40848 41936
rect 1104 41862 1950 41914
rect 2002 41862 2014 41914
rect 2066 41862 2078 41914
rect 2130 41862 2142 41914
rect 2194 41862 2206 41914
rect 2258 41862 6950 41914
rect 7002 41862 7014 41914
rect 7066 41862 7078 41914
rect 7130 41862 7142 41914
rect 7194 41862 7206 41914
rect 7258 41862 11950 41914
rect 12002 41862 12014 41914
rect 12066 41862 12078 41914
rect 12130 41862 12142 41914
rect 12194 41862 12206 41914
rect 12258 41862 16950 41914
rect 17002 41862 17014 41914
rect 17066 41862 17078 41914
rect 17130 41862 17142 41914
rect 17194 41862 17206 41914
rect 17258 41862 21950 41914
rect 22002 41862 22014 41914
rect 22066 41862 22078 41914
rect 22130 41862 22142 41914
rect 22194 41862 22206 41914
rect 22258 41862 26950 41914
rect 27002 41862 27014 41914
rect 27066 41862 27078 41914
rect 27130 41862 27142 41914
rect 27194 41862 27206 41914
rect 27258 41862 31950 41914
rect 32002 41862 32014 41914
rect 32066 41862 32078 41914
rect 32130 41862 32142 41914
rect 32194 41862 32206 41914
rect 32258 41862 36950 41914
rect 37002 41862 37014 41914
rect 37066 41862 37078 41914
rect 37130 41862 37142 41914
rect 37194 41862 37206 41914
rect 37258 41862 40848 41914
rect 1104 41840 40848 41862
rect 9122 41760 9128 41812
rect 9180 41800 9186 41812
rect 9490 41800 9496 41812
rect 9180 41772 9496 41800
rect 9180 41760 9186 41772
rect 9490 41760 9496 41772
rect 9548 41760 9554 41812
rect 27338 41800 27344 41812
rect 16546 41772 27344 41800
rect 8938 41692 8944 41744
rect 8996 41732 9002 41744
rect 16546 41732 16574 41772
rect 27338 41760 27344 41772
rect 27396 41760 27402 41812
rect 8996 41704 16574 41732
rect 8996 41692 9002 41704
rect 29730 41624 29736 41676
rect 29788 41664 29794 41676
rect 29788 41636 33088 41664
rect 29788 41624 29794 41636
rect 15562 41556 15568 41608
rect 15620 41596 15626 41608
rect 16482 41596 16488 41608
rect 15620 41568 16488 41596
rect 15620 41556 15626 41568
rect 16482 41556 16488 41568
rect 16540 41596 16546 41608
rect 32677 41599 32735 41605
rect 32677 41596 32689 41599
rect 16540 41568 32689 41596
rect 16540 41556 16546 41568
rect 32677 41565 32689 41568
rect 32723 41596 32735 41599
rect 32766 41596 32772 41608
rect 32723 41568 32772 41596
rect 32723 41565 32735 41568
rect 32677 41559 32735 41565
rect 32766 41556 32772 41568
rect 32824 41556 32830 41608
rect 33060 41605 33088 41636
rect 33226 41624 33232 41676
rect 33284 41624 33290 41676
rect 33045 41599 33103 41605
rect 33045 41565 33057 41599
rect 33091 41565 33103 41599
rect 33045 41559 33103 41565
rect 33781 41599 33839 41605
rect 33781 41565 33793 41599
rect 33827 41596 33839 41599
rect 34974 41596 34980 41608
rect 33827 41568 34980 41596
rect 33827 41565 33839 41568
rect 33781 41559 33839 41565
rect 34974 41556 34980 41568
rect 35032 41556 35038 41608
rect 8478 41488 8484 41540
rect 8536 41528 8542 41540
rect 8938 41528 8944 41540
rect 8536 41500 8944 41528
rect 8536 41488 8542 41500
rect 8938 41488 8944 41500
rect 8996 41488 9002 41540
rect 28258 41488 28264 41540
rect 28316 41528 28322 41540
rect 32306 41528 32312 41540
rect 28316 41500 32312 41528
rect 28316 41488 28322 41500
rect 32306 41488 32312 41500
rect 32364 41488 32370 41540
rect 8754 41420 8760 41472
rect 8812 41460 8818 41472
rect 11790 41460 11796 41472
rect 8812 41432 11796 41460
rect 8812 41420 8818 41432
rect 11790 41420 11796 41432
rect 11848 41420 11854 41472
rect 23106 41420 23112 41472
rect 23164 41460 23170 41472
rect 23750 41460 23756 41472
rect 23164 41432 23756 41460
rect 23164 41420 23170 41432
rect 23750 41420 23756 41432
rect 23808 41420 23814 41472
rect 28350 41420 28356 41472
rect 28408 41460 28414 41472
rect 28810 41460 28816 41472
rect 28408 41432 28816 41460
rect 28408 41420 28414 41432
rect 28810 41420 28816 41432
rect 28868 41420 28874 41472
rect 31110 41420 31116 41472
rect 31168 41460 31174 41472
rect 33318 41460 33324 41472
rect 31168 41432 33324 41460
rect 31168 41420 31174 41432
rect 33318 41420 33324 41432
rect 33376 41420 33382 41472
rect 36630 41420 36636 41472
rect 36688 41460 36694 41472
rect 38654 41460 38660 41472
rect 36688 41432 38660 41460
rect 36688 41420 36694 41432
rect 38654 41420 38660 41432
rect 38712 41420 38718 41472
rect 1104 41370 40848 41392
rect 1104 41318 2610 41370
rect 2662 41318 2674 41370
rect 2726 41318 2738 41370
rect 2790 41318 2802 41370
rect 2854 41318 2866 41370
rect 2918 41318 7610 41370
rect 7662 41318 7674 41370
rect 7726 41318 7738 41370
rect 7790 41318 7802 41370
rect 7854 41318 7866 41370
rect 7918 41318 12610 41370
rect 12662 41318 12674 41370
rect 12726 41318 12738 41370
rect 12790 41318 12802 41370
rect 12854 41318 12866 41370
rect 12918 41318 17610 41370
rect 17662 41318 17674 41370
rect 17726 41318 17738 41370
rect 17790 41318 17802 41370
rect 17854 41318 17866 41370
rect 17918 41318 22610 41370
rect 22662 41318 22674 41370
rect 22726 41318 22738 41370
rect 22790 41318 22802 41370
rect 22854 41318 22866 41370
rect 22918 41318 27610 41370
rect 27662 41318 27674 41370
rect 27726 41318 27738 41370
rect 27790 41318 27802 41370
rect 27854 41318 27866 41370
rect 27918 41318 32610 41370
rect 32662 41318 32674 41370
rect 32726 41318 32738 41370
rect 32790 41318 32802 41370
rect 32854 41318 32866 41370
rect 32918 41318 37610 41370
rect 37662 41318 37674 41370
rect 37726 41318 37738 41370
rect 37790 41318 37802 41370
rect 37854 41318 37866 41370
rect 37918 41318 40848 41370
rect 1104 41296 40848 41318
rect 16574 41216 16580 41268
rect 16632 41256 16638 41268
rect 17310 41256 17316 41268
rect 16632 41228 17316 41256
rect 16632 41216 16638 41228
rect 17310 41216 17316 41228
rect 17368 41216 17374 41268
rect 19978 41216 19984 41268
rect 20036 41256 20042 41268
rect 20036 41228 29592 41256
rect 20036 41216 20042 41228
rect 21542 41188 21548 41200
rect 8036 41160 21548 41188
rect 2777 41123 2835 41129
rect 2777 41089 2789 41123
rect 2823 41120 2835 41123
rect 5534 41120 5540 41132
rect 2823 41092 5540 41120
rect 2823 41089 2835 41092
rect 2777 41083 2835 41089
rect 5534 41080 5540 41092
rect 5592 41080 5598 41132
rect 8036 41129 8064 41160
rect 21542 41148 21548 41160
rect 21600 41148 21606 41200
rect 29178 41188 29184 41200
rect 22066 41160 29184 41188
rect 8021 41123 8079 41129
rect 8021 41089 8033 41123
rect 8067 41089 8079 41123
rect 8021 41083 8079 41089
rect 8389 41123 8447 41129
rect 8389 41089 8401 41123
rect 8435 41120 8447 41123
rect 17310 41120 17316 41132
rect 8435 41092 17316 41120
rect 8435 41089 8447 41092
rect 8389 41083 8447 41089
rect 17310 41080 17316 41092
rect 17368 41080 17374 41132
rect 3418 41012 3424 41064
rect 3476 41052 3482 41064
rect 3878 41052 3884 41064
rect 3476 41024 3884 41052
rect 3476 41012 3482 41024
rect 3878 41012 3884 41024
rect 3936 41012 3942 41064
rect 8481 41055 8539 41061
rect 8481 41021 8493 41055
rect 8527 41052 8539 41055
rect 10410 41052 10416 41064
rect 8527 41024 10416 41052
rect 8527 41021 8539 41024
rect 8481 41015 8539 41021
rect 10410 41012 10416 41024
rect 10468 41012 10474 41064
rect 21560 41052 21588 41148
rect 22066 41052 22094 41160
rect 29178 41148 29184 41160
rect 29236 41148 29242 41200
rect 22830 41080 22836 41132
rect 22888 41120 22894 41132
rect 23382 41120 23388 41132
rect 22888 41092 23388 41120
rect 22888 41080 22894 41092
rect 23382 41080 23388 41092
rect 23440 41080 23446 41132
rect 25130 41080 25136 41132
rect 25188 41120 25194 41132
rect 25866 41120 25872 41132
rect 25188 41092 25872 41120
rect 25188 41080 25194 41092
rect 25866 41080 25872 41092
rect 25924 41080 25930 41132
rect 27982 41080 27988 41132
rect 28040 41120 28046 41132
rect 28537 41123 28595 41129
rect 28537 41120 28549 41123
rect 28040 41092 28549 41120
rect 28040 41080 28046 41092
rect 28537 41089 28549 41092
rect 28583 41089 28595 41123
rect 28537 41083 28595 41089
rect 29270 41080 29276 41132
rect 29328 41080 29334 41132
rect 29564 41129 29592 41228
rect 29638 41216 29644 41268
rect 29696 41256 29702 41268
rect 29914 41256 29920 41268
rect 29696 41228 29920 41256
rect 29696 41216 29702 41228
rect 29914 41216 29920 41228
rect 29972 41216 29978 41268
rect 34054 41188 34060 41200
rect 31726 41160 34060 41188
rect 29549 41123 29607 41129
rect 29549 41089 29561 41123
rect 29595 41089 29607 41123
rect 29549 41083 29607 41089
rect 29914 41080 29920 41132
rect 29972 41080 29978 41132
rect 30558 41080 30564 41132
rect 30616 41080 30622 41132
rect 30834 41080 30840 41132
rect 30892 41120 30898 41132
rect 30929 41123 30987 41129
rect 30929 41120 30941 41123
rect 30892 41092 30941 41120
rect 30892 41080 30898 41092
rect 30929 41089 30941 41092
rect 30975 41089 30987 41123
rect 30929 41083 30987 41089
rect 30101 41055 30159 41061
rect 30101 41052 30113 41055
rect 21560 41024 22094 41052
rect 23032 41024 30113 41052
rect 7837 40987 7895 40993
rect 7837 40953 7849 40987
rect 7883 40984 7895 40987
rect 22738 40984 22744 40996
rect 7883 40956 22744 40984
rect 7883 40953 7895 40956
rect 7837 40947 7895 40953
rect 22738 40944 22744 40956
rect 22796 40944 22802 40996
rect 10594 40876 10600 40928
rect 10652 40916 10658 40928
rect 23032 40916 23060 41024
rect 30101 41021 30113 41024
rect 30147 41021 30159 41055
rect 30101 41015 30159 41021
rect 31018 41012 31024 41064
rect 31076 41012 31082 41064
rect 23658 40944 23664 40996
rect 23716 40984 23722 40996
rect 28629 40987 28687 40993
rect 28629 40984 28641 40987
rect 23716 40956 28641 40984
rect 23716 40944 23722 40956
rect 28629 40953 28641 40956
rect 28675 40953 28687 40987
rect 28629 40947 28687 40953
rect 29270 40944 29276 40996
rect 29328 40984 29334 40996
rect 31726 40984 31754 41160
rect 34054 41148 34060 41160
rect 34112 41148 34118 41200
rect 29328 40956 31754 40984
rect 29328 40944 29334 40956
rect 10652 40888 23060 40916
rect 10652 40876 10658 40888
rect 23106 40876 23112 40928
rect 23164 40916 23170 40928
rect 25685 40919 25743 40925
rect 25685 40916 25697 40919
rect 23164 40888 25697 40916
rect 23164 40876 23170 40888
rect 25685 40885 25697 40888
rect 25731 40885 25743 40919
rect 25685 40879 25743 40885
rect 29178 40876 29184 40928
rect 29236 40916 29242 40928
rect 30098 40916 30104 40928
rect 29236 40888 30104 40916
rect 29236 40876 29242 40888
rect 30098 40876 30104 40888
rect 30156 40876 30162 40928
rect 1104 40826 40848 40848
rect 1104 40774 1950 40826
rect 2002 40774 2014 40826
rect 2066 40774 2078 40826
rect 2130 40774 2142 40826
rect 2194 40774 2206 40826
rect 2258 40774 6950 40826
rect 7002 40774 7014 40826
rect 7066 40774 7078 40826
rect 7130 40774 7142 40826
rect 7194 40774 7206 40826
rect 7258 40774 11950 40826
rect 12002 40774 12014 40826
rect 12066 40774 12078 40826
rect 12130 40774 12142 40826
rect 12194 40774 12206 40826
rect 12258 40774 16950 40826
rect 17002 40774 17014 40826
rect 17066 40774 17078 40826
rect 17130 40774 17142 40826
rect 17194 40774 17206 40826
rect 17258 40774 21950 40826
rect 22002 40774 22014 40826
rect 22066 40774 22078 40826
rect 22130 40774 22142 40826
rect 22194 40774 22206 40826
rect 22258 40774 26950 40826
rect 27002 40774 27014 40826
rect 27066 40774 27078 40826
rect 27130 40774 27142 40826
rect 27194 40774 27206 40826
rect 27258 40774 31950 40826
rect 32002 40774 32014 40826
rect 32066 40774 32078 40826
rect 32130 40774 32142 40826
rect 32194 40774 32206 40826
rect 32258 40774 36950 40826
rect 37002 40774 37014 40826
rect 37066 40774 37078 40826
rect 37130 40774 37142 40826
rect 37194 40774 37206 40826
rect 37258 40774 40848 40826
rect 1104 40752 40848 40774
rect 13262 40672 13268 40724
rect 13320 40712 13326 40724
rect 17129 40715 17187 40721
rect 17129 40712 17141 40715
rect 13320 40684 17141 40712
rect 13320 40672 13326 40684
rect 17129 40681 17141 40684
rect 17175 40681 17187 40715
rect 17129 40675 17187 40681
rect 21358 40672 21364 40724
rect 21416 40712 21422 40724
rect 22465 40715 22523 40721
rect 22465 40712 22477 40715
rect 21416 40684 22477 40712
rect 21416 40672 21422 40684
rect 22465 40681 22477 40684
rect 22511 40712 22523 40715
rect 23014 40712 23020 40724
rect 22511 40684 23020 40712
rect 22511 40681 22523 40684
rect 22465 40675 22523 40681
rect 23014 40672 23020 40684
rect 23072 40672 23078 40724
rect 10962 40604 10968 40656
rect 11020 40644 11026 40656
rect 11020 40616 31616 40644
rect 11020 40604 11026 40616
rect 17221 40579 17279 40585
rect 17221 40545 17233 40579
rect 17267 40576 17279 40579
rect 29362 40576 29368 40588
rect 17267 40548 29368 40576
rect 17267 40545 17279 40548
rect 17221 40539 17279 40545
rect 29362 40536 29368 40548
rect 29420 40536 29426 40588
rect 31588 40585 31616 40616
rect 31573 40579 31631 40585
rect 31573 40545 31585 40579
rect 31619 40545 31631 40579
rect 31573 40539 31631 40545
rect 36262 40536 36268 40588
rect 36320 40576 36326 40588
rect 39209 40579 39267 40585
rect 39209 40576 39221 40579
rect 36320 40548 39221 40576
rect 36320 40536 36326 40548
rect 39209 40545 39221 40548
rect 39255 40576 39267 40579
rect 39298 40576 39304 40588
rect 39255 40548 39304 40576
rect 39255 40545 39267 40548
rect 39209 40539 39267 40545
rect 39298 40536 39304 40548
rect 39356 40536 39362 40588
rect 1762 40468 1768 40520
rect 1820 40508 1826 40520
rect 2225 40511 2283 40517
rect 2225 40508 2237 40511
rect 1820 40480 2237 40508
rect 1820 40468 1826 40480
rect 2225 40477 2237 40480
rect 2271 40477 2283 40511
rect 2225 40471 2283 40477
rect 2869 40511 2927 40517
rect 2869 40477 2881 40511
rect 2915 40508 2927 40511
rect 2958 40508 2964 40520
rect 2915 40480 2964 40508
rect 2915 40477 2927 40480
rect 2869 40471 2927 40477
rect 2958 40468 2964 40480
rect 3016 40468 3022 40520
rect 3510 40468 3516 40520
rect 3568 40468 3574 40520
rect 16758 40468 16764 40520
rect 16816 40508 16822 40520
rect 16945 40511 17003 40517
rect 16945 40508 16957 40511
rect 16816 40480 16957 40508
rect 16816 40468 16822 40480
rect 16945 40477 16957 40480
rect 16991 40477 17003 40511
rect 16945 40471 17003 40477
rect 22281 40511 22339 40517
rect 22281 40477 22293 40511
rect 22327 40508 22339 40511
rect 22462 40508 22468 40520
rect 22327 40480 22468 40508
rect 22327 40477 22339 40480
rect 22281 40471 22339 40477
rect 22462 40468 22468 40480
rect 22520 40468 22526 40520
rect 23106 40468 23112 40520
rect 23164 40468 23170 40520
rect 23566 40468 23572 40520
rect 23624 40508 23630 40520
rect 24670 40508 24676 40520
rect 23624 40480 24676 40508
rect 23624 40468 23630 40480
rect 24670 40468 24676 40480
rect 24728 40468 24734 40520
rect 25130 40468 25136 40520
rect 25188 40468 25194 40520
rect 31846 40468 31852 40520
rect 31904 40508 31910 40520
rect 32033 40511 32091 40517
rect 32033 40508 32045 40511
rect 31904 40480 32045 40508
rect 31904 40468 31910 40480
rect 32033 40477 32045 40480
rect 32079 40477 32091 40511
rect 32033 40471 32091 40477
rect 32125 40511 32183 40517
rect 32125 40477 32137 40511
rect 32171 40508 32183 40511
rect 32398 40508 32404 40520
rect 32171 40480 32404 40508
rect 32171 40477 32183 40480
rect 32125 40471 32183 40477
rect 32398 40468 32404 40480
rect 32456 40468 32462 40520
rect 3050 40400 3056 40452
rect 3108 40400 3114 40452
rect 24394 40400 24400 40452
rect 24452 40440 24458 40452
rect 24581 40443 24639 40449
rect 24581 40440 24593 40443
rect 24452 40412 24593 40440
rect 24452 40400 24458 40412
rect 24581 40409 24593 40412
rect 24627 40409 24639 40443
rect 24581 40403 24639 40409
rect 13538 40332 13544 40384
rect 13596 40372 13602 40384
rect 16761 40375 16819 40381
rect 16761 40372 16773 40375
rect 13596 40344 16773 40372
rect 13596 40332 13602 40344
rect 16761 40341 16773 40344
rect 16807 40341 16819 40375
rect 16761 40335 16819 40341
rect 22738 40332 22744 40384
rect 22796 40372 22802 40384
rect 29454 40372 29460 40384
rect 22796 40344 29460 40372
rect 22796 40332 22802 40344
rect 29454 40332 29460 40344
rect 29512 40332 29518 40384
rect 38654 40332 38660 40384
rect 38712 40332 38718 40384
rect 1104 40282 40848 40304
rect 1104 40230 2610 40282
rect 2662 40230 2674 40282
rect 2726 40230 2738 40282
rect 2790 40230 2802 40282
rect 2854 40230 2866 40282
rect 2918 40230 7610 40282
rect 7662 40230 7674 40282
rect 7726 40230 7738 40282
rect 7790 40230 7802 40282
rect 7854 40230 7866 40282
rect 7918 40230 12610 40282
rect 12662 40230 12674 40282
rect 12726 40230 12738 40282
rect 12790 40230 12802 40282
rect 12854 40230 12866 40282
rect 12918 40230 17610 40282
rect 17662 40230 17674 40282
rect 17726 40230 17738 40282
rect 17790 40230 17802 40282
rect 17854 40230 17866 40282
rect 17918 40230 22610 40282
rect 22662 40230 22674 40282
rect 22726 40230 22738 40282
rect 22790 40230 22802 40282
rect 22854 40230 22866 40282
rect 22918 40230 27610 40282
rect 27662 40230 27674 40282
rect 27726 40230 27738 40282
rect 27790 40230 27802 40282
rect 27854 40230 27866 40282
rect 27918 40230 32610 40282
rect 32662 40230 32674 40282
rect 32726 40230 32738 40282
rect 32790 40230 32802 40282
rect 32854 40230 32866 40282
rect 32918 40230 37610 40282
rect 37662 40230 37674 40282
rect 37726 40230 37738 40282
rect 37790 40230 37802 40282
rect 37854 40230 37866 40282
rect 37918 40230 40848 40282
rect 1104 40208 40848 40230
rect 16482 40128 16488 40180
rect 16540 40168 16546 40180
rect 16758 40168 16764 40180
rect 16540 40140 16764 40168
rect 16540 40128 16546 40140
rect 16758 40128 16764 40140
rect 16816 40128 16822 40180
rect 842 40060 848 40112
rect 900 40100 906 40112
rect 1397 40103 1455 40109
rect 1397 40100 1409 40103
rect 900 40072 1409 40100
rect 900 40060 906 40072
rect 1397 40069 1409 40072
rect 1443 40069 1455 40103
rect 1397 40063 1455 40069
rect 10594 40060 10600 40112
rect 10652 40100 10658 40112
rect 10870 40100 10876 40112
rect 10652 40072 10876 40100
rect 10652 40060 10658 40072
rect 10870 40060 10876 40072
rect 10928 40060 10934 40112
rect 17310 40060 17316 40112
rect 17368 40100 17374 40112
rect 24854 40100 24860 40112
rect 17368 40072 24860 40100
rect 17368 40060 17374 40072
rect 24854 40060 24860 40072
rect 24912 40100 24918 40112
rect 24912 40072 26188 40100
rect 24912 40060 24918 40072
rect 26160 40032 26188 40072
rect 39298 40060 39304 40112
rect 39356 40060 39362 40112
rect 40862 40100 40868 40112
rect 40604 40072 40868 40100
rect 32306 40032 32312 40044
rect 26160 40004 32312 40032
rect 32306 39992 32312 40004
rect 32364 39992 32370 40044
rect 40497 40035 40555 40041
rect 40497 40001 40509 40035
rect 40543 40032 40555 40035
rect 40604 40032 40632 40072
rect 40862 40060 40868 40072
rect 40920 40060 40926 40112
rect 40543 40004 40632 40032
rect 40543 40001 40555 40004
rect 40497 39995 40555 40001
rect 2225 39967 2283 39973
rect 2225 39933 2237 39967
rect 2271 39964 2283 39967
rect 8294 39964 8300 39976
rect 2271 39936 8300 39964
rect 2271 39933 2283 39936
rect 2225 39927 2283 39933
rect 8294 39924 8300 39936
rect 8352 39924 8358 39976
rect 10410 39856 10416 39908
rect 10468 39896 10474 39908
rect 30558 39896 30564 39908
rect 10468 39868 30564 39896
rect 10468 39856 10474 39868
rect 30558 39856 30564 39868
rect 30616 39856 30622 39908
rect 2498 39788 2504 39840
rect 2556 39828 2562 39840
rect 13446 39828 13452 39840
rect 2556 39800 13452 39828
rect 2556 39788 2562 39800
rect 13446 39788 13452 39800
rect 13504 39788 13510 39840
rect 15010 39788 15016 39840
rect 15068 39828 15074 39840
rect 23382 39828 23388 39840
rect 15068 39800 23388 39828
rect 15068 39788 15074 39800
rect 23382 39788 23388 39800
rect 23440 39788 23446 39840
rect 23658 39788 23664 39840
rect 23716 39828 23722 39840
rect 36722 39828 36728 39840
rect 23716 39800 36728 39828
rect 23716 39788 23722 39800
rect 36722 39788 36728 39800
rect 36780 39788 36786 39840
rect 1104 39738 40848 39760
rect 1104 39686 1950 39738
rect 2002 39686 2014 39738
rect 2066 39686 2078 39738
rect 2130 39686 2142 39738
rect 2194 39686 2206 39738
rect 2258 39686 6950 39738
rect 7002 39686 7014 39738
rect 7066 39686 7078 39738
rect 7130 39686 7142 39738
rect 7194 39686 7206 39738
rect 7258 39686 11950 39738
rect 12002 39686 12014 39738
rect 12066 39686 12078 39738
rect 12130 39686 12142 39738
rect 12194 39686 12206 39738
rect 12258 39686 16950 39738
rect 17002 39686 17014 39738
rect 17066 39686 17078 39738
rect 17130 39686 17142 39738
rect 17194 39686 17206 39738
rect 17258 39686 21950 39738
rect 22002 39686 22014 39738
rect 22066 39686 22078 39738
rect 22130 39686 22142 39738
rect 22194 39686 22206 39738
rect 22258 39686 26950 39738
rect 27002 39686 27014 39738
rect 27066 39686 27078 39738
rect 27130 39686 27142 39738
rect 27194 39686 27206 39738
rect 27258 39686 31950 39738
rect 32002 39686 32014 39738
rect 32066 39686 32078 39738
rect 32130 39686 32142 39738
rect 32194 39686 32206 39738
rect 32258 39686 36950 39738
rect 37002 39686 37014 39738
rect 37066 39686 37078 39738
rect 37130 39686 37142 39738
rect 37194 39686 37206 39738
rect 37258 39686 40848 39738
rect 1104 39664 40848 39686
rect 12805 39627 12863 39633
rect 12805 39593 12817 39627
rect 12851 39624 12863 39627
rect 14550 39624 14556 39636
rect 12851 39596 14556 39624
rect 12851 39593 12863 39596
rect 12805 39587 12863 39593
rect 14550 39584 14556 39596
rect 14608 39584 14614 39636
rect 23566 39624 23572 39636
rect 22066 39596 23572 39624
rect 4246 39516 4252 39568
rect 4304 39556 4310 39568
rect 14918 39556 14924 39568
rect 4304 39528 14924 39556
rect 4304 39516 4310 39528
rect 14918 39516 14924 39528
rect 14976 39516 14982 39568
rect 16298 39448 16304 39500
rect 16356 39488 16362 39500
rect 22066 39488 22094 39596
rect 23566 39584 23572 39596
rect 23624 39584 23630 39636
rect 30469 39627 30527 39633
rect 30469 39593 30481 39627
rect 30515 39624 30527 39627
rect 30742 39624 30748 39636
rect 30515 39596 30748 39624
rect 30515 39593 30527 39596
rect 30469 39587 30527 39593
rect 30742 39584 30748 39596
rect 30800 39584 30806 39636
rect 23382 39516 23388 39568
rect 23440 39556 23446 39568
rect 23440 39528 26004 39556
rect 23440 39516 23446 39528
rect 16356 39460 22094 39488
rect 25976 39488 26004 39528
rect 26234 39516 26240 39568
rect 26292 39556 26298 39568
rect 28629 39559 28687 39565
rect 28629 39556 28641 39559
rect 26292 39528 28641 39556
rect 26292 39516 26298 39528
rect 28629 39525 28641 39528
rect 28675 39525 28687 39559
rect 28629 39519 28687 39525
rect 28718 39516 28724 39568
rect 28776 39556 28782 39568
rect 29730 39556 29736 39568
rect 28776 39528 29736 39556
rect 28776 39516 28782 39528
rect 29730 39516 29736 39528
rect 29788 39516 29794 39568
rect 33134 39516 33140 39568
rect 33192 39516 33198 39568
rect 31297 39491 31355 39497
rect 25976 39460 28948 39488
rect 16356 39448 16362 39460
rect 12989 39423 13047 39429
rect 12989 39389 13001 39423
rect 13035 39389 13047 39423
rect 12989 39383 13047 39389
rect 13081 39423 13139 39429
rect 13081 39389 13093 39423
rect 13127 39389 13139 39423
rect 13081 39383 13139 39389
rect 13004 39284 13032 39383
rect 13096 39352 13124 39383
rect 13262 39380 13268 39432
rect 13320 39380 13326 39432
rect 13357 39423 13415 39429
rect 13357 39389 13369 39423
rect 13403 39420 13415 39423
rect 19426 39420 19432 39432
rect 13403 39392 19432 39420
rect 13403 39389 13415 39392
rect 13357 39383 13415 39389
rect 19426 39380 19432 39392
rect 19484 39380 19490 39432
rect 19610 39380 19616 39432
rect 19668 39420 19674 39432
rect 19794 39420 19800 39432
rect 19668 39392 19800 39420
rect 19668 39380 19674 39392
rect 19794 39380 19800 39392
rect 19852 39420 19858 39432
rect 19852 39392 21588 39420
rect 19852 39380 19858 39392
rect 21450 39352 21456 39364
rect 13096 39324 21456 39352
rect 21450 39312 21456 39324
rect 21508 39312 21514 39364
rect 21560 39352 21588 39392
rect 23198 39380 23204 39432
rect 23256 39380 23262 39432
rect 23290 39380 23296 39432
rect 23348 39380 23354 39432
rect 23477 39423 23535 39429
rect 23477 39389 23489 39423
rect 23523 39420 23535 39423
rect 23566 39420 23572 39432
rect 23523 39392 23572 39420
rect 23523 39389 23535 39392
rect 23477 39383 23535 39389
rect 23566 39380 23572 39392
rect 23624 39380 23630 39432
rect 23658 39380 23664 39432
rect 23716 39380 23722 39432
rect 25593 39423 25651 39429
rect 25593 39389 25605 39423
rect 25639 39420 25651 39423
rect 25866 39420 25872 39432
rect 25639 39392 25872 39420
rect 25639 39389 25651 39392
rect 25593 39383 25651 39389
rect 25866 39380 25872 39392
rect 25924 39380 25930 39432
rect 25976 39429 26004 39460
rect 25961 39423 26019 39429
rect 25961 39389 25973 39423
rect 26007 39389 26019 39423
rect 25961 39383 26019 39389
rect 26142 39380 26148 39432
rect 26200 39380 26206 39432
rect 23385 39355 23443 39361
rect 23385 39352 23397 39355
rect 21560 39324 23397 39352
rect 23385 39321 23397 39324
rect 23431 39352 23443 39355
rect 23431 39324 25820 39352
rect 23431 39321 23443 39324
rect 23385 39315 23443 39321
rect 22186 39284 22192 39296
rect 13004 39256 22192 39284
rect 22186 39244 22192 39256
rect 22244 39244 22250 39296
rect 23014 39244 23020 39296
rect 23072 39244 23078 39296
rect 23750 39244 23756 39296
rect 23808 39284 23814 39296
rect 25685 39287 25743 39293
rect 25685 39284 25697 39287
rect 23808 39256 25697 39284
rect 23808 39244 23814 39256
rect 25685 39253 25697 39256
rect 25731 39253 25743 39287
rect 25792 39284 25820 39324
rect 28626 39312 28632 39364
rect 28684 39352 28690 39364
rect 28813 39355 28871 39361
rect 28813 39352 28825 39355
rect 28684 39324 28825 39352
rect 28684 39312 28690 39324
rect 28813 39321 28825 39324
rect 28859 39321 28871 39355
rect 28920 39352 28948 39460
rect 31297 39457 31309 39491
rect 31343 39488 31355 39491
rect 33152 39488 33180 39516
rect 31343 39460 33180 39488
rect 31343 39457 31355 39460
rect 31297 39451 31355 39457
rect 30009 39423 30067 39429
rect 30009 39389 30021 39423
rect 30055 39420 30067 39423
rect 30190 39420 30196 39432
rect 30055 39392 30196 39420
rect 30055 39389 30067 39392
rect 30009 39383 30067 39389
rect 30190 39380 30196 39392
rect 30248 39380 30254 39432
rect 30742 39380 30748 39432
rect 30800 39380 30806 39432
rect 33134 39380 33140 39432
rect 33192 39420 33198 39432
rect 38194 39420 38200 39432
rect 33192 39392 38200 39420
rect 33192 39380 33198 39392
rect 38194 39380 38200 39392
rect 38252 39380 38258 39432
rect 32950 39352 32956 39364
rect 28920 39324 32956 39352
rect 28813 39315 28871 39321
rect 32950 39312 32956 39324
rect 33008 39312 33014 39364
rect 29914 39284 29920 39296
rect 25792 39256 29920 39284
rect 25685 39247 25743 39253
rect 29914 39244 29920 39256
rect 29972 39244 29978 39296
rect 31846 39244 31852 39296
rect 31904 39284 31910 39296
rect 32677 39287 32735 39293
rect 32677 39284 32689 39287
rect 31904 39256 32689 39284
rect 31904 39244 31910 39256
rect 32677 39253 32689 39256
rect 32723 39253 32735 39287
rect 32677 39247 32735 39253
rect 1104 39194 40848 39216
rect 1104 39142 2610 39194
rect 2662 39142 2674 39194
rect 2726 39142 2738 39194
rect 2790 39142 2802 39194
rect 2854 39142 2866 39194
rect 2918 39142 7610 39194
rect 7662 39142 7674 39194
rect 7726 39142 7738 39194
rect 7790 39142 7802 39194
rect 7854 39142 7866 39194
rect 7918 39142 12610 39194
rect 12662 39142 12674 39194
rect 12726 39142 12738 39194
rect 12790 39142 12802 39194
rect 12854 39142 12866 39194
rect 12918 39142 17610 39194
rect 17662 39142 17674 39194
rect 17726 39142 17738 39194
rect 17790 39142 17802 39194
rect 17854 39142 17866 39194
rect 17918 39142 22610 39194
rect 22662 39142 22674 39194
rect 22726 39142 22738 39194
rect 22790 39142 22802 39194
rect 22854 39142 22866 39194
rect 22918 39142 27610 39194
rect 27662 39142 27674 39194
rect 27726 39142 27738 39194
rect 27790 39142 27802 39194
rect 27854 39142 27866 39194
rect 27918 39142 32610 39194
rect 32662 39142 32674 39194
rect 32726 39142 32738 39194
rect 32790 39142 32802 39194
rect 32854 39142 32866 39194
rect 32918 39142 37610 39194
rect 37662 39142 37674 39194
rect 37726 39142 37738 39194
rect 37790 39142 37802 39194
rect 37854 39142 37866 39194
rect 37918 39142 40848 39194
rect 1104 39120 40848 39142
rect 9858 39040 9864 39092
rect 9916 39080 9922 39092
rect 16298 39080 16304 39092
rect 9916 39052 16304 39080
rect 9916 39040 9922 39052
rect 16298 39040 16304 39052
rect 16356 39040 16362 39092
rect 20438 39040 20444 39092
rect 20496 39080 20502 39092
rect 28718 39080 28724 39092
rect 20496 39052 28724 39080
rect 20496 39040 20502 39052
rect 28718 39040 28724 39052
rect 28776 39040 28782 39092
rect 30098 39040 30104 39092
rect 30156 39080 30162 39092
rect 32325 39083 32383 39089
rect 32325 39080 32337 39083
rect 30156 39052 32337 39080
rect 30156 39040 30162 39052
rect 32325 39049 32337 39052
rect 32371 39049 32383 39083
rect 32325 39043 32383 39049
rect 32493 39083 32551 39089
rect 32493 39049 32505 39083
rect 32539 39080 32551 39083
rect 33134 39080 33140 39092
rect 32539 39052 33140 39080
rect 32539 39049 32551 39052
rect 32493 39043 32551 39049
rect 33134 39040 33140 39052
rect 33192 39040 33198 39092
rect 26234 39012 26240 39024
rect 21284 38984 26240 39012
rect 20438 38904 20444 38956
rect 20496 38904 20502 38956
rect 21284 38953 21312 38984
rect 26234 38972 26240 38984
rect 26292 38972 26298 39024
rect 28810 38972 28816 39024
rect 28868 39012 28874 39024
rect 28948 39012 28954 39024
rect 28868 38984 28954 39012
rect 28868 38972 28874 38984
rect 28948 38972 28954 38984
rect 29006 38972 29012 39024
rect 30377 39015 30435 39021
rect 30377 38981 30389 39015
rect 30423 39012 30435 39015
rect 30466 39012 30472 39024
rect 30423 38984 30472 39012
rect 30423 38981 30435 38984
rect 30377 38975 30435 38981
rect 30466 38972 30472 38984
rect 30524 38972 30530 39024
rect 30558 38972 30564 39024
rect 30616 39012 30622 39024
rect 32125 39015 32183 39021
rect 32125 39012 32137 39015
rect 30616 38984 32137 39012
rect 30616 38972 30622 38984
rect 32125 38981 32137 38984
rect 32171 39012 32183 39015
rect 32769 39015 32827 39021
rect 32769 39012 32781 39015
rect 32171 38984 32781 39012
rect 32171 38981 32183 38984
rect 32125 38975 32183 38981
rect 32769 38981 32781 38984
rect 32815 38981 32827 39015
rect 32769 38975 32827 38981
rect 21269 38947 21327 38953
rect 21269 38913 21281 38947
rect 21315 38913 21327 38947
rect 21269 38907 21327 38913
rect 28626 38904 28632 38956
rect 28684 38944 28690 38956
rect 29086 38944 29092 38956
rect 28684 38916 29092 38944
rect 28684 38904 28690 38916
rect 29086 38904 29092 38916
rect 29144 38904 29150 38956
rect 29178 38904 29184 38956
rect 29236 38904 29242 38956
rect 29273 38947 29331 38953
rect 29273 38913 29285 38947
rect 29319 38944 29331 38947
rect 29641 38947 29699 38953
rect 29319 38916 29408 38944
rect 29319 38913 29331 38916
rect 29273 38907 29331 38913
rect 20352 38888 20404 38894
rect 29380 38888 29408 38916
rect 29641 38913 29653 38947
rect 29687 38944 29699 38947
rect 29730 38944 29736 38956
rect 29687 38916 29736 38944
rect 29687 38913 29699 38916
rect 29641 38907 29699 38913
rect 29730 38904 29736 38916
rect 29788 38904 29794 38956
rect 30742 38904 30748 38956
rect 30800 38904 30806 38956
rect 30926 38904 30932 38956
rect 30984 38904 30990 38956
rect 21545 38879 21603 38885
rect 21545 38845 21557 38879
rect 21591 38876 21603 38879
rect 21591 38848 23796 38876
rect 21591 38845 21603 38848
rect 21545 38839 21603 38845
rect 20352 38830 20404 38836
rect 20162 38768 20168 38820
rect 20220 38808 20226 38820
rect 20257 38811 20315 38817
rect 20257 38808 20269 38811
rect 20220 38780 20269 38808
rect 20220 38768 20226 38780
rect 20257 38777 20269 38780
rect 20303 38777 20315 38811
rect 20257 38771 20315 38777
rect 5074 38700 5080 38752
rect 5132 38740 5138 38752
rect 10226 38740 10232 38752
rect 5132 38712 10232 38740
rect 5132 38700 5138 38712
rect 10226 38700 10232 38712
rect 10284 38700 10290 38752
rect 23382 38700 23388 38752
rect 23440 38700 23446 38752
rect 23768 38740 23796 38848
rect 23842 38836 23848 38888
rect 23900 38836 23906 38888
rect 24302 38836 24308 38888
rect 24360 38876 24366 38888
rect 24360 38848 29132 38876
rect 24360 38836 24366 38848
rect 24578 38768 24584 38820
rect 24636 38808 24642 38820
rect 28994 38808 29000 38820
rect 24636 38780 29000 38808
rect 24636 38768 24642 38780
rect 28994 38768 29000 38780
rect 29052 38768 29058 38820
rect 29104 38752 29132 38848
rect 29362 38836 29368 38888
rect 29420 38836 29426 38888
rect 29546 38836 29552 38888
rect 29604 38836 29610 38888
rect 29178 38768 29184 38820
rect 29236 38808 29242 38820
rect 30760 38808 30788 38904
rect 29236 38780 30788 38808
rect 29236 38768 29242 38780
rect 28810 38740 28816 38752
rect 23768 38712 28816 38740
rect 28810 38700 28816 38712
rect 28868 38700 28874 38752
rect 29086 38700 29092 38752
rect 29144 38700 29150 38752
rect 30190 38700 30196 38752
rect 30248 38700 30254 38752
rect 32306 38700 32312 38752
rect 32364 38700 32370 38752
rect 1104 38650 40848 38672
rect 1104 38598 1950 38650
rect 2002 38598 2014 38650
rect 2066 38598 2078 38650
rect 2130 38598 2142 38650
rect 2194 38598 2206 38650
rect 2258 38598 6950 38650
rect 7002 38598 7014 38650
rect 7066 38598 7078 38650
rect 7130 38598 7142 38650
rect 7194 38598 7206 38650
rect 7258 38598 11950 38650
rect 12002 38598 12014 38650
rect 12066 38598 12078 38650
rect 12130 38598 12142 38650
rect 12194 38598 12206 38650
rect 12258 38598 16950 38650
rect 17002 38598 17014 38650
rect 17066 38598 17078 38650
rect 17130 38598 17142 38650
rect 17194 38598 17206 38650
rect 17258 38598 21950 38650
rect 22002 38598 22014 38650
rect 22066 38598 22078 38650
rect 22130 38598 22142 38650
rect 22194 38598 22206 38650
rect 22258 38598 26950 38650
rect 27002 38598 27014 38650
rect 27066 38598 27078 38650
rect 27130 38598 27142 38650
rect 27194 38598 27206 38650
rect 27258 38598 31950 38650
rect 32002 38598 32014 38650
rect 32066 38598 32078 38650
rect 32130 38598 32142 38650
rect 32194 38598 32206 38650
rect 32258 38598 36950 38650
rect 37002 38598 37014 38650
rect 37066 38598 37078 38650
rect 37130 38598 37142 38650
rect 37194 38598 37206 38650
rect 37258 38598 40848 38650
rect 1104 38576 40848 38598
rect 19518 38496 19524 38548
rect 19576 38496 19582 38548
rect 24118 38496 24124 38548
rect 24176 38536 24182 38548
rect 25133 38539 25191 38545
rect 25133 38536 25145 38539
rect 24176 38508 25145 38536
rect 24176 38496 24182 38508
rect 25133 38505 25145 38508
rect 25179 38505 25191 38539
rect 25133 38499 25191 38505
rect 32306 38496 32312 38548
rect 32364 38536 32370 38548
rect 33042 38536 33048 38548
rect 32364 38508 33048 38536
rect 32364 38496 32370 38508
rect 33042 38496 33048 38508
rect 33100 38496 33106 38548
rect 6454 38428 6460 38480
rect 6512 38468 6518 38480
rect 6512 38440 24900 38468
rect 6512 38428 6518 38440
rect 23842 38360 23848 38412
rect 23900 38400 23906 38412
rect 24762 38400 24768 38412
rect 23900 38372 24768 38400
rect 23900 38360 23906 38372
rect 24762 38360 24768 38372
rect 24820 38360 24826 38412
rect 19794 38292 19800 38344
rect 19852 38292 19858 38344
rect 24397 38335 24455 38341
rect 24397 38332 24409 38335
rect 22066 38304 24409 38332
rect 14826 38224 14832 38276
rect 14884 38264 14890 38276
rect 22066 38264 22094 38304
rect 24397 38301 24409 38304
rect 24443 38301 24455 38335
rect 24397 38295 24455 38301
rect 24578 38292 24584 38344
rect 24636 38292 24642 38344
rect 24673 38335 24731 38341
rect 24673 38301 24685 38335
rect 24719 38332 24731 38335
rect 24872 38332 24900 38440
rect 24719 38304 24900 38332
rect 24949 38335 25007 38341
rect 24719 38301 24731 38304
rect 24673 38295 24731 38301
rect 24949 38301 24961 38335
rect 24995 38332 25007 38335
rect 33686 38332 33692 38344
rect 24995 38304 33692 38332
rect 24995 38301 25007 38304
rect 24949 38295 25007 38301
rect 14884 38236 22094 38264
rect 24688 38264 24716 38295
rect 33686 38292 33692 38304
rect 33744 38292 33750 38344
rect 25866 38264 25872 38276
rect 24688 38236 25872 38264
rect 14884 38224 14890 38236
rect 25866 38224 25872 38236
rect 25924 38224 25930 38276
rect 10318 38156 10324 38208
rect 10376 38196 10382 38208
rect 19337 38199 19395 38205
rect 19337 38196 19349 38199
rect 10376 38168 19349 38196
rect 10376 38156 10382 38168
rect 19337 38165 19349 38168
rect 19383 38165 19395 38199
rect 19337 38159 19395 38165
rect 1104 38106 40848 38128
rect 1104 38054 2610 38106
rect 2662 38054 2674 38106
rect 2726 38054 2738 38106
rect 2790 38054 2802 38106
rect 2854 38054 2866 38106
rect 2918 38054 7610 38106
rect 7662 38054 7674 38106
rect 7726 38054 7738 38106
rect 7790 38054 7802 38106
rect 7854 38054 7866 38106
rect 7918 38054 12610 38106
rect 12662 38054 12674 38106
rect 12726 38054 12738 38106
rect 12790 38054 12802 38106
rect 12854 38054 12866 38106
rect 12918 38054 17610 38106
rect 17662 38054 17674 38106
rect 17726 38054 17738 38106
rect 17790 38054 17802 38106
rect 17854 38054 17866 38106
rect 17918 38054 22610 38106
rect 22662 38054 22674 38106
rect 22726 38054 22738 38106
rect 22790 38054 22802 38106
rect 22854 38054 22866 38106
rect 22918 38054 27610 38106
rect 27662 38054 27674 38106
rect 27726 38054 27738 38106
rect 27790 38054 27802 38106
rect 27854 38054 27866 38106
rect 27918 38054 32610 38106
rect 32662 38054 32674 38106
rect 32726 38054 32738 38106
rect 32790 38054 32802 38106
rect 32854 38054 32866 38106
rect 32918 38054 37610 38106
rect 37662 38054 37674 38106
rect 37726 38054 37738 38106
rect 37790 38054 37802 38106
rect 37854 38054 37866 38106
rect 37918 38054 40848 38106
rect 1104 38032 40848 38054
rect 32398 37952 32404 38004
rect 32456 37992 32462 38004
rect 37369 37995 37427 38001
rect 37369 37992 37381 37995
rect 32456 37964 37381 37992
rect 32456 37952 32462 37964
rect 37369 37961 37381 37964
rect 37415 37961 37427 37995
rect 37369 37955 37427 37961
rect 37553 37995 37611 38001
rect 37553 37961 37565 37995
rect 37599 37992 37611 37995
rect 38378 37992 38384 38004
rect 37599 37964 38384 37992
rect 37599 37961 37611 37964
rect 37553 37955 37611 37961
rect 38378 37952 38384 37964
rect 38436 37952 38442 38004
rect 11054 37884 11060 37936
rect 11112 37924 11118 37936
rect 14553 37927 14611 37933
rect 14553 37924 14565 37927
rect 11112 37896 14565 37924
rect 11112 37884 11118 37896
rect 14553 37893 14565 37896
rect 14599 37924 14611 37927
rect 15286 37924 15292 37936
rect 14599 37896 15292 37924
rect 14599 37893 14611 37896
rect 14553 37887 14611 37893
rect 15286 37884 15292 37896
rect 15344 37884 15350 37936
rect 25222 37884 25228 37936
rect 25280 37884 25286 37936
rect 25498 37884 25504 37936
rect 25556 37924 25562 37936
rect 25556 37896 26832 37924
rect 25556 37884 25562 37896
rect 26804 37868 26832 37896
rect 35526 37884 35532 37936
rect 35584 37924 35590 37936
rect 37645 37927 37703 37933
rect 37645 37924 37657 37927
rect 35584 37896 37657 37924
rect 35584 37884 35590 37896
rect 37645 37893 37657 37896
rect 37691 37893 37703 37927
rect 37645 37887 37703 37893
rect 8294 37816 8300 37868
rect 8352 37856 8358 37868
rect 12805 37859 12863 37865
rect 12805 37856 12817 37859
rect 8352 37828 12817 37856
rect 8352 37816 8358 37828
rect 12805 37825 12817 37828
rect 12851 37856 12863 37859
rect 16850 37856 16856 37868
rect 12851 37828 16856 37856
rect 12851 37825 12863 37828
rect 12805 37819 12863 37825
rect 16850 37816 16856 37828
rect 16908 37816 16914 37868
rect 25682 37816 25688 37868
rect 25740 37816 25746 37868
rect 25777 37859 25835 37865
rect 25777 37825 25789 37859
rect 25823 37825 25835 37859
rect 25777 37819 25835 37825
rect 25498 37748 25504 37800
rect 25556 37788 25562 37800
rect 25792 37788 25820 37819
rect 26786 37816 26792 37868
rect 26844 37856 26850 37868
rect 27065 37859 27123 37865
rect 27065 37856 27077 37859
rect 26844 37828 27077 37856
rect 26844 37816 26850 37828
rect 27065 37825 27077 37828
rect 27111 37825 27123 37859
rect 27065 37819 27123 37825
rect 27341 37859 27399 37865
rect 27341 37825 27353 37859
rect 27387 37856 27399 37859
rect 27430 37856 27436 37868
rect 27387 37828 27436 37856
rect 27387 37825 27399 37828
rect 27341 37819 27399 37825
rect 27430 37816 27436 37828
rect 27488 37816 27494 37868
rect 37737 37859 37795 37865
rect 37737 37825 37749 37859
rect 37783 37825 37795 37859
rect 37737 37819 37795 37825
rect 25556 37760 25820 37788
rect 25556 37748 25562 37760
rect 32582 37748 32588 37800
rect 32640 37788 32646 37800
rect 37752 37788 37780 37819
rect 32640 37760 37780 37788
rect 32640 37748 32646 37760
rect 18046 37680 18052 37732
rect 18104 37720 18110 37732
rect 27065 37723 27123 37729
rect 27065 37720 27077 37723
rect 18104 37692 27077 37720
rect 18104 37680 18110 37692
rect 27065 37689 27077 37692
rect 27111 37689 27123 37723
rect 27065 37683 27123 37689
rect 30466 37680 30472 37732
rect 30524 37720 30530 37732
rect 37921 37723 37979 37729
rect 37921 37720 37933 37723
rect 30524 37692 37933 37720
rect 30524 37680 30530 37692
rect 37921 37689 37933 37692
rect 37967 37689 37979 37723
rect 37921 37683 37979 37689
rect 25961 37655 26019 37661
rect 25961 37621 25973 37655
rect 26007 37652 26019 37655
rect 29546 37652 29552 37664
rect 26007 37624 29552 37652
rect 26007 37621 26019 37624
rect 25961 37615 26019 37621
rect 29546 37612 29552 37624
rect 29604 37612 29610 37664
rect 1104 37562 40848 37584
rect 1104 37510 1950 37562
rect 2002 37510 2014 37562
rect 2066 37510 2078 37562
rect 2130 37510 2142 37562
rect 2194 37510 2206 37562
rect 2258 37510 6950 37562
rect 7002 37510 7014 37562
rect 7066 37510 7078 37562
rect 7130 37510 7142 37562
rect 7194 37510 7206 37562
rect 7258 37510 11950 37562
rect 12002 37510 12014 37562
rect 12066 37510 12078 37562
rect 12130 37510 12142 37562
rect 12194 37510 12206 37562
rect 12258 37510 16950 37562
rect 17002 37510 17014 37562
rect 17066 37510 17078 37562
rect 17130 37510 17142 37562
rect 17194 37510 17206 37562
rect 17258 37510 21950 37562
rect 22002 37510 22014 37562
rect 22066 37510 22078 37562
rect 22130 37510 22142 37562
rect 22194 37510 22206 37562
rect 22258 37510 26950 37562
rect 27002 37510 27014 37562
rect 27066 37510 27078 37562
rect 27130 37510 27142 37562
rect 27194 37510 27206 37562
rect 27258 37510 31950 37562
rect 32002 37510 32014 37562
rect 32066 37510 32078 37562
rect 32130 37510 32142 37562
rect 32194 37510 32206 37562
rect 32258 37510 36950 37562
rect 37002 37510 37014 37562
rect 37066 37510 37078 37562
rect 37130 37510 37142 37562
rect 37194 37510 37206 37562
rect 37258 37510 40848 37562
rect 1104 37488 40848 37510
rect 18417 37451 18475 37457
rect 18417 37417 18429 37451
rect 18463 37448 18475 37451
rect 18598 37448 18604 37460
rect 18463 37420 18604 37448
rect 18463 37417 18475 37420
rect 18417 37411 18475 37417
rect 18598 37408 18604 37420
rect 18656 37408 18662 37460
rect 28074 37408 28080 37460
rect 28132 37448 28138 37460
rect 28132 37420 35894 37448
rect 28132 37408 28138 37420
rect 8386 37340 8392 37392
rect 8444 37380 8450 37392
rect 25498 37380 25504 37392
rect 8444 37352 25504 37380
rect 8444 37340 8450 37352
rect 25498 37340 25504 37352
rect 25556 37340 25562 37392
rect 26602 37340 26608 37392
rect 26660 37380 26666 37392
rect 28534 37380 28540 37392
rect 26660 37352 28540 37380
rect 26660 37340 26666 37352
rect 28534 37340 28540 37352
rect 28592 37340 28598 37392
rect 32490 37380 32496 37392
rect 31726 37352 32496 37380
rect 17402 37272 17408 37324
rect 17460 37312 17466 37324
rect 18966 37312 18972 37324
rect 17460 37284 18972 37312
rect 17460 37272 17466 37284
rect 18966 37272 18972 37284
rect 19024 37272 19030 37324
rect 31726 37312 31754 37352
rect 32490 37340 32496 37352
rect 32548 37340 32554 37392
rect 35866 37380 35894 37420
rect 39393 37383 39451 37389
rect 39393 37380 39405 37383
rect 35866 37352 39405 37380
rect 39393 37349 39405 37352
rect 39439 37349 39451 37383
rect 39393 37343 39451 37349
rect 19076 37284 31754 37312
rect 18509 37247 18567 37253
rect 18509 37244 18521 37247
rect 17604 37216 18521 37244
rect 16758 37068 16764 37120
rect 16816 37108 16822 37120
rect 17604 37117 17632 37216
rect 18509 37213 18521 37216
rect 18555 37244 18567 37247
rect 19076 37244 19104 37284
rect 18555 37216 19104 37244
rect 18555 37213 18567 37216
rect 18509 37207 18567 37213
rect 34698 37204 34704 37256
rect 34756 37244 34762 37256
rect 34882 37244 34888 37256
rect 34756 37216 34888 37244
rect 34756 37204 34762 37216
rect 34882 37204 34888 37216
rect 34940 37244 34946 37256
rect 35161 37247 35219 37253
rect 35161 37244 35173 37247
rect 34940 37216 35173 37244
rect 34940 37204 34946 37216
rect 35161 37213 35173 37216
rect 35207 37213 35219 37247
rect 35161 37207 35219 37213
rect 38838 37204 38844 37256
rect 38896 37204 38902 37256
rect 39022 37204 39028 37256
rect 39080 37204 39086 37256
rect 39209 37247 39267 37253
rect 39209 37213 39221 37247
rect 39255 37213 39267 37247
rect 39209 37207 39267 37213
rect 31202 37136 31208 37188
rect 31260 37176 31266 37188
rect 39224 37176 39252 37207
rect 31260 37148 39252 37176
rect 31260 37136 31266 37148
rect 17589 37111 17647 37117
rect 17589 37108 17601 37111
rect 16816 37080 17601 37108
rect 16816 37068 16822 37080
rect 17589 37077 17601 37080
rect 17635 37077 17647 37111
rect 17589 37071 17647 37077
rect 17954 37068 17960 37120
rect 18012 37108 18018 37120
rect 18049 37111 18107 37117
rect 18049 37108 18061 37111
rect 18012 37080 18061 37108
rect 18012 37068 18018 37080
rect 18049 37077 18061 37080
rect 18095 37077 18107 37111
rect 18049 37071 18107 37077
rect 35621 37111 35679 37117
rect 35621 37077 35633 37111
rect 35667 37108 35679 37111
rect 38010 37108 38016 37120
rect 35667 37080 38016 37108
rect 35667 37077 35679 37080
rect 35621 37071 35679 37077
rect 38010 37068 38016 37080
rect 38068 37068 38074 37120
rect 1104 37018 40848 37040
rect 1104 36966 2610 37018
rect 2662 36966 2674 37018
rect 2726 36966 2738 37018
rect 2790 36966 2802 37018
rect 2854 36966 2866 37018
rect 2918 36966 7610 37018
rect 7662 36966 7674 37018
rect 7726 36966 7738 37018
rect 7790 36966 7802 37018
rect 7854 36966 7866 37018
rect 7918 36966 12610 37018
rect 12662 36966 12674 37018
rect 12726 36966 12738 37018
rect 12790 36966 12802 37018
rect 12854 36966 12866 37018
rect 12918 36966 17610 37018
rect 17662 36966 17674 37018
rect 17726 36966 17738 37018
rect 17790 36966 17802 37018
rect 17854 36966 17866 37018
rect 17918 36966 22610 37018
rect 22662 36966 22674 37018
rect 22726 36966 22738 37018
rect 22790 36966 22802 37018
rect 22854 36966 22866 37018
rect 22918 36966 27610 37018
rect 27662 36966 27674 37018
rect 27726 36966 27738 37018
rect 27790 36966 27802 37018
rect 27854 36966 27866 37018
rect 27918 36966 32610 37018
rect 32662 36966 32674 37018
rect 32726 36966 32738 37018
rect 32790 36966 32802 37018
rect 32854 36966 32866 37018
rect 32918 36966 37610 37018
rect 37662 36966 37674 37018
rect 37726 36966 37738 37018
rect 37790 36966 37802 37018
rect 37854 36966 37866 37018
rect 37918 36966 40848 37018
rect 1104 36944 40848 36966
rect 24949 36839 25007 36845
rect 24949 36805 24961 36839
rect 24995 36836 25007 36839
rect 26602 36836 26608 36848
rect 24995 36808 26608 36836
rect 24995 36805 25007 36808
rect 24949 36799 25007 36805
rect 26602 36796 26608 36808
rect 26660 36796 26666 36848
rect 38102 36796 38108 36848
rect 38160 36836 38166 36848
rect 38197 36839 38255 36845
rect 38197 36836 38209 36839
rect 38160 36808 38209 36836
rect 38160 36796 38166 36808
rect 38197 36805 38209 36808
rect 38243 36805 38255 36839
rect 38197 36799 38255 36805
rect 23474 36728 23480 36780
rect 23532 36768 23538 36780
rect 23934 36768 23940 36780
rect 23532 36740 23940 36768
rect 23532 36728 23538 36740
rect 23934 36728 23940 36740
rect 23992 36728 23998 36780
rect 24397 36771 24455 36777
rect 24397 36737 24409 36771
rect 24443 36768 24455 36771
rect 30374 36768 30380 36780
rect 24443 36740 30380 36768
rect 24443 36737 24455 36740
rect 24397 36731 24455 36737
rect 30374 36728 30380 36740
rect 30432 36728 30438 36780
rect 37921 36771 37979 36777
rect 37921 36737 37933 36771
rect 37967 36737 37979 36771
rect 37921 36731 37979 36737
rect 37936 36700 37964 36731
rect 38010 36728 38016 36780
rect 38068 36728 38074 36780
rect 38562 36700 38568 36712
rect 37936 36672 38568 36700
rect 38562 36660 38568 36672
rect 38620 36660 38626 36712
rect 15286 36524 15292 36576
rect 15344 36564 15350 36576
rect 18690 36564 18696 36576
rect 15344 36536 18696 36564
rect 15344 36524 15350 36536
rect 18690 36524 18696 36536
rect 18748 36524 18754 36576
rect 1104 36474 40848 36496
rect 1104 36422 1950 36474
rect 2002 36422 2014 36474
rect 2066 36422 2078 36474
rect 2130 36422 2142 36474
rect 2194 36422 2206 36474
rect 2258 36422 6950 36474
rect 7002 36422 7014 36474
rect 7066 36422 7078 36474
rect 7130 36422 7142 36474
rect 7194 36422 7206 36474
rect 7258 36422 11950 36474
rect 12002 36422 12014 36474
rect 12066 36422 12078 36474
rect 12130 36422 12142 36474
rect 12194 36422 12206 36474
rect 12258 36422 16950 36474
rect 17002 36422 17014 36474
rect 17066 36422 17078 36474
rect 17130 36422 17142 36474
rect 17194 36422 17206 36474
rect 17258 36422 21950 36474
rect 22002 36422 22014 36474
rect 22066 36422 22078 36474
rect 22130 36422 22142 36474
rect 22194 36422 22206 36474
rect 22258 36422 26950 36474
rect 27002 36422 27014 36474
rect 27066 36422 27078 36474
rect 27130 36422 27142 36474
rect 27194 36422 27206 36474
rect 27258 36422 31950 36474
rect 32002 36422 32014 36474
rect 32066 36422 32078 36474
rect 32130 36422 32142 36474
rect 32194 36422 32206 36474
rect 32258 36422 36950 36474
rect 37002 36422 37014 36474
rect 37066 36422 37078 36474
rect 37130 36422 37142 36474
rect 37194 36422 37206 36474
rect 37258 36422 40848 36474
rect 1104 36400 40848 36422
rect 9861 36363 9919 36369
rect 9861 36329 9873 36363
rect 9907 36360 9919 36363
rect 11698 36360 11704 36372
rect 9907 36332 11704 36360
rect 9907 36329 9919 36332
rect 9861 36323 9919 36329
rect 11698 36320 11704 36332
rect 11756 36320 11762 36372
rect 30282 36252 30288 36304
rect 30340 36292 30346 36304
rect 30742 36292 30748 36304
rect 30340 36264 30748 36292
rect 30340 36252 30346 36264
rect 30742 36252 30748 36264
rect 30800 36292 30806 36304
rect 35437 36295 35495 36301
rect 35437 36292 35449 36295
rect 30800 36264 35449 36292
rect 30800 36252 30806 36264
rect 35437 36261 35449 36264
rect 35483 36261 35495 36295
rect 35437 36255 35495 36261
rect 10962 36224 10968 36236
rect 9692 36196 10968 36224
rect 9582 36116 9588 36168
rect 9640 36156 9646 36168
rect 9692 36165 9720 36196
rect 10962 36184 10968 36196
rect 11020 36184 11026 36236
rect 20070 36184 20076 36236
rect 20128 36224 20134 36236
rect 20128 36196 34928 36224
rect 20128 36184 20134 36196
rect 9677 36159 9735 36165
rect 9677 36156 9689 36159
rect 9640 36128 9689 36156
rect 9640 36116 9646 36128
rect 9677 36125 9689 36128
rect 9723 36125 9735 36159
rect 9677 36119 9735 36125
rect 9861 36159 9919 36165
rect 9861 36125 9873 36159
rect 9907 36156 9919 36159
rect 28258 36156 28264 36168
rect 9907 36128 28264 36156
rect 9907 36125 9919 36128
rect 9861 36119 9919 36125
rect 28258 36116 28264 36128
rect 28316 36116 28322 36168
rect 34900 36165 34928 36196
rect 34885 36159 34943 36165
rect 34885 36125 34897 36159
rect 34931 36125 34943 36159
rect 34885 36119 34943 36125
rect 35066 36116 35072 36168
rect 35124 36116 35130 36168
rect 35250 36116 35256 36168
rect 35308 36116 35314 36168
rect 1104 35930 40848 35952
rect 1104 35878 2610 35930
rect 2662 35878 2674 35930
rect 2726 35878 2738 35930
rect 2790 35878 2802 35930
rect 2854 35878 2866 35930
rect 2918 35878 7610 35930
rect 7662 35878 7674 35930
rect 7726 35878 7738 35930
rect 7790 35878 7802 35930
rect 7854 35878 7866 35930
rect 7918 35878 12610 35930
rect 12662 35878 12674 35930
rect 12726 35878 12738 35930
rect 12790 35878 12802 35930
rect 12854 35878 12866 35930
rect 12918 35878 17610 35930
rect 17662 35878 17674 35930
rect 17726 35878 17738 35930
rect 17790 35878 17802 35930
rect 17854 35878 17866 35930
rect 17918 35878 22610 35930
rect 22662 35878 22674 35930
rect 22726 35878 22738 35930
rect 22790 35878 22802 35930
rect 22854 35878 22866 35930
rect 22918 35878 27610 35930
rect 27662 35878 27674 35930
rect 27726 35878 27738 35930
rect 27790 35878 27802 35930
rect 27854 35878 27866 35930
rect 27918 35878 32610 35930
rect 32662 35878 32674 35930
rect 32726 35878 32738 35930
rect 32790 35878 32802 35930
rect 32854 35878 32866 35930
rect 32918 35878 37610 35930
rect 37662 35878 37674 35930
rect 37726 35878 37738 35930
rect 37790 35878 37802 35930
rect 37854 35878 37866 35930
rect 37918 35878 40848 35930
rect 1104 35856 40848 35878
rect 3881 35819 3939 35825
rect 3881 35785 3893 35819
rect 3927 35816 3939 35819
rect 3970 35816 3976 35828
rect 3927 35788 3976 35816
rect 3927 35785 3939 35788
rect 3881 35779 3939 35785
rect 3970 35776 3976 35788
rect 4028 35776 4034 35828
rect 7466 35776 7472 35828
rect 7524 35816 7530 35828
rect 7650 35816 7656 35828
rect 7524 35788 7656 35816
rect 7524 35776 7530 35788
rect 7650 35776 7656 35788
rect 7708 35776 7714 35828
rect 10226 35776 10232 35828
rect 10284 35816 10290 35828
rect 23198 35816 23204 35828
rect 10284 35788 23204 35816
rect 10284 35776 10290 35788
rect 23198 35776 23204 35788
rect 23256 35816 23262 35828
rect 23382 35816 23388 35828
rect 23256 35788 23388 35816
rect 23256 35776 23262 35788
rect 23382 35776 23388 35788
rect 23440 35776 23446 35828
rect 31754 35816 31760 35828
rect 26896 35788 31760 35816
rect 9766 35708 9772 35760
rect 9824 35748 9830 35760
rect 9824 35720 16620 35748
rect 9824 35708 9830 35720
rect 4065 35683 4123 35689
rect 4065 35649 4077 35683
rect 4111 35649 4123 35683
rect 4065 35643 4123 35649
rect 4080 35612 4108 35643
rect 4154 35640 4160 35692
rect 4212 35640 4218 35692
rect 4433 35683 4491 35689
rect 4433 35649 4445 35683
rect 4479 35680 4491 35683
rect 14182 35680 14188 35692
rect 4479 35652 14188 35680
rect 4479 35649 4491 35652
rect 4433 35643 4491 35649
rect 14182 35640 14188 35652
rect 14240 35680 14246 35692
rect 15010 35680 15016 35692
rect 14240 35652 15016 35680
rect 14240 35640 14246 35652
rect 15010 35640 15016 35652
rect 15068 35640 15074 35692
rect 16592 35680 16620 35720
rect 16666 35708 16672 35760
rect 16724 35748 16730 35760
rect 26896 35748 26924 35788
rect 31754 35776 31760 35788
rect 31812 35776 31818 35828
rect 16724 35720 26924 35748
rect 29825 35751 29883 35757
rect 16724 35708 16730 35720
rect 29825 35717 29837 35751
rect 29871 35748 29883 35751
rect 31846 35748 31852 35760
rect 29871 35720 31852 35748
rect 29871 35717 29883 35720
rect 29825 35711 29883 35717
rect 31846 35708 31852 35720
rect 31904 35708 31910 35760
rect 16592 35652 16988 35680
rect 6086 35612 6092 35624
rect 4080 35584 6092 35612
rect 6086 35572 6092 35584
rect 6144 35612 6150 35624
rect 16482 35612 16488 35624
rect 6144 35584 16488 35612
rect 6144 35572 6150 35584
rect 16482 35572 16488 35584
rect 16540 35612 16546 35624
rect 16850 35612 16856 35624
rect 16540 35584 16856 35612
rect 16540 35572 16546 35584
rect 16850 35572 16856 35584
rect 16908 35572 16914 35624
rect 16960 35612 16988 35652
rect 17218 35640 17224 35692
rect 17276 35680 17282 35692
rect 17586 35680 17592 35692
rect 17276 35652 17592 35680
rect 17276 35640 17282 35652
rect 17586 35640 17592 35652
rect 17644 35640 17650 35692
rect 24946 35640 24952 35692
rect 25004 35680 25010 35692
rect 26142 35680 26148 35692
rect 25004 35652 26148 35680
rect 25004 35640 25010 35652
rect 26142 35640 26148 35652
rect 26200 35640 26206 35692
rect 26602 35640 26608 35692
rect 26660 35680 26666 35692
rect 30193 35683 30251 35689
rect 30193 35680 30205 35683
rect 26660 35652 30205 35680
rect 26660 35640 26666 35652
rect 30193 35649 30205 35652
rect 30239 35649 30251 35683
rect 30193 35643 30251 35649
rect 30285 35683 30343 35689
rect 30285 35649 30297 35683
rect 30331 35680 30343 35683
rect 30466 35680 30472 35692
rect 30331 35652 30472 35680
rect 30331 35649 30343 35652
rect 30285 35643 30343 35649
rect 16960 35584 17356 35612
rect 3970 35504 3976 35556
rect 4028 35544 4034 35556
rect 16390 35544 16396 35556
rect 4028 35516 16396 35544
rect 4028 35504 4034 35516
rect 16390 35504 16396 35516
rect 16448 35504 16454 35556
rect 17328 35544 17356 35584
rect 17678 35572 17684 35624
rect 17736 35612 17742 35624
rect 17736 35584 25084 35612
rect 17736 35572 17742 35584
rect 19242 35544 19248 35556
rect 17328 35516 19248 35544
rect 19242 35504 19248 35516
rect 19300 35504 19306 35556
rect 4341 35479 4399 35485
rect 4341 35445 4353 35479
rect 4387 35476 4399 35479
rect 24946 35476 24952 35488
rect 4387 35448 24952 35476
rect 4387 35445 4399 35448
rect 4341 35439 4399 35445
rect 24946 35436 24952 35448
rect 25004 35436 25010 35488
rect 25056 35476 25084 35584
rect 29454 35572 29460 35624
rect 29512 35612 29518 35624
rect 30101 35615 30159 35621
rect 30101 35612 30113 35615
rect 29512 35584 30113 35612
rect 29512 35572 29518 35584
rect 30101 35581 30113 35584
rect 30147 35581 30159 35615
rect 30101 35575 30159 35581
rect 25130 35504 25136 35556
rect 25188 35544 25194 35556
rect 29365 35547 29423 35553
rect 29365 35544 29377 35547
rect 25188 35516 29377 35544
rect 25188 35504 25194 35516
rect 29365 35513 29377 35516
rect 29411 35513 29423 35547
rect 30208 35544 30236 35643
rect 30466 35640 30472 35652
rect 30524 35640 30530 35692
rect 36538 35612 36544 35624
rect 31726 35584 36544 35612
rect 31726 35544 31754 35584
rect 36538 35572 36544 35584
rect 36596 35572 36602 35624
rect 30208 35516 31754 35544
rect 29365 35507 29423 35513
rect 30466 35476 30472 35488
rect 25056 35448 30472 35476
rect 30466 35436 30472 35448
rect 30524 35436 30530 35488
rect 1104 35386 40848 35408
rect 1104 35334 1950 35386
rect 2002 35334 2014 35386
rect 2066 35334 2078 35386
rect 2130 35334 2142 35386
rect 2194 35334 2206 35386
rect 2258 35334 6950 35386
rect 7002 35334 7014 35386
rect 7066 35334 7078 35386
rect 7130 35334 7142 35386
rect 7194 35334 7206 35386
rect 7258 35334 11950 35386
rect 12002 35334 12014 35386
rect 12066 35334 12078 35386
rect 12130 35334 12142 35386
rect 12194 35334 12206 35386
rect 12258 35334 16950 35386
rect 17002 35334 17014 35386
rect 17066 35334 17078 35386
rect 17130 35334 17142 35386
rect 17194 35334 17206 35386
rect 17258 35334 21950 35386
rect 22002 35334 22014 35386
rect 22066 35334 22078 35386
rect 22130 35334 22142 35386
rect 22194 35334 22206 35386
rect 22258 35334 26950 35386
rect 27002 35334 27014 35386
rect 27066 35334 27078 35386
rect 27130 35334 27142 35386
rect 27194 35334 27206 35386
rect 27258 35334 31950 35386
rect 32002 35334 32014 35386
rect 32066 35334 32078 35386
rect 32130 35334 32142 35386
rect 32194 35334 32206 35386
rect 32258 35334 36950 35386
rect 37002 35334 37014 35386
rect 37066 35334 37078 35386
rect 37130 35334 37142 35386
rect 37194 35334 37206 35386
rect 37258 35334 40848 35386
rect 1104 35312 40848 35334
rect 3786 35232 3792 35284
rect 3844 35272 3850 35284
rect 3881 35275 3939 35281
rect 3881 35272 3893 35275
rect 3844 35244 3893 35272
rect 3844 35232 3850 35244
rect 3881 35241 3893 35244
rect 3927 35241 3939 35275
rect 3881 35235 3939 35241
rect 4065 35275 4123 35281
rect 4065 35241 4077 35275
rect 4111 35272 4123 35275
rect 6730 35272 6736 35284
rect 4111 35244 6736 35272
rect 4111 35241 4123 35244
rect 4065 35235 4123 35241
rect 6730 35232 6736 35244
rect 6788 35232 6794 35284
rect 7190 35232 7196 35284
rect 7248 35272 7254 35284
rect 9766 35272 9772 35284
rect 7248 35244 9772 35272
rect 7248 35232 7254 35244
rect 9766 35232 9772 35244
rect 9824 35232 9830 35284
rect 10413 35275 10471 35281
rect 10413 35241 10425 35275
rect 10459 35272 10471 35275
rect 10502 35272 10508 35284
rect 10459 35244 10508 35272
rect 10459 35241 10471 35244
rect 10413 35235 10471 35241
rect 10502 35232 10508 35244
rect 10560 35232 10566 35284
rect 3513 35207 3571 35213
rect 3513 35173 3525 35207
rect 3559 35204 3571 35207
rect 6638 35204 6644 35216
rect 3559 35176 6644 35204
rect 3559 35173 3571 35176
rect 3513 35167 3571 35173
rect 6638 35164 6644 35176
rect 6696 35164 6702 35216
rect 19886 35164 19892 35216
rect 19944 35204 19950 35216
rect 19944 35176 22094 35204
rect 19944 35164 19950 35176
rect 5994 35136 6000 35148
rect 3344 35108 6000 35136
rect 3344 35077 3372 35108
rect 5994 35096 6000 35108
rect 6052 35136 6058 35148
rect 11054 35136 11060 35148
rect 6052 35108 11060 35136
rect 6052 35096 6058 35108
rect 3237 35071 3295 35077
rect 3237 35037 3249 35071
rect 3283 35037 3295 35071
rect 3237 35031 3295 35037
rect 3329 35071 3387 35077
rect 3329 35037 3341 35071
rect 3375 35037 3387 35071
rect 3329 35031 3387 35037
rect 3513 35071 3571 35077
rect 3513 35037 3525 35071
rect 3559 35068 3571 35071
rect 6454 35068 6460 35080
rect 3559 35040 6460 35068
rect 3559 35037 3571 35040
rect 3513 35031 3571 35037
rect 3252 35000 3280 35031
rect 6454 35028 6460 35040
rect 6512 35028 6518 35080
rect 7466 35028 7472 35080
rect 7524 35068 7530 35080
rect 7650 35068 7656 35080
rect 7524 35040 7656 35068
rect 7524 35028 7530 35040
rect 7650 35028 7656 35040
rect 7708 35028 7714 35080
rect 9766 35028 9772 35080
rect 9824 35028 9830 35080
rect 9858 35028 9864 35080
rect 9916 35028 9922 35080
rect 10060 35077 10088 35108
rect 11054 35096 11060 35108
rect 11112 35096 11118 35148
rect 12434 35096 12440 35148
rect 12492 35096 12498 35148
rect 13998 35136 14004 35148
rect 13188 35108 14004 35136
rect 10045 35071 10103 35077
rect 10045 35037 10057 35071
rect 10091 35037 10103 35071
rect 10045 35031 10103 35037
rect 10226 35028 10232 35080
rect 10284 35028 10290 35080
rect 12980 35071 13038 35077
rect 12980 35037 12992 35071
rect 13026 35068 13038 35071
rect 13078 35068 13084 35080
rect 13026 35040 13084 35068
rect 13026 35037 13038 35040
rect 12980 35031 13038 35037
rect 13078 35028 13084 35040
rect 13136 35028 13142 35080
rect 13188 35077 13216 35108
rect 13998 35096 14004 35108
rect 14056 35136 14062 35148
rect 14826 35136 14832 35148
rect 14056 35108 14832 35136
rect 14056 35096 14062 35108
rect 14826 35096 14832 35108
rect 14884 35096 14890 35148
rect 16390 35096 16396 35148
rect 16448 35136 16454 35148
rect 16448 35108 16620 35136
rect 16448 35096 16454 35108
rect 13173 35071 13231 35077
rect 13173 35037 13185 35071
rect 13219 35037 13231 35071
rect 13173 35031 13231 35037
rect 13538 35028 13544 35080
rect 13596 35028 13602 35080
rect 13722 35028 13728 35080
rect 13780 35028 13786 35080
rect 13814 35028 13820 35080
rect 13872 35028 13878 35080
rect 16485 35071 16543 35077
rect 16485 35037 16497 35071
rect 16531 35037 16543 35071
rect 16592 35068 16620 35108
rect 16666 35096 16672 35148
rect 16724 35096 16730 35148
rect 22066 35136 22094 35176
rect 23106 35164 23112 35216
rect 23164 35204 23170 35216
rect 23164 35176 27200 35204
rect 23164 35164 23170 35176
rect 27172 35145 27200 35176
rect 33134 35164 33140 35216
rect 33192 35204 33198 35216
rect 34146 35204 34152 35216
rect 33192 35176 34152 35204
rect 33192 35164 33198 35176
rect 34146 35164 34152 35176
rect 34204 35204 34210 35216
rect 38930 35204 38936 35216
rect 34204 35176 38936 35204
rect 34204 35164 34210 35176
rect 38930 35164 38936 35176
rect 38988 35164 38994 35216
rect 27157 35139 27215 35145
rect 22066 35108 27016 35136
rect 17037 35071 17095 35077
rect 17037 35068 17049 35071
rect 16592 35040 17049 35068
rect 16485 35031 16543 35037
rect 17037 35037 17049 35040
rect 17083 35068 17095 35071
rect 17678 35068 17684 35080
rect 17083 35040 17684 35068
rect 17083 35037 17095 35040
rect 17037 35031 17095 35037
rect 4249 35003 4307 35009
rect 3252 34972 4200 35000
rect 4062 34892 4068 34944
rect 4120 34892 4126 34944
rect 4172 34932 4200 34972
rect 4249 34969 4261 35003
rect 4295 35000 4307 35003
rect 8110 35000 8116 35012
rect 4295 34972 8116 35000
rect 4295 34969 4307 34972
rect 4249 34963 4307 34969
rect 8110 34960 8116 34972
rect 8168 34960 8174 35012
rect 10137 35003 10195 35009
rect 10137 34969 10149 35003
rect 10183 34969 10195 35003
rect 10137 34963 10195 34969
rect 6454 34932 6460 34944
rect 4172 34904 6460 34932
rect 6454 34892 6460 34904
rect 6512 34932 6518 34944
rect 10152 34932 10180 34963
rect 16500 34932 16528 35031
rect 17678 35028 17684 35040
rect 17736 35028 17742 35080
rect 25866 35028 25872 35080
rect 25924 35068 25930 35080
rect 26988 35077 27016 35108
rect 27157 35105 27169 35139
rect 27203 35136 27215 35139
rect 27203 35108 31754 35136
rect 27203 35105 27215 35108
rect 27157 35099 27215 35105
rect 26605 35071 26663 35077
rect 26605 35068 26617 35071
rect 25924 35040 26617 35068
rect 25924 35028 25930 35040
rect 26605 35037 26617 35040
rect 26651 35068 26663 35071
rect 26973 35071 27031 35077
rect 26651 35040 26832 35068
rect 26651 35037 26663 35040
rect 26605 35031 26663 35037
rect 17586 34960 17592 35012
rect 17644 35000 17650 35012
rect 26697 35003 26755 35009
rect 26697 35000 26709 35003
rect 17644 34972 26709 35000
rect 17644 34960 17650 34972
rect 26697 34969 26709 34972
rect 26743 34969 26755 35003
rect 26697 34963 26755 34969
rect 26602 34932 26608 34944
rect 6512 34904 26608 34932
rect 6512 34892 6518 34904
rect 26602 34892 26608 34904
rect 26660 34892 26666 34944
rect 26804 34932 26832 35040
rect 26973 35037 26985 35071
rect 27019 35037 27031 35071
rect 31726 35068 31754 35108
rect 31726 35040 35894 35068
rect 26973 35031 27031 35037
rect 26988 35000 27016 35031
rect 35434 35000 35440 35012
rect 26988 34972 35440 35000
rect 35434 34960 35440 34972
rect 35492 34960 35498 35012
rect 29638 34932 29644 34944
rect 26804 34904 29644 34932
rect 29638 34892 29644 34904
rect 29696 34892 29702 34944
rect 35866 34932 35894 35040
rect 38378 34932 38384 34944
rect 35866 34904 38384 34932
rect 38378 34892 38384 34904
rect 38436 34892 38442 34944
rect 1104 34842 40848 34864
rect 1104 34790 2610 34842
rect 2662 34790 2674 34842
rect 2726 34790 2738 34842
rect 2790 34790 2802 34842
rect 2854 34790 2866 34842
rect 2918 34790 7610 34842
rect 7662 34790 7674 34842
rect 7726 34790 7738 34842
rect 7790 34790 7802 34842
rect 7854 34790 7866 34842
rect 7918 34790 12610 34842
rect 12662 34790 12674 34842
rect 12726 34790 12738 34842
rect 12790 34790 12802 34842
rect 12854 34790 12866 34842
rect 12918 34790 17610 34842
rect 17662 34790 17674 34842
rect 17726 34790 17738 34842
rect 17790 34790 17802 34842
rect 17854 34790 17866 34842
rect 17918 34790 22610 34842
rect 22662 34790 22674 34842
rect 22726 34790 22738 34842
rect 22790 34790 22802 34842
rect 22854 34790 22866 34842
rect 22918 34790 27610 34842
rect 27662 34790 27674 34842
rect 27726 34790 27738 34842
rect 27790 34790 27802 34842
rect 27854 34790 27866 34842
rect 27918 34790 32610 34842
rect 32662 34790 32674 34842
rect 32726 34790 32738 34842
rect 32790 34790 32802 34842
rect 32854 34790 32866 34842
rect 32918 34790 37610 34842
rect 37662 34790 37674 34842
rect 37726 34790 37738 34842
rect 37790 34790 37802 34842
rect 37854 34790 37866 34842
rect 37918 34790 40848 34842
rect 1104 34768 40848 34790
rect 7561 34731 7619 34737
rect 7561 34697 7573 34731
rect 7607 34728 7619 34731
rect 7607 34700 12434 34728
rect 7607 34697 7619 34700
rect 7561 34691 7619 34697
rect 7190 34620 7196 34672
rect 7248 34620 7254 34672
rect 7285 34663 7343 34669
rect 7285 34629 7297 34663
rect 7331 34660 7343 34663
rect 7466 34660 7472 34672
rect 7331 34632 7472 34660
rect 7331 34629 7343 34632
rect 7285 34623 7343 34629
rect 7466 34620 7472 34632
rect 7524 34660 7530 34672
rect 8110 34660 8116 34672
rect 7524 34632 8116 34660
rect 7524 34620 7530 34632
rect 8110 34620 8116 34632
rect 8168 34620 8174 34672
rect 7009 34595 7067 34601
rect 7009 34561 7021 34595
rect 7055 34561 7067 34595
rect 7009 34555 7067 34561
rect 7024 34524 7052 34555
rect 7374 34552 7380 34604
rect 7432 34552 7438 34604
rect 12406 34592 12434 34700
rect 18690 34688 18696 34740
rect 18748 34728 18754 34740
rect 23106 34728 23112 34740
rect 18748 34700 23112 34728
rect 18748 34688 18754 34700
rect 23106 34688 23112 34700
rect 23164 34688 23170 34740
rect 36722 34688 36728 34740
rect 36780 34728 36786 34740
rect 38105 34731 38163 34737
rect 38105 34728 38117 34731
rect 36780 34700 38117 34728
rect 36780 34688 36786 34700
rect 38105 34697 38117 34700
rect 38151 34697 38163 34731
rect 38105 34691 38163 34697
rect 16850 34620 16856 34672
rect 16908 34660 16914 34672
rect 16908 34632 22094 34660
rect 16908 34620 16914 34632
rect 12986 34592 12992 34604
rect 12406 34564 12992 34592
rect 12986 34552 12992 34564
rect 13044 34552 13050 34604
rect 13538 34552 13544 34604
rect 13596 34592 13602 34604
rect 15562 34592 15568 34604
rect 13596 34564 15568 34592
rect 13596 34552 13602 34564
rect 15562 34552 15568 34564
rect 15620 34552 15626 34604
rect 15746 34552 15752 34604
rect 15804 34552 15810 34604
rect 15933 34595 15991 34601
rect 15933 34561 15945 34595
rect 15979 34592 15991 34595
rect 21634 34592 21640 34604
rect 15979 34564 21640 34592
rect 15979 34561 15991 34564
rect 15933 34555 15991 34561
rect 21634 34552 21640 34564
rect 21692 34552 21698 34604
rect 21726 34552 21732 34604
rect 21784 34592 21790 34604
rect 21821 34595 21879 34601
rect 21821 34592 21833 34595
rect 21784 34564 21833 34592
rect 21784 34552 21790 34564
rect 21821 34561 21833 34564
rect 21867 34561 21879 34595
rect 22066 34592 22094 34632
rect 29914 34620 29920 34672
rect 29972 34660 29978 34672
rect 34238 34660 34244 34672
rect 29972 34632 34244 34660
rect 29972 34620 29978 34632
rect 34238 34620 34244 34632
rect 34296 34660 34302 34672
rect 34296 34632 38700 34660
rect 34296 34620 34302 34632
rect 38672 34601 38700 34632
rect 38289 34595 38347 34601
rect 38289 34592 38301 34595
rect 22066 34564 38301 34592
rect 21821 34555 21879 34561
rect 38289 34561 38301 34564
rect 38335 34561 38347 34595
rect 38289 34555 38347 34561
rect 38381 34595 38439 34601
rect 38381 34561 38393 34595
rect 38427 34561 38439 34595
rect 38381 34555 38439 34561
rect 38657 34595 38715 34601
rect 38657 34561 38669 34595
rect 38703 34561 38715 34595
rect 38657 34555 38715 34561
rect 16666 34524 16672 34536
rect 7024 34496 16672 34524
rect 16666 34484 16672 34496
rect 16724 34524 16730 34536
rect 23017 34527 23075 34533
rect 23017 34524 23029 34527
rect 16724 34496 23029 34524
rect 16724 34484 16730 34496
rect 23017 34493 23029 34496
rect 23063 34524 23075 34527
rect 33134 34524 33140 34536
rect 23063 34496 33140 34524
rect 23063 34493 23075 34496
rect 23017 34487 23075 34493
rect 33134 34484 33140 34496
rect 33192 34484 33198 34536
rect 36170 34484 36176 34536
rect 36228 34524 36234 34536
rect 38396 34524 38424 34555
rect 36228 34496 38424 34524
rect 36228 34484 36234 34496
rect 38562 34484 38568 34536
rect 38620 34484 38626 34536
rect 13722 34416 13728 34468
rect 13780 34456 13786 34468
rect 19610 34456 19616 34468
rect 13780 34428 19616 34456
rect 13780 34416 13786 34428
rect 19610 34416 19616 34428
rect 19668 34416 19674 34468
rect 1104 34298 40848 34320
rect 1104 34246 1950 34298
rect 2002 34246 2014 34298
rect 2066 34246 2078 34298
rect 2130 34246 2142 34298
rect 2194 34246 2206 34298
rect 2258 34246 6950 34298
rect 7002 34246 7014 34298
rect 7066 34246 7078 34298
rect 7130 34246 7142 34298
rect 7194 34246 7206 34298
rect 7258 34246 11950 34298
rect 12002 34246 12014 34298
rect 12066 34246 12078 34298
rect 12130 34246 12142 34298
rect 12194 34246 12206 34298
rect 12258 34246 16950 34298
rect 17002 34246 17014 34298
rect 17066 34246 17078 34298
rect 17130 34246 17142 34298
rect 17194 34246 17206 34298
rect 17258 34246 21950 34298
rect 22002 34246 22014 34298
rect 22066 34246 22078 34298
rect 22130 34246 22142 34298
rect 22194 34246 22206 34298
rect 22258 34246 26950 34298
rect 27002 34246 27014 34298
rect 27066 34246 27078 34298
rect 27130 34246 27142 34298
rect 27194 34246 27206 34298
rect 27258 34246 31950 34298
rect 32002 34246 32014 34298
rect 32066 34246 32078 34298
rect 32130 34246 32142 34298
rect 32194 34246 32206 34298
rect 32258 34246 36950 34298
rect 37002 34246 37014 34298
rect 37066 34246 37078 34298
rect 37130 34246 37142 34298
rect 37194 34246 37206 34298
rect 37258 34246 40848 34298
rect 1104 34224 40848 34246
rect 14734 34144 14740 34196
rect 14792 34184 14798 34196
rect 25406 34184 25412 34196
rect 14792 34156 25412 34184
rect 14792 34144 14798 34156
rect 25406 34144 25412 34156
rect 25464 34144 25470 34196
rect 2409 34119 2467 34125
rect 2409 34085 2421 34119
rect 2455 34116 2467 34119
rect 2958 34116 2964 34128
rect 2455 34088 2964 34116
rect 2455 34085 2467 34088
rect 2409 34079 2467 34085
rect 2958 34076 2964 34088
rect 3016 34116 3022 34128
rect 5534 34116 5540 34128
rect 3016 34088 5540 34116
rect 3016 34076 3022 34088
rect 5534 34076 5540 34088
rect 5592 34076 5598 34128
rect 21818 34076 21824 34128
rect 21876 34116 21882 34128
rect 21876 34088 32628 34116
rect 21876 34076 21882 34088
rect 7466 34008 7472 34060
rect 7524 34048 7530 34060
rect 24854 34048 24860 34060
rect 7524 34020 24860 34048
rect 7524 34008 7530 34020
rect 24854 34008 24860 34020
rect 24912 34008 24918 34060
rect 1762 33940 1768 33992
rect 1820 33980 1826 33992
rect 2225 33983 2283 33989
rect 2225 33980 2237 33983
rect 1820 33952 2237 33980
rect 1820 33940 1826 33952
rect 2225 33949 2237 33952
rect 2271 33949 2283 33983
rect 2225 33943 2283 33949
rect 2501 33983 2559 33989
rect 2501 33949 2513 33983
rect 2547 33949 2559 33983
rect 2501 33943 2559 33949
rect 2516 33912 2544 33943
rect 14918 33940 14924 33992
rect 14976 33980 14982 33992
rect 15654 33980 15660 33992
rect 14976 33952 15660 33980
rect 14976 33940 14982 33952
rect 15654 33940 15660 33952
rect 15712 33980 15718 33992
rect 32600 33989 32628 34088
rect 17037 33983 17095 33989
rect 17037 33980 17049 33983
rect 15712 33952 17049 33980
rect 15712 33940 15718 33952
rect 17037 33949 17049 33952
rect 17083 33949 17095 33983
rect 17037 33943 17095 33949
rect 32585 33983 32643 33989
rect 32585 33949 32597 33983
rect 32631 33949 32643 33983
rect 32585 33943 32643 33949
rect 3510 33912 3516 33924
rect 2516 33884 3516 33912
rect 3510 33872 3516 33884
rect 3568 33912 3574 33924
rect 11698 33912 11704 33924
rect 3568 33884 11704 33912
rect 3568 33872 3574 33884
rect 11698 33872 11704 33884
rect 11756 33872 11762 33924
rect 13262 33872 13268 33924
rect 13320 33912 13326 33924
rect 17310 33912 17316 33924
rect 13320 33884 17316 33912
rect 13320 33872 13326 33884
rect 17310 33872 17316 33884
rect 17368 33872 17374 33924
rect 23566 33872 23572 33924
rect 23624 33912 23630 33924
rect 24118 33912 24124 33924
rect 23624 33884 24124 33912
rect 23624 33872 23630 33884
rect 24118 33872 24124 33884
rect 24176 33912 24182 33924
rect 33321 33915 33379 33921
rect 33321 33912 33333 33915
rect 24176 33884 33333 33912
rect 24176 33872 24182 33884
rect 33321 33881 33333 33884
rect 33367 33912 33379 33915
rect 36446 33912 36452 33924
rect 33367 33884 36452 33912
rect 33367 33881 33379 33884
rect 33321 33875 33379 33881
rect 36446 33872 36452 33884
rect 36504 33872 36510 33924
rect 2041 33847 2099 33853
rect 2041 33813 2053 33847
rect 2087 33844 2099 33847
rect 16114 33844 16120 33856
rect 2087 33816 16120 33844
rect 2087 33813 2099 33816
rect 2041 33807 2099 33813
rect 16114 33804 16120 33816
rect 16172 33804 16178 33856
rect 17221 33847 17279 33853
rect 17221 33813 17233 33847
rect 17267 33844 17279 33847
rect 27982 33844 27988 33856
rect 17267 33816 27988 33844
rect 17267 33813 17279 33816
rect 17221 33807 17279 33813
rect 27982 33804 27988 33816
rect 28040 33804 28046 33856
rect 1104 33754 40848 33776
rect 1104 33702 2610 33754
rect 2662 33702 2674 33754
rect 2726 33702 2738 33754
rect 2790 33702 2802 33754
rect 2854 33702 2866 33754
rect 2918 33702 7610 33754
rect 7662 33702 7674 33754
rect 7726 33702 7738 33754
rect 7790 33702 7802 33754
rect 7854 33702 7866 33754
rect 7918 33702 12610 33754
rect 12662 33702 12674 33754
rect 12726 33702 12738 33754
rect 12790 33702 12802 33754
rect 12854 33702 12866 33754
rect 12918 33702 17610 33754
rect 17662 33702 17674 33754
rect 17726 33702 17738 33754
rect 17790 33702 17802 33754
rect 17854 33702 17866 33754
rect 17918 33702 22610 33754
rect 22662 33702 22674 33754
rect 22726 33702 22738 33754
rect 22790 33702 22802 33754
rect 22854 33702 22866 33754
rect 22918 33702 27610 33754
rect 27662 33702 27674 33754
rect 27726 33702 27738 33754
rect 27790 33702 27802 33754
rect 27854 33702 27866 33754
rect 27918 33702 32610 33754
rect 32662 33702 32674 33754
rect 32726 33702 32738 33754
rect 32790 33702 32802 33754
rect 32854 33702 32866 33754
rect 32918 33702 37610 33754
rect 37662 33702 37674 33754
rect 37726 33702 37738 33754
rect 37790 33702 37802 33754
rect 37854 33702 37866 33754
rect 37918 33702 40848 33754
rect 1104 33680 40848 33702
rect 7374 33600 7380 33652
rect 7432 33640 7438 33652
rect 14826 33640 14832 33652
rect 7432 33612 14832 33640
rect 7432 33600 7438 33612
rect 14826 33600 14832 33612
rect 14884 33600 14890 33652
rect 14918 33600 14924 33652
rect 14976 33640 14982 33652
rect 14976 33612 15148 33640
rect 14976 33600 14982 33612
rect 6362 33532 6368 33584
rect 6420 33532 6426 33584
rect 6549 33507 6607 33513
rect 6549 33473 6561 33507
rect 6595 33504 6607 33507
rect 13538 33504 13544 33516
rect 6595 33476 13544 33504
rect 6595 33473 6607 33476
rect 6549 33467 6607 33473
rect 13538 33464 13544 33476
rect 13596 33464 13602 33516
rect 13722 33464 13728 33516
rect 13780 33464 13786 33516
rect 14182 33464 14188 33516
rect 14240 33464 14246 33516
rect 14645 33507 14703 33513
rect 14645 33473 14657 33507
rect 14691 33504 14703 33507
rect 14826 33504 14832 33516
rect 14691 33476 14832 33504
rect 14691 33473 14703 33476
rect 14645 33467 14703 33473
rect 14826 33464 14832 33476
rect 14884 33464 14890 33516
rect 15120 33513 15148 33612
rect 17494 33600 17500 33652
rect 17552 33640 17558 33652
rect 18417 33643 18475 33649
rect 18417 33640 18429 33643
rect 17552 33612 18429 33640
rect 17552 33600 17558 33612
rect 18417 33609 18429 33612
rect 18463 33609 18475 33643
rect 18585 33643 18643 33649
rect 18585 33640 18597 33643
rect 18417 33603 18475 33609
rect 18524 33612 18597 33640
rect 17310 33532 17316 33584
rect 17368 33572 17374 33584
rect 17773 33575 17831 33581
rect 17773 33572 17785 33575
rect 17368 33544 17785 33572
rect 17368 33532 17374 33544
rect 17773 33541 17785 33544
rect 17819 33541 17831 33575
rect 17773 33535 17831 33541
rect 18230 33532 18236 33584
rect 18288 33572 18294 33584
rect 18524 33572 18552 33612
rect 18585 33609 18597 33612
rect 18631 33640 18643 33643
rect 19242 33640 19248 33652
rect 18631 33612 19248 33640
rect 18631 33609 18643 33612
rect 18585 33603 18643 33609
rect 19242 33600 19248 33612
rect 19300 33600 19306 33652
rect 22376 33584 22428 33590
rect 18288 33544 18552 33572
rect 18785 33575 18843 33581
rect 18288 33532 18294 33544
rect 18785 33541 18797 33575
rect 18831 33572 18843 33575
rect 19334 33572 19340 33584
rect 18831 33544 19340 33572
rect 18831 33541 18843 33544
rect 18785 33535 18843 33541
rect 19334 33532 19340 33544
rect 19392 33572 19398 33584
rect 19886 33572 19892 33584
rect 19392 33544 19892 33572
rect 19392 33532 19398 33544
rect 19886 33532 19892 33544
rect 19944 33532 19950 33584
rect 24210 33572 24216 33584
rect 22376 33526 22428 33532
rect 23216 33544 24216 33572
rect 15105 33507 15163 33513
rect 15105 33473 15117 33507
rect 15151 33473 15163 33507
rect 15105 33467 15163 33473
rect 17681 33507 17739 33513
rect 17681 33473 17693 33507
rect 17727 33473 17739 33507
rect 17681 33467 17739 33473
rect 7374 33396 7380 33448
rect 7432 33436 7438 33448
rect 8386 33436 8392 33448
rect 7432 33408 8392 33436
rect 7432 33396 7438 33408
rect 8386 33396 8392 33408
rect 8444 33396 8450 33448
rect 14274 33396 14280 33448
rect 14332 33436 14338 33448
rect 15010 33436 15016 33448
rect 14332 33408 15016 33436
rect 14332 33396 14338 33408
rect 15010 33396 15016 33408
rect 15068 33396 15074 33448
rect 17696 33436 17724 33467
rect 17862 33464 17868 33516
rect 17920 33464 17926 33516
rect 23216 33513 23244 33544
rect 24210 33532 24216 33544
rect 24268 33532 24274 33584
rect 24854 33532 24860 33584
rect 24912 33532 24918 33584
rect 23201 33507 23259 33513
rect 23201 33473 23213 33507
rect 23247 33473 23259 33507
rect 23201 33467 23259 33473
rect 23290 33464 23296 33516
rect 23348 33504 23354 33516
rect 23477 33507 23535 33513
rect 23477 33504 23489 33507
rect 23348 33476 23489 33504
rect 23348 33464 23354 33476
rect 23477 33473 23489 33476
rect 23523 33473 23535 33507
rect 23477 33467 23535 33473
rect 25406 33464 25412 33516
rect 25464 33464 25470 33516
rect 25866 33464 25872 33516
rect 25924 33504 25930 33516
rect 26142 33504 26148 33516
rect 25924 33476 26148 33504
rect 25924 33464 25930 33476
rect 26142 33464 26148 33476
rect 26200 33464 26206 33516
rect 18874 33436 18880 33448
rect 17696 33408 18880 33436
rect 18874 33396 18880 33408
rect 18932 33396 18938 33448
rect 6362 33328 6368 33380
rect 6420 33368 6426 33380
rect 12986 33368 12992 33380
rect 6420 33340 12992 33368
rect 6420 33328 6426 33340
rect 12986 33328 12992 33340
rect 13044 33368 13050 33380
rect 15746 33368 15752 33380
rect 13044 33340 15752 33368
rect 13044 33328 13050 33340
rect 15746 33328 15752 33340
rect 15804 33328 15810 33380
rect 19978 33368 19984 33380
rect 15856 33340 19984 33368
rect 6641 33303 6699 33309
rect 6641 33269 6653 33303
rect 6687 33300 6699 33303
rect 13998 33300 14004 33312
rect 6687 33272 14004 33300
rect 6687 33269 6699 33272
rect 6641 33263 6699 33269
rect 13998 33260 14004 33272
rect 14056 33300 14062 33312
rect 14642 33300 14648 33312
rect 14056 33272 14648 33300
rect 14056 33260 14062 33272
rect 14642 33260 14648 33272
rect 14700 33260 14706 33312
rect 14826 33260 14832 33312
rect 14884 33300 14890 33312
rect 15856 33300 15884 33340
rect 19978 33328 19984 33340
rect 20036 33328 20042 33380
rect 14884 33272 15884 33300
rect 14884 33260 14890 33272
rect 18414 33260 18420 33312
rect 18472 33300 18478 33312
rect 18601 33303 18659 33309
rect 18601 33300 18613 33303
rect 18472 33272 18613 33300
rect 18472 33260 18478 33272
rect 18601 33269 18613 33272
rect 18647 33300 18659 33303
rect 18690 33300 18696 33312
rect 18647 33272 18696 33300
rect 18647 33269 18659 33272
rect 18601 33263 18659 33269
rect 18690 33260 18696 33272
rect 18748 33260 18754 33312
rect 1104 33210 40848 33232
rect 1104 33158 1950 33210
rect 2002 33158 2014 33210
rect 2066 33158 2078 33210
rect 2130 33158 2142 33210
rect 2194 33158 2206 33210
rect 2258 33158 6950 33210
rect 7002 33158 7014 33210
rect 7066 33158 7078 33210
rect 7130 33158 7142 33210
rect 7194 33158 7206 33210
rect 7258 33158 11950 33210
rect 12002 33158 12014 33210
rect 12066 33158 12078 33210
rect 12130 33158 12142 33210
rect 12194 33158 12206 33210
rect 12258 33158 16950 33210
rect 17002 33158 17014 33210
rect 17066 33158 17078 33210
rect 17130 33158 17142 33210
rect 17194 33158 17206 33210
rect 17258 33158 21950 33210
rect 22002 33158 22014 33210
rect 22066 33158 22078 33210
rect 22130 33158 22142 33210
rect 22194 33158 22206 33210
rect 22258 33158 26950 33210
rect 27002 33158 27014 33210
rect 27066 33158 27078 33210
rect 27130 33158 27142 33210
rect 27194 33158 27206 33210
rect 27258 33158 31950 33210
rect 32002 33158 32014 33210
rect 32066 33158 32078 33210
rect 32130 33158 32142 33210
rect 32194 33158 32206 33210
rect 32258 33158 36950 33210
rect 37002 33158 37014 33210
rect 37066 33158 37078 33210
rect 37130 33158 37142 33210
rect 37194 33158 37206 33210
rect 37258 33158 40848 33210
rect 1104 33136 40848 33158
rect 4890 33056 4896 33108
rect 4948 33096 4954 33108
rect 10226 33096 10232 33108
rect 4948 33068 10232 33096
rect 4948 33056 4954 33068
rect 10226 33056 10232 33068
rect 10284 33056 10290 33108
rect 13078 33056 13084 33108
rect 13136 33096 13142 33108
rect 14182 33096 14188 33108
rect 13136 33068 14188 33096
rect 13136 33056 13142 33068
rect 14182 33056 14188 33068
rect 14240 33056 14246 33108
rect 24486 33056 24492 33108
rect 24544 33096 24550 33108
rect 35986 33096 35992 33108
rect 24544 33068 35992 33096
rect 24544 33056 24550 33068
rect 35986 33056 35992 33068
rect 36044 33056 36050 33108
rect 36096 33068 37412 33096
rect 3142 32988 3148 33040
rect 3200 33028 3206 33040
rect 11514 33028 11520 33040
rect 3200 33000 11520 33028
rect 3200 32988 3206 33000
rect 11514 32988 11520 33000
rect 11572 32988 11578 33040
rect 13538 32988 13544 33040
rect 13596 33028 13602 33040
rect 13722 33028 13728 33040
rect 13596 33000 13728 33028
rect 13596 32988 13602 33000
rect 13722 32988 13728 33000
rect 13780 32988 13786 33040
rect 15930 32988 15936 33040
rect 15988 33028 15994 33040
rect 16577 33031 16635 33037
rect 16577 33028 16589 33031
rect 15988 33000 16589 33028
rect 15988 32988 15994 33000
rect 16577 32997 16589 33000
rect 16623 32997 16635 33031
rect 16577 32991 16635 32997
rect 30374 32988 30380 33040
rect 30432 33028 30438 33040
rect 31478 33028 31484 33040
rect 30432 33000 31484 33028
rect 30432 32988 30438 33000
rect 31478 32988 31484 33000
rect 31536 33028 31542 33040
rect 36096 33028 36124 33068
rect 31536 33000 36124 33028
rect 37277 33031 37335 33037
rect 31536 32988 31542 33000
rect 37277 32997 37289 33031
rect 37323 32997 37335 33031
rect 37277 32991 37335 32997
rect 5718 32920 5724 32972
rect 5776 32960 5782 32972
rect 11606 32960 11612 32972
rect 5776 32932 11612 32960
rect 5776 32920 5782 32932
rect 11606 32920 11612 32932
rect 11664 32920 11670 32972
rect 13814 32920 13820 32972
rect 13872 32960 13878 32972
rect 18046 32960 18052 32972
rect 13872 32932 18052 32960
rect 13872 32920 13878 32932
rect 18046 32920 18052 32932
rect 18104 32920 18110 32972
rect 37292 32960 37320 32991
rect 33336 32932 37320 32960
rect 37384 32946 37412 33068
rect 39209 33031 39267 33037
rect 39209 33028 39221 33031
rect 38672 33000 39221 33028
rect 38672 32969 38700 33000
rect 39209 32997 39221 33000
rect 39255 32997 39267 33031
rect 39209 32991 39267 32997
rect 38657 32963 38715 32969
rect 17402 32852 17408 32904
rect 17460 32892 17466 32904
rect 33226 32892 33232 32904
rect 17460 32864 33232 32892
rect 17460 32852 17466 32864
rect 33226 32852 33232 32864
rect 33284 32852 33290 32904
rect 16761 32827 16819 32833
rect 16761 32793 16773 32827
rect 16807 32824 16819 32827
rect 16850 32824 16856 32836
rect 16807 32796 16856 32824
rect 16807 32793 16819 32796
rect 16761 32787 16819 32793
rect 16850 32784 16856 32796
rect 16908 32824 16914 32836
rect 33336 32824 33364 32932
rect 38657 32929 38669 32963
rect 38703 32929 38715 32963
rect 38657 32923 38715 32929
rect 33505 32895 33563 32901
rect 33505 32861 33517 32895
rect 33551 32892 33563 32895
rect 33551 32864 35894 32892
rect 33551 32861 33563 32864
rect 33505 32855 33563 32861
rect 16908 32796 33364 32824
rect 16908 32784 16914 32796
rect 35866 32756 35894 32864
rect 36538 32852 36544 32904
rect 36596 32892 36602 32904
rect 37461 32895 37519 32901
rect 37461 32892 37473 32895
rect 36596 32864 37473 32892
rect 36596 32852 36602 32864
rect 37461 32861 37473 32864
rect 37507 32861 37519 32895
rect 37461 32855 37519 32861
rect 38105 32895 38163 32901
rect 38105 32861 38117 32895
rect 38151 32861 38163 32895
rect 38105 32855 38163 32861
rect 35986 32784 35992 32836
rect 36044 32824 36050 32836
rect 38120 32824 38148 32855
rect 38194 32852 38200 32904
rect 38252 32892 38258 32904
rect 38749 32895 38807 32901
rect 38749 32892 38761 32895
rect 38252 32864 38761 32892
rect 38252 32852 38258 32864
rect 38749 32861 38761 32864
rect 38795 32861 38807 32895
rect 38749 32855 38807 32861
rect 36044 32796 38148 32824
rect 36044 32784 36050 32796
rect 38194 32756 38200 32768
rect 35866 32728 38200 32756
rect 38194 32716 38200 32728
rect 38252 32716 38258 32768
rect 1104 32666 40848 32688
rect 1104 32614 2610 32666
rect 2662 32614 2674 32666
rect 2726 32614 2738 32666
rect 2790 32614 2802 32666
rect 2854 32614 2866 32666
rect 2918 32614 7610 32666
rect 7662 32614 7674 32666
rect 7726 32614 7738 32666
rect 7790 32614 7802 32666
rect 7854 32614 7866 32666
rect 7918 32614 12610 32666
rect 12662 32614 12674 32666
rect 12726 32614 12738 32666
rect 12790 32614 12802 32666
rect 12854 32614 12866 32666
rect 12918 32614 17610 32666
rect 17662 32614 17674 32666
rect 17726 32614 17738 32666
rect 17790 32614 17802 32666
rect 17854 32614 17866 32666
rect 17918 32614 22610 32666
rect 22662 32614 22674 32666
rect 22726 32614 22738 32666
rect 22790 32614 22802 32666
rect 22854 32614 22866 32666
rect 22918 32614 27610 32666
rect 27662 32614 27674 32666
rect 27726 32614 27738 32666
rect 27790 32614 27802 32666
rect 27854 32614 27866 32666
rect 27918 32614 32610 32666
rect 32662 32614 32674 32666
rect 32726 32614 32738 32666
rect 32790 32614 32802 32666
rect 32854 32614 32866 32666
rect 32918 32614 37610 32666
rect 37662 32614 37674 32666
rect 37726 32614 37738 32666
rect 37790 32614 37802 32666
rect 37854 32614 37866 32666
rect 37918 32614 40848 32666
rect 1104 32592 40848 32614
rect 6917 32555 6975 32561
rect 6917 32521 6929 32555
rect 6963 32552 6975 32555
rect 9766 32552 9772 32564
rect 6963 32524 9772 32552
rect 6963 32521 6975 32524
rect 6917 32515 6975 32521
rect 9766 32512 9772 32524
rect 9824 32512 9830 32564
rect 16022 32512 16028 32564
rect 16080 32552 16086 32564
rect 19058 32552 19064 32564
rect 16080 32524 19064 32552
rect 16080 32512 16086 32524
rect 6086 32444 6092 32496
rect 6144 32484 6150 32496
rect 6144 32456 6776 32484
rect 6144 32444 6150 32456
rect 6748 32428 6776 32456
rect 11422 32444 11428 32496
rect 11480 32484 11486 32496
rect 16942 32484 16948 32496
rect 11480 32456 16948 32484
rect 11480 32444 11486 32456
rect 16942 32444 16948 32456
rect 17000 32444 17006 32496
rect 17052 32493 17080 32524
rect 19058 32512 19064 32524
rect 19116 32512 19122 32564
rect 17037 32487 17095 32493
rect 17037 32453 17049 32487
rect 17083 32453 17095 32487
rect 17037 32447 17095 32453
rect 17126 32444 17132 32496
rect 17184 32484 17190 32496
rect 29273 32487 29331 32493
rect 17184 32456 29224 32484
rect 17184 32444 17190 32456
rect 5994 32376 6000 32428
rect 6052 32416 6058 32428
rect 6362 32416 6368 32428
rect 6052 32388 6368 32416
rect 6052 32376 6058 32388
rect 6362 32376 6368 32388
rect 6420 32376 6426 32428
rect 6638 32376 6644 32428
rect 6696 32376 6702 32428
rect 6730 32376 6736 32428
rect 6788 32376 6794 32428
rect 16853 32419 16911 32425
rect 16853 32385 16865 32419
rect 16899 32416 16911 32419
rect 19889 32419 19947 32425
rect 16899 32388 19288 32416
rect 16899 32385 16911 32388
rect 16853 32379 16911 32385
rect 19260 32360 19288 32388
rect 19889 32385 19901 32419
rect 19935 32385 19947 32419
rect 19889 32379 19947 32385
rect 19981 32419 20039 32425
rect 19981 32385 19993 32419
rect 20027 32385 20039 32419
rect 19981 32379 20039 32385
rect 6454 32308 6460 32360
rect 6512 32308 6518 32360
rect 19242 32308 19248 32360
rect 19300 32348 19306 32360
rect 19904 32348 19932 32379
rect 19300 32320 19932 32348
rect 19300 32308 19306 32320
rect 17221 32283 17279 32289
rect 17221 32249 17233 32283
rect 17267 32280 17279 32283
rect 18966 32280 18972 32292
rect 17267 32252 18972 32280
rect 17267 32249 17279 32252
rect 17221 32243 17279 32249
rect 18966 32240 18972 32252
rect 19024 32240 19030 32292
rect 19058 32240 19064 32292
rect 19116 32280 19122 32292
rect 19996 32280 20024 32379
rect 28626 32376 28632 32428
rect 28684 32376 28690 32428
rect 28810 32376 28816 32428
rect 28868 32376 28874 32428
rect 28905 32419 28963 32425
rect 28905 32385 28917 32419
rect 28951 32385 28963 32419
rect 28905 32379 28963 32385
rect 20165 32351 20223 32357
rect 20165 32317 20177 32351
rect 20211 32348 20223 32351
rect 24302 32348 24308 32360
rect 20211 32320 24308 32348
rect 20211 32317 20223 32320
rect 20165 32311 20223 32317
rect 24302 32308 24308 32320
rect 24360 32308 24366 32360
rect 28718 32308 28724 32360
rect 28776 32348 28782 32360
rect 28920 32348 28948 32379
rect 28994 32376 29000 32428
rect 29052 32416 29058 32428
rect 29196 32416 29224 32456
rect 29273 32453 29285 32487
rect 29319 32484 29331 32487
rect 30926 32484 30932 32496
rect 29319 32456 30932 32484
rect 29319 32453 29331 32456
rect 29273 32447 29331 32453
rect 30926 32444 30932 32456
rect 30984 32444 30990 32496
rect 30466 32416 30472 32428
rect 29052 32388 29097 32416
rect 29196 32388 30472 32416
rect 29052 32376 29058 32388
rect 30466 32376 30472 32388
rect 30524 32376 30530 32428
rect 28776 32320 28948 32348
rect 28776 32308 28782 32320
rect 19116 32252 20024 32280
rect 19116 32240 19122 32252
rect 18046 32172 18052 32224
rect 18104 32212 18110 32224
rect 18322 32212 18328 32224
rect 18104 32184 18328 32212
rect 18104 32172 18110 32184
rect 18322 32172 18328 32184
rect 18380 32172 18386 32224
rect 1104 32122 40848 32144
rect 1104 32070 1950 32122
rect 2002 32070 2014 32122
rect 2066 32070 2078 32122
rect 2130 32070 2142 32122
rect 2194 32070 2206 32122
rect 2258 32070 6950 32122
rect 7002 32070 7014 32122
rect 7066 32070 7078 32122
rect 7130 32070 7142 32122
rect 7194 32070 7206 32122
rect 7258 32070 11950 32122
rect 12002 32070 12014 32122
rect 12066 32070 12078 32122
rect 12130 32070 12142 32122
rect 12194 32070 12206 32122
rect 12258 32070 16950 32122
rect 17002 32070 17014 32122
rect 17066 32070 17078 32122
rect 17130 32070 17142 32122
rect 17194 32070 17206 32122
rect 17258 32070 21950 32122
rect 22002 32070 22014 32122
rect 22066 32070 22078 32122
rect 22130 32070 22142 32122
rect 22194 32070 22206 32122
rect 22258 32070 26950 32122
rect 27002 32070 27014 32122
rect 27066 32070 27078 32122
rect 27130 32070 27142 32122
rect 27194 32070 27206 32122
rect 27258 32070 31950 32122
rect 32002 32070 32014 32122
rect 32066 32070 32078 32122
rect 32130 32070 32142 32122
rect 32194 32070 32206 32122
rect 32258 32070 36950 32122
rect 37002 32070 37014 32122
rect 37066 32070 37078 32122
rect 37130 32070 37142 32122
rect 37194 32070 37206 32122
rect 37258 32070 40848 32122
rect 1104 32048 40848 32070
rect 18322 31968 18328 32020
rect 18380 32008 18386 32020
rect 18380 31980 18644 32008
rect 18380 31968 18386 31980
rect 16390 31900 16396 31952
rect 16448 31940 16454 31952
rect 16758 31940 16764 31952
rect 16448 31912 16764 31940
rect 16448 31900 16454 31912
rect 16758 31900 16764 31912
rect 16816 31900 16822 31952
rect 16945 31943 17003 31949
rect 16945 31909 16957 31943
rect 16991 31940 17003 31943
rect 17310 31940 17316 31952
rect 16991 31912 17316 31940
rect 16991 31909 17003 31912
rect 16945 31903 17003 31909
rect 17310 31900 17316 31912
rect 17368 31900 17374 31952
rect 18616 31949 18644 31980
rect 18509 31943 18567 31949
rect 18509 31909 18521 31943
rect 18555 31909 18567 31943
rect 18509 31903 18567 31909
rect 18601 31943 18659 31949
rect 18601 31909 18613 31943
rect 18647 31909 18659 31943
rect 18601 31903 18659 31909
rect 7374 31832 7380 31884
rect 7432 31832 7438 31884
rect 9306 31832 9312 31884
rect 9364 31872 9370 31884
rect 9677 31875 9735 31881
rect 9677 31872 9689 31875
rect 9364 31844 9689 31872
rect 9364 31832 9370 31844
rect 9677 31841 9689 31844
rect 9723 31872 9735 31875
rect 10226 31872 10232 31884
rect 9723 31844 10232 31872
rect 9723 31841 9735 31844
rect 9677 31835 9735 31841
rect 10226 31832 10232 31844
rect 10284 31832 10290 31884
rect 18524 31872 18552 31903
rect 18690 31900 18696 31952
rect 18748 31940 18754 31952
rect 19334 31940 19340 31952
rect 18748 31912 19340 31940
rect 18748 31900 18754 31912
rect 19334 31900 19340 31912
rect 19392 31900 19398 31952
rect 18874 31872 18880 31884
rect 18524 31844 18880 31872
rect 18874 31832 18880 31844
rect 18932 31832 18938 31884
rect 24578 31872 24584 31884
rect 19306 31844 24584 31872
rect 1394 31764 1400 31816
rect 1452 31764 1458 31816
rect 1670 31764 1676 31816
rect 1728 31764 1734 31816
rect 7392 31668 7420 31832
rect 9030 31764 9036 31816
rect 9088 31764 9094 31816
rect 17402 31764 17408 31816
rect 17460 31764 17466 31816
rect 18969 31739 19027 31745
rect 18969 31705 18981 31739
rect 19015 31736 19027 31739
rect 19306 31736 19334 31844
rect 24578 31832 24584 31844
rect 24636 31832 24642 31884
rect 30558 31832 30564 31884
rect 30616 31872 30622 31884
rect 30616 31844 31156 31872
rect 30616 31832 30622 31844
rect 31128 31816 31156 31844
rect 27338 31764 27344 31816
rect 27396 31804 27402 31816
rect 30929 31807 30987 31813
rect 30929 31804 30941 31807
rect 27396 31776 30941 31804
rect 27396 31764 27402 31776
rect 30929 31773 30941 31776
rect 30975 31773 30987 31807
rect 30929 31767 30987 31773
rect 31110 31764 31116 31816
rect 31168 31764 31174 31816
rect 31297 31807 31355 31813
rect 31297 31773 31309 31807
rect 31343 31804 31355 31807
rect 32490 31804 32496 31816
rect 31343 31776 32496 31804
rect 31343 31773 31355 31776
rect 31297 31767 31355 31773
rect 32490 31764 32496 31776
rect 32548 31804 32554 31816
rect 34054 31804 34060 31816
rect 32548 31776 34060 31804
rect 32548 31764 32554 31776
rect 34054 31764 34060 31776
rect 34112 31764 34118 31816
rect 19015 31708 19334 31736
rect 19015 31705 19027 31708
rect 18969 31699 19027 31705
rect 7466 31668 7472 31680
rect 7392 31640 7472 31668
rect 7466 31628 7472 31640
rect 7524 31628 7530 31680
rect 16850 31628 16856 31680
rect 16908 31668 16914 31680
rect 18984 31668 19012 31699
rect 16908 31640 19012 31668
rect 16908 31628 16914 31640
rect 1104 31578 40848 31600
rect 1104 31526 2610 31578
rect 2662 31526 2674 31578
rect 2726 31526 2738 31578
rect 2790 31526 2802 31578
rect 2854 31526 2866 31578
rect 2918 31526 7610 31578
rect 7662 31526 7674 31578
rect 7726 31526 7738 31578
rect 7790 31526 7802 31578
rect 7854 31526 7866 31578
rect 7918 31526 12610 31578
rect 12662 31526 12674 31578
rect 12726 31526 12738 31578
rect 12790 31526 12802 31578
rect 12854 31526 12866 31578
rect 12918 31526 17610 31578
rect 17662 31526 17674 31578
rect 17726 31526 17738 31578
rect 17790 31526 17802 31578
rect 17854 31526 17866 31578
rect 17918 31526 22610 31578
rect 22662 31526 22674 31578
rect 22726 31526 22738 31578
rect 22790 31526 22802 31578
rect 22854 31526 22866 31578
rect 22918 31526 27610 31578
rect 27662 31526 27674 31578
rect 27726 31526 27738 31578
rect 27790 31526 27802 31578
rect 27854 31526 27866 31578
rect 27918 31526 32610 31578
rect 32662 31526 32674 31578
rect 32726 31526 32738 31578
rect 32790 31526 32802 31578
rect 32854 31526 32866 31578
rect 32918 31526 37610 31578
rect 37662 31526 37674 31578
rect 37726 31526 37738 31578
rect 37790 31526 37802 31578
rect 37854 31526 37866 31578
rect 37918 31526 40848 31578
rect 1104 31504 40848 31526
rect 16666 31424 16672 31476
rect 16724 31464 16730 31476
rect 16724 31436 17080 31464
rect 16724 31424 16730 31436
rect 17052 31405 17080 31436
rect 16837 31399 16895 31405
rect 16837 31365 16849 31399
rect 16883 31396 16895 31399
rect 17037 31399 17095 31405
rect 16883 31368 16988 31396
rect 16883 31365 16895 31368
rect 16837 31359 16895 31365
rect 16960 31328 16988 31368
rect 17037 31365 17049 31399
rect 17083 31365 17095 31399
rect 17037 31359 17095 31365
rect 17402 31328 17408 31340
rect 16960 31300 17408 31328
rect 17402 31288 17408 31300
rect 17460 31288 17466 31340
rect 18322 31288 18328 31340
rect 18380 31328 18386 31340
rect 31570 31328 31576 31340
rect 18380 31300 31576 31328
rect 18380 31288 18386 31300
rect 31570 31288 31576 31300
rect 31628 31288 31634 31340
rect 40494 31288 40500 31340
rect 40552 31288 40558 31340
rect 10226 31220 10232 31272
rect 10284 31260 10290 31272
rect 24578 31260 24584 31272
rect 10284 31232 24584 31260
rect 10284 31220 10290 31232
rect 24578 31220 24584 31232
rect 24636 31220 24642 31272
rect 24762 31220 24768 31272
rect 24820 31260 24826 31272
rect 33778 31260 33784 31272
rect 24820 31232 33784 31260
rect 24820 31220 24826 31232
rect 33778 31220 33784 31232
rect 33836 31220 33842 31272
rect 38286 31220 38292 31272
rect 38344 31260 38350 31272
rect 39669 31263 39727 31269
rect 39669 31260 39681 31263
rect 38344 31232 39681 31260
rect 38344 31220 38350 31232
rect 39669 31229 39681 31232
rect 39715 31229 39727 31263
rect 39669 31223 39727 31229
rect 8294 31152 8300 31204
rect 8352 31192 8358 31204
rect 24946 31192 24952 31204
rect 8352 31164 24952 31192
rect 8352 31152 8358 31164
rect 24946 31152 24952 31164
rect 25004 31152 25010 31204
rect 15930 31084 15936 31136
rect 15988 31124 15994 31136
rect 16669 31127 16727 31133
rect 16669 31124 16681 31127
rect 15988 31096 16681 31124
rect 15988 31084 15994 31096
rect 16669 31093 16681 31096
rect 16715 31093 16727 31127
rect 16669 31087 16727 31093
rect 16853 31127 16911 31133
rect 16853 31093 16865 31127
rect 16899 31124 16911 31127
rect 18506 31124 18512 31136
rect 16899 31096 18512 31124
rect 16899 31093 16911 31096
rect 16853 31087 16911 31093
rect 18506 31084 18512 31096
rect 18564 31084 18570 31136
rect 31202 31084 31208 31136
rect 31260 31124 31266 31136
rect 31386 31124 31392 31136
rect 31260 31096 31392 31124
rect 31260 31084 31266 31096
rect 31386 31084 31392 31096
rect 31444 31084 31450 31136
rect 1104 31034 40848 31056
rect 1104 30982 1950 31034
rect 2002 30982 2014 31034
rect 2066 30982 2078 31034
rect 2130 30982 2142 31034
rect 2194 30982 2206 31034
rect 2258 30982 6950 31034
rect 7002 30982 7014 31034
rect 7066 30982 7078 31034
rect 7130 30982 7142 31034
rect 7194 30982 7206 31034
rect 7258 30982 11950 31034
rect 12002 30982 12014 31034
rect 12066 30982 12078 31034
rect 12130 30982 12142 31034
rect 12194 30982 12206 31034
rect 12258 30982 16950 31034
rect 17002 30982 17014 31034
rect 17066 30982 17078 31034
rect 17130 30982 17142 31034
rect 17194 30982 17206 31034
rect 17258 30982 21950 31034
rect 22002 30982 22014 31034
rect 22066 30982 22078 31034
rect 22130 30982 22142 31034
rect 22194 30982 22206 31034
rect 22258 30982 26950 31034
rect 27002 30982 27014 31034
rect 27066 30982 27078 31034
rect 27130 30982 27142 31034
rect 27194 30982 27206 31034
rect 27258 30982 31950 31034
rect 32002 30982 32014 31034
rect 32066 30982 32078 31034
rect 32130 30982 32142 31034
rect 32194 30982 32206 31034
rect 32258 30982 36950 31034
rect 37002 30982 37014 31034
rect 37066 30982 37078 31034
rect 37130 30982 37142 31034
rect 37194 30982 37206 31034
rect 37258 30982 40848 31034
rect 1104 30960 40848 30982
rect 16114 30880 16120 30932
rect 16172 30920 16178 30932
rect 16482 30920 16488 30932
rect 16172 30892 16488 30920
rect 16172 30880 16178 30892
rect 16482 30880 16488 30892
rect 16540 30880 16546 30932
rect 17862 30880 17868 30932
rect 17920 30920 17926 30932
rect 24762 30920 24768 30932
rect 17920 30892 24768 30920
rect 17920 30880 17926 30892
rect 24762 30880 24768 30892
rect 24820 30880 24826 30932
rect 35986 30880 35992 30932
rect 36044 30920 36050 30932
rect 36354 30920 36360 30932
rect 36044 30892 36360 30920
rect 36044 30880 36050 30892
rect 36354 30880 36360 30892
rect 36412 30880 36418 30932
rect 36722 30812 36728 30864
rect 36780 30852 36786 30864
rect 36817 30855 36875 30861
rect 36817 30852 36829 30855
rect 36780 30824 36829 30852
rect 36780 30812 36786 30824
rect 36817 30821 36829 30824
rect 36863 30821 36875 30855
rect 36817 30815 36875 30821
rect 2498 30784 2504 30796
rect 2332 30756 2504 30784
rect 1854 30676 1860 30728
rect 1912 30716 1918 30728
rect 2332 30725 2360 30756
rect 2498 30744 2504 30756
rect 2556 30744 2562 30796
rect 17954 30744 17960 30796
rect 18012 30784 18018 30796
rect 18230 30784 18236 30796
rect 18012 30756 18236 30784
rect 18012 30744 18018 30756
rect 18230 30744 18236 30756
rect 18288 30744 18294 30796
rect 2041 30719 2099 30725
rect 2041 30716 2053 30719
rect 1912 30688 2053 30716
rect 1912 30676 1918 30688
rect 2041 30685 2053 30688
rect 2087 30685 2099 30719
rect 2041 30679 2099 30685
rect 2133 30719 2191 30725
rect 2133 30685 2145 30719
rect 2179 30685 2191 30719
rect 2133 30679 2191 30685
rect 2317 30719 2375 30725
rect 2317 30685 2329 30719
rect 2363 30685 2375 30719
rect 2317 30679 2375 30685
rect 2409 30719 2467 30725
rect 2409 30685 2421 30719
rect 2455 30716 2467 30719
rect 3510 30716 3516 30728
rect 2455 30688 3516 30716
rect 2455 30685 2467 30688
rect 2409 30679 2467 30685
rect 1486 30608 1492 30660
rect 1544 30648 1550 30660
rect 2148 30648 2176 30679
rect 3510 30676 3516 30688
rect 3568 30716 3574 30728
rect 9858 30716 9864 30728
rect 3568 30688 9864 30716
rect 3568 30676 3574 30688
rect 9858 30676 9864 30688
rect 9916 30676 9922 30728
rect 27430 30676 27436 30728
rect 27488 30716 27494 30728
rect 36387 30719 36445 30725
rect 36387 30716 36399 30719
rect 27488 30688 36399 30716
rect 27488 30676 27494 30688
rect 36387 30685 36399 30688
rect 36433 30685 36445 30719
rect 36387 30679 36445 30685
rect 36814 30676 36820 30728
rect 36872 30716 36878 30728
rect 36909 30719 36967 30725
rect 36909 30716 36921 30719
rect 36872 30688 36921 30716
rect 36872 30676 36878 30688
rect 36909 30685 36921 30688
rect 36955 30685 36967 30719
rect 36909 30679 36967 30685
rect 1544 30620 2176 30648
rect 1544 30608 1550 30620
rect 1857 30583 1915 30589
rect 1857 30549 1869 30583
rect 1903 30580 1915 30583
rect 13170 30580 13176 30592
rect 1903 30552 13176 30580
rect 1903 30549 1915 30552
rect 1857 30543 1915 30549
rect 13170 30540 13176 30552
rect 13228 30540 13234 30592
rect 36262 30540 36268 30592
rect 36320 30540 36326 30592
rect 36446 30540 36452 30592
rect 36504 30540 36510 30592
rect 1104 30490 40848 30512
rect 1104 30438 2610 30490
rect 2662 30438 2674 30490
rect 2726 30438 2738 30490
rect 2790 30438 2802 30490
rect 2854 30438 2866 30490
rect 2918 30438 7610 30490
rect 7662 30438 7674 30490
rect 7726 30438 7738 30490
rect 7790 30438 7802 30490
rect 7854 30438 7866 30490
rect 7918 30438 12610 30490
rect 12662 30438 12674 30490
rect 12726 30438 12738 30490
rect 12790 30438 12802 30490
rect 12854 30438 12866 30490
rect 12918 30438 17610 30490
rect 17662 30438 17674 30490
rect 17726 30438 17738 30490
rect 17790 30438 17802 30490
rect 17854 30438 17866 30490
rect 17918 30438 22610 30490
rect 22662 30438 22674 30490
rect 22726 30438 22738 30490
rect 22790 30438 22802 30490
rect 22854 30438 22866 30490
rect 22918 30438 27610 30490
rect 27662 30438 27674 30490
rect 27726 30438 27738 30490
rect 27790 30438 27802 30490
rect 27854 30438 27866 30490
rect 27918 30438 32610 30490
rect 32662 30438 32674 30490
rect 32726 30438 32738 30490
rect 32790 30438 32802 30490
rect 32854 30438 32866 30490
rect 32918 30438 37610 30490
rect 37662 30438 37674 30490
rect 37726 30438 37738 30490
rect 37790 30438 37802 30490
rect 37854 30438 37866 30490
rect 37918 30438 40848 30490
rect 1104 30416 40848 30438
rect 9122 30268 9128 30320
rect 9180 30308 9186 30320
rect 35434 30308 35440 30320
rect 9180 30280 35440 30308
rect 9180 30268 9186 30280
rect 35434 30268 35440 30280
rect 35492 30268 35498 30320
rect 16666 30200 16672 30252
rect 16724 30240 16730 30252
rect 31205 30243 31263 30249
rect 31205 30240 31217 30243
rect 16724 30212 31217 30240
rect 16724 30200 16730 30212
rect 31205 30209 31217 30212
rect 31251 30240 31263 30243
rect 33410 30240 33416 30252
rect 31251 30212 33416 30240
rect 31251 30209 31263 30212
rect 31205 30203 31263 30209
rect 33410 30200 33416 30212
rect 33468 30200 33474 30252
rect 8846 30132 8852 30184
rect 8904 30172 8910 30184
rect 8904 30144 30328 30172
rect 8904 30132 8910 30144
rect 11330 30064 11336 30116
rect 11388 30104 11394 30116
rect 30098 30104 30104 30116
rect 11388 30076 30104 30104
rect 11388 30064 11394 30076
rect 30098 30064 30104 30076
rect 30156 30064 30162 30116
rect 30300 30104 30328 30144
rect 30374 30132 30380 30184
rect 30432 30132 30438 30184
rect 30466 30132 30472 30184
rect 30524 30132 30530 30184
rect 31297 30175 31355 30181
rect 31297 30141 31309 30175
rect 31343 30141 31355 30175
rect 31297 30135 31355 30141
rect 31202 30104 31208 30116
rect 30300 30076 31208 30104
rect 31202 30064 31208 30076
rect 31260 30104 31266 30116
rect 31312 30104 31340 30135
rect 31260 30076 31340 30104
rect 31260 30064 31266 30076
rect 15010 29996 15016 30048
rect 15068 30036 15074 30048
rect 36078 30036 36084 30048
rect 15068 30008 36084 30036
rect 15068 29996 15074 30008
rect 36078 29996 36084 30008
rect 36136 29996 36142 30048
rect 1104 29946 40848 29968
rect 1104 29894 1950 29946
rect 2002 29894 2014 29946
rect 2066 29894 2078 29946
rect 2130 29894 2142 29946
rect 2194 29894 2206 29946
rect 2258 29894 6950 29946
rect 7002 29894 7014 29946
rect 7066 29894 7078 29946
rect 7130 29894 7142 29946
rect 7194 29894 7206 29946
rect 7258 29894 11950 29946
rect 12002 29894 12014 29946
rect 12066 29894 12078 29946
rect 12130 29894 12142 29946
rect 12194 29894 12206 29946
rect 12258 29894 16950 29946
rect 17002 29894 17014 29946
rect 17066 29894 17078 29946
rect 17130 29894 17142 29946
rect 17194 29894 17206 29946
rect 17258 29894 21950 29946
rect 22002 29894 22014 29946
rect 22066 29894 22078 29946
rect 22130 29894 22142 29946
rect 22194 29894 22206 29946
rect 22258 29894 26950 29946
rect 27002 29894 27014 29946
rect 27066 29894 27078 29946
rect 27130 29894 27142 29946
rect 27194 29894 27206 29946
rect 27258 29894 31950 29946
rect 32002 29894 32014 29946
rect 32066 29894 32078 29946
rect 32130 29894 32142 29946
rect 32194 29894 32206 29946
rect 32258 29894 36950 29946
rect 37002 29894 37014 29946
rect 37066 29894 37078 29946
rect 37130 29894 37142 29946
rect 37194 29894 37206 29946
rect 37258 29894 40848 29946
rect 1104 29872 40848 29894
rect 9214 29792 9220 29844
rect 9272 29832 9278 29844
rect 23566 29832 23572 29844
rect 9272 29804 23572 29832
rect 9272 29792 9278 29804
rect 23566 29792 23572 29804
rect 23624 29792 23630 29844
rect 35434 29792 35440 29844
rect 35492 29832 35498 29844
rect 35621 29835 35679 29841
rect 35621 29832 35633 29835
rect 35492 29804 35633 29832
rect 35492 29792 35498 29804
rect 35621 29801 35633 29804
rect 35667 29801 35679 29835
rect 35621 29795 35679 29801
rect 36170 29792 36176 29844
rect 36228 29832 36234 29844
rect 36449 29835 36507 29841
rect 36449 29832 36461 29835
rect 36228 29804 36461 29832
rect 36228 29792 36234 29804
rect 36449 29801 36461 29804
rect 36495 29801 36507 29835
rect 36449 29795 36507 29801
rect 30926 29764 30932 29776
rect 20916 29736 30932 29764
rect 20916 29708 20944 29736
rect 30926 29724 30932 29736
rect 30984 29724 30990 29776
rect 17402 29656 17408 29708
rect 17460 29696 17466 29708
rect 18322 29696 18328 29708
rect 17460 29668 18328 29696
rect 17460 29656 17466 29668
rect 18322 29656 18328 29668
rect 18380 29656 18386 29708
rect 20898 29656 20904 29708
rect 20956 29656 20962 29708
rect 22462 29696 22468 29708
rect 22020 29668 22468 29696
rect 21634 29588 21640 29640
rect 21692 29588 21698 29640
rect 21729 29631 21787 29637
rect 21729 29597 21741 29631
rect 21775 29628 21787 29631
rect 21818 29628 21824 29640
rect 21775 29600 21824 29628
rect 21775 29597 21787 29600
rect 21729 29591 21787 29597
rect 21818 29588 21824 29600
rect 21876 29588 21882 29640
rect 22020 29637 22048 29668
rect 22462 29656 22468 29668
rect 22520 29696 22526 29708
rect 26050 29696 26056 29708
rect 22520 29668 26056 29696
rect 22520 29656 22526 29668
rect 26050 29656 26056 29668
rect 26108 29656 26114 29708
rect 28626 29656 28632 29708
rect 28684 29696 28690 29708
rect 32585 29699 32643 29705
rect 32585 29696 32597 29699
rect 28684 29668 32597 29696
rect 28684 29656 28690 29668
rect 32585 29665 32597 29668
rect 32631 29696 32643 29699
rect 38930 29696 38936 29708
rect 32631 29668 38936 29696
rect 32631 29665 32643 29668
rect 32585 29659 32643 29665
rect 38930 29656 38936 29668
rect 38988 29656 38994 29708
rect 22005 29631 22063 29637
rect 22005 29597 22017 29631
rect 22051 29597 22063 29631
rect 22005 29591 22063 29597
rect 22097 29631 22155 29637
rect 22097 29597 22109 29631
rect 22143 29628 22155 29631
rect 23198 29628 23204 29640
rect 22143 29600 23204 29628
rect 22143 29597 22155 29600
rect 22097 29591 22155 29597
rect 23198 29588 23204 29600
rect 23256 29588 23262 29640
rect 31202 29588 31208 29640
rect 31260 29628 31266 29640
rect 31297 29631 31355 29637
rect 31297 29628 31309 29631
rect 31260 29600 31309 29628
rect 31260 29588 31266 29600
rect 31297 29597 31309 29600
rect 31343 29597 31355 29631
rect 31297 29591 31355 29597
rect 35434 29588 35440 29640
rect 35492 29628 35498 29640
rect 35989 29631 36047 29637
rect 35989 29628 36001 29631
rect 35492 29600 36001 29628
rect 35492 29588 35498 29600
rect 35989 29597 36001 29600
rect 36035 29597 36047 29631
rect 35989 29591 36047 29597
rect 36078 29588 36084 29640
rect 36136 29588 36142 29640
rect 36170 29588 36176 29640
rect 36228 29628 36234 29640
rect 36265 29631 36323 29637
rect 36265 29628 36277 29631
rect 36228 29600 36277 29628
rect 36228 29588 36234 29600
rect 36265 29597 36277 29600
rect 36311 29628 36323 29631
rect 36817 29631 36875 29637
rect 36817 29628 36829 29631
rect 36311 29600 36829 29628
rect 36311 29597 36323 29600
rect 36265 29591 36323 29597
rect 36817 29597 36829 29600
rect 36863 29597 36875 29631
rect 36817 29591 36875 29597
rect 16942 29520 16948 29572
rect 17000 29560 17006 29572
rect 17862 29560 17868 29572
rect 17000 29532 17868 29560
rect 17000 29520 17006 29532
rect 17862 29520 17868 29532
rect 17920 29520 17926 29572
rect 21913 29563 21971 29569
rect 21913 29529 21925 29563
rect 21959 29560 21971 29563
rect 25590 29560 25596 29572
rect 21959 29532 22094 29560
rect 21959 29529 21971 29532
rect 21913 29523 21971 29529
rect 8662 29452 8668 29504
rect 8720 29492 8726 29504
rect 8938 29492 8944 29504
rect 8720 29464 8944 29492
rect 8720 29452 8726 29464
rect 8938 29452 8944 29464
rect 8996 29452 9002 29504
rect 15838 29452 15844 29504
rect 15896 29492 15902 29504
rect 20441 29495 20499 29501
rect 20441 29492 20453 29495
rect 15896 29464 20453 29492
rect 15896 29452 15902 29464
rect 20441 29461 20453 29464
rect 20487 29461 20499 29495
rect 22066 29492 22094 29532
rect 22204 29532 25596 29560
rect 22204 29492 22232 29532
rect 25590 29520 25596 29532
rect 25648 29560 25654 29572
rect 27430 29560 27436 29572
rect 25648 29532 27436 29560
rect 25648 29520 25654 29532
rect 27430 29520 27436 29532
rect 27488 29520 27494 29572
rect 31849 29563 31907 29569
rect 31849 29529 31861 29563
rect 31895 29560 31907 29563
rect 32490 29560 32496 29572
rect 31895 29532 32496 29560
rect 31895 29529 31907 29532
rect 31849 29523 31907 29529
rect 32490 29520 32496 29532
rect 32548 29520 32554 29572
rect 22066 29464 22232 29492
rect 22281 29495 22339 29501
rect 20441 29455 20499 29461
rect 22281 29461 22293 29495
rect 22327 29492 22339 29495
rect 23290 29492 23296 29504
rect 22327 29464 23296 29492
rect 22327 29461 22339 29464
rect 22281 29455 22339 29461
rect 23290 29452 23296 29464
rect 23348 29452 23354 29504
rect 31938 29452 31944 29504
rect 31996 29492 32002 29504
rect 32125 29495 32183 29501
rect 32125 29492 32137 29495
rect 31996 29464 32137 29492
rect 31996 29452 32002 29464
rect 32125 29461 32137 29464
rect 32171 29461 32183 29495
rect 32125 29455 32183 29461
rect 1104 29402 40848 29424
rect 1104 29350 2610 29402
rect 2662 29350 2674 29402
rect 2726 29350 2738 29402
rect 2790 29350 2802 29402
rect 2854 29350 2866 29402
rect 2918 29350 7610 29402
rect 7662 29350 7674 29402
rect 7726 29350 7738 29402
rect 7790 29350 7802 29402
rect 7854 29350 7866 29402
rect 7918 29350 12610 29402
rect 12662 29350 12674 29402
rect 12726 29350 12738 29402
rect 12790 29350 12802 29402
rect 12854 29350 12866 29402
rect 12918 29350 17610 29402
rect 17662 29350 17674 29402
rect 17726 29350 17738 29402
rect 17790 29350 17802 29402
rect 17854 29350 17866 29402
rect 17918 29350 22610 29402
rect 22662 29350 22674 29402
rect 22726 29350 22738 29402
rect 22790 29350 22802 29402
rect 22854 29350 22866 29402
rect 22918 29350 27610 29402
rect 27662 29350 27674 29402
rect 27726 29350 27738 29402
rect 27790 29350 27802 29402
rect 27854 29350 27866 29402
rect 27918 29350 32610 29402
rect 32662 29350 32674 29402
rect 32726 29350 32738 29402
rect 32790 29350 32802 29402
rect 32854 29350 32866 29402
rect 32918 29350 37610 29402
rect 37662 29350 37674 29402
rect 37726 29350 37738 29402
rect 37790 29350 37802 29402
rect 37854 29350 37866 29402
rect 37918 29350 40848 29402
rect 1104 29328 40848 29350
rect 12250 29288 12256 29300
rect 9048 29260 12256 29288
rect 8846 29112 8852 29164
rect 8904 29152 8910 29164
rect 9048 29161 9076 29260
rect 12250 29248 12256 29260
rect 12308 29248 12314 29300
rect 23566 29248 23572 29300
rect 23624 29288 23630 29300
rect 24486 29288 24492 29300
rect 23624 29260 24492 29288
rect 23624 29248 23630 29260
rect 24486 29248 24492 29260
rect 24544 29288 24550 29300
rect 36170 29288 36176 29300
rect 24544 29260 36176 29288
rect 24544 29248 24550 29260
rect 36170 29248 36176 29260
rect 36228 29248 36234 29300
rect 38930 29248 38936 29300
rect 38988 29248 38994 29300
rect 12526 29180 12532 29232
rect 12584 29220 12590 29232
rect 31662 29220 31668 29232
rect 12584 29192 31668 29220
rect 12584 29180 12590 29192
rect 31662 29180 31668 29192
rect 31720 29180 31726 29232
rect 9033 29155 9091 29161
rect 9033 29152 9045 29155
rect 8904 29124 9045 29152
rect 8904 29112 8910 29124
rect 9033 29121 9045 29124
rect 9079 29121 9091 29155
rect 9033 29115 9091 29121
rect 9401 29155 9459 29161
rect 9401 29121 9413 29155
rect 9447 29121 9459 29155
rect 9401 29115 9459 29121
rect 9677 29155 9735 29161
rect 9677 29121 9689 29155
rect 9723 29152 9735 29155
rect 11974 29152 11980 29164
rect 9723 29124 11980 29152
rect 9723 29121 9735 29124
rect 9677 29115 9735 29121
rect 4706 29044 4712 29096
rect 4764 29084 4770 29096
rect 6822 29084 6828 29096
rect 4764 29056 6828 29084
rect 4764 29044 4770 29056
rect 6822 29044 6828 29056
rect 6880 29044 6886 29096
rect 9416 29016 9444 29115
rect 11974 29112 11980 29124
rect 12032 29112 12038 29164
rect 12250 29112 12256 29164
rect 12308 29152 12314 29164
rect 12345 29155 12403 29161
rect 12345 29152 12357 29155
rect 12308 29124 12357 29152
rect 12308 29112 12314 29124
rect 12345 29121 12357 29124
rect 12391 29152 12403 29155
rect 17402 29152 17408 29164
rect 12391 29124 17408 29152
rect 12391 29121 12403 29124
rect 12345 29115 12403 29121
rect 17402 29112 17408 29124
rect 17460 29112 17466 29164
rect 30926 29112 30932 29164
rect 30984 29152 30990 29164
rect 38473 29155 38531 29161
rect 38473 29152 38485 29155
rect 30984 29124 38485 29152
rect 30984 29112 30990 29124
rect 38473 29121 38485 29124
rect 38519 29121 38531 29155
rect 38473 29115 38531 29121
rect 38749 29155 38807 29161
rect 38749 29121 38761 29155
rect 38795 29121 38807 29155
rect 38749 29115 38807 29121
rect 10594 29044 10600 29096
rect 10652 29084 10658 29096
rect 10689 29087 10747 29093
rect 10689 29084 10701 29087
rect 10652 29056 10701 29084
rect 10652 29044 10658 29056
rect 10689 29053 10701 29056
rect 10735 29053 10747 29087
rect 10689 29047 10747 29053
rect 11330 29044 11336 29096
rect 11388 29044 11394 29096
rect 12437 29087 12495 29093
rect 12437 29084 12449 29087
rect 11440 29056 12449 29084
rect 11440 29016 11468 29056
rect 12437 29053 12449 29056
rect 12483 29084 12495 29087
rect 16298 29084 16304 29096
rect 12483 29056 16304 29084
rect 12483 29053 12495 29056
rect 12437 29047 12495 29053
rect 16298 29044 16304 29056
rect 16356 29084 16362 29096
rect 16942 29084 16948 29096
rect 16356 29056 16948 29084
rect 16356 29044 16362 29056
rect 16942 29044 16948 29056
rect 17000 29044 17006 29096
rect 30098 29044 30104 29096
rect 30156 29084 30162 29096
rect 38565 29087 38623 29093
rect 38565 29084 38577 29087
rect 30156 29056 38577 29084
rect 30156 29044 30162 29056
rect 38565 29053 38577 29056
rect 38611 29053 38623 29087
rect 38565 29047 38623 29053
rect 9416 28988 11468 29016
rect 11514 28976 11520 29028
rect 11572 29016 11578 29028
rect 11790 29016 11796 29028
rect 11572 28988 11796 29016
rect 11572 28976 11578 28988
rect 11790 28976 11796 28988
rect 11848 28976 11854 29028
rect 11974 28976 11980 29028
rect 12032 29016 12038 29028
rect 12526 29016 12532 29028
rect 12032 28988 12532 29016
rect 12032 28976 12038 28988
rect 12526 28976 12532 28988
rect 12584 28976 12590 29028
rect 16666 28976 16672 29028
rect 16724 29016 16730 29028
rect 17862 29016 17868 29028
rect 16724 28988 17868 29016
rect 16724 28976 16730 28988
rect 17862 28976 17868 28988
rect 17920 28976 17926 29028
rect 33226 28976 33232 29028
rect 33284 29016 33290 29028
rect 33962 29016 33968 29028
rect 33284 28988 33968 29016
rect 33284 28976 33290 28988
rect 33962 28976 33968 28988
rect 34020 29016 34026 29028
rect 38764 29016 38792 29115
rect 34020 28988 38792 29016
rect 34020 28976 34026 28988
rect 9122 28908 9128 28960
rect 9180 28908 9186 28960
rect 9674 28908 9680 28960
rect 9732 28948 9738 28960
rect 10042 28948 10048 28960
rect 9732 28920 10048 28948
rect 9732 28908 9738 28920
rect 10042 28908 10048 28920
rect 10100 28948 10106 28960
rect 17770 28948 17776 28960
rect 10100 28920 17776 28948
rect 10100 28908 10106 28920
rect 17770 28908 17776 28920
rect 17828 28908 17834 28960
rect 25314 28908 25320 28960
rect 25372 28948 25378 28960
rect 25958 28948 25964 28960
rect 25372 28920 25964 28948
rect 25372 28908 25378 28920
rect 25958 28908 25964 28920
rect 26016 28908 26022 28960
rect 1104 28858 40848 28880
rect 1104 28806 1950 28858
rect 2002 28806 2014 28858
rect 2066 28806 2078 28858
rect 2130 28806 2142 28858
rect 2194 28806 2206 28858
rect 2258 28806 6950 28858
rect 7002 28806 7014 28858
rect 7066 28806 7078 28858
rect 7130 28806 7142 28858
rect 7194 28806 7206 28858
rect 7258 28806 11950 28858
rect 12002 28806 12014 28858
rect 12066 28806 12078 28858
rect 12130 28806 12142 28858
rect 12194 28806 12206 28858
rect 12258 28806 16950 28858
rect 17002 28806 17014 28858
rect 17066 28806 17078 28858
rect 17130 28806 17142 28858
rect 17194 28806 17206 28858
rect 17258 28806 21950 28858
rect 22002 28806 22014 28858
rect 22066 28806 22078 28858
rect 22130 28806 22142 28858
rect 22194 28806 22206 28858
rect 22258 28806 26950 28858
rect 27002 28806 27014 28858
rect 27066 28806 27078 28858
rect 27130 28806 27142 28858
rect 27194 28806 27206 28858
rect 27258 28806 31950 28858
rect 32002 28806 32014 28858
rect 32066 28806 32078 28858
rect 32130 28806 32142 28858
rect 32194 28806 32206 28858
rect 32258 28806 36950 28858
rect 37002 28806 37014 28858
rect 37066 28806 37078 28858
rect 37130 28806 37142 28858
rect 37194 28806 37206 28858
rect 37258 28806 40848 28858
rect 1104 28784 40848 28806
rect 10873 28747 10931 28753
rect 10873 28713 10885 28747
rect 10919 28744 10931 28747
rect 16850 28744 16856 28756
rect 10919 28716 16856 28744
rect 10919 28713 10931 28716
rect 10873 28707 10931 28713
rect 16850 28704 16856 28716
rect 16908 28704 16914 28756
rect 16942 28704 16948 28756
rect 17000 28744 17006 28756
rect 18690 28744 18696 28756
rect 17000 28716 18696 28744
rect 17000 28704 17006 28716
rect 18690 28704 18696 28716
rect 18748 28704 18754 28756
rect 23934 28744 23940 28756
rect 22066 28716 23940 28744
rect 22066 28676 22094 28716
rect 23934 28704 23940 28716
rect 23992 28704 23998 28756
rect 12406 28648 22094 28676
rect 10778 28500 10784 28552
rect 10836 28500 10842 28552
rect 10965 28543 11023 28549
rect 10965 28509 10977 28543
rect 11011 28540 11023 28543
rect 12406 28540 12434 28648
rect 17402 28568 17408 28620
rect 17460 28568 17466 28620
rect 17770 28568 17776 28620
rect 17828 28568 17834 28620
rect 24394 28568 24400 28620
rect 24452 28608 24458 28620
rect 24489 28611 24547 28617
rect 24489 28608 24501 28611
rect 24452 28580 24501 28608
rect 24452 28568 24458 28580
rect 24489 28577 24501 28580
rect 24535 28577 24547 28611
rect 24489 28571 24547 28577
rect 11011 28512 12434 28540
rect 11011 28509 11023 28512
rect 10965 28503 11023 28509
rect 15930 28500 15936 28552
rect 15988 28540 15994 28552
rect 16301 28543 16359 28549
rect 16301 28540 16313 28543
rect 15988 28512 16313 28540
rect 15988 28500 15994 28512
rect 16301 28509 16313 28512
rect 16347 28509 16359 28543
rect 16301 28503 16359 28509
rect 16393 28543 16451 28549
rect 16393 28509 16405 28543
rect 16439 28509 16451 28543
rect 16393 28503 16451 28509
rect 16577 28543 16635 28549
rect 16577 28509 16589 28543
rect 16623 28540 16635 28543
rect 16942 28540 16948 28552
rect 16623 28512 16948 28540
rect 16623 28509 16635 28512
rect 16577 28503 16635 28509
rect 10686 28432 10692 28484
rect 10744 28472 10750 28484
rect 16408 28472 16436 28503
rect 16942 28500 16948 28512
rect 17000 28500 17006 28552
rect 17313 28543 17371 28549
rect 17313 28509 17325 28543
rect 17359 28509 17371 28543
rect 17313 28503 17371 28509
rect 10744 28444 16436 28472
rect 10744 28432 10750 28444
rect 16666 28432 16672 28484
rect 16724 28472 16730 28484
rect 17129 28475 17187 28481
rect 17129 28472 17141 28475
rect 16724 28444 17141 28472
rect 16724 28432 16730 28444
rect 17129 28441 17141 28444
rect 17175 28441 17187 28475
rect 17328 28472 17356 28503
rect 20714 28500 20720 28552
rect 20772 28540 20778 28552
rect 24765 28543 24823 28549
rect 24765 28540 24777 28543
rect 20772 28512 24777 28540
rect 20772 28500 20778 28512
rect 24765 28509 24777 28512
rect 24811 28509 24823 28543
rect 24765 28503 24823 28509
rect 25314 28472 25320 28484
rect 17328 28444 25320 28472
rect 17129 28435 17187 28441
rect 25314 28432 25320 28444
rect 25372 28432 25378 28484
rect 16761 28407 16819 28413
rect 16761 28373 16773 28407
rect 16807 28404 16819 28407
rect 19794 28404 19800 28416
rect 16807 28376 19800 28404
rect 16807 28373 16819 28376
rect 16761 28367 16819 28373
rect 19794 28364 19800 28376
rect 19852 28364 19858 28416
rect 1104 28314 40848 28336
rect 1104 28262 2610 28314
rect 2662 28262 2674 28314
rect 2726 28262 2738 28314
rect 2790 28262 2802 28314
rect 2854 28262 2866 28314
rect 2918 28262 7610 28314
rect 7662 28262 7674 28314
rect 7726 28262 7738 28314
rect 7790 28262 7802 28314
rect 7854 28262 7866 28314
rect 7918 28262 12610 28314
rect 12662 28262 12674 28314
rect 12726 28262 12738 28314
rect 12790 28262 12802 28314
rect 12854 28262 12866 28314
rect 12918 28262 17610 28314
rect 17662 28262 17674 28314
rect 17726 28262 17738 28314
rect 17790 28262 17802 28314
rect 17854 28262 17866 28314
rect 17918 28262 22610 28314
rect 22662 28262 22674 28314
rect 22726 28262 22738 28314
rect 22790 28262 22802 28314
rect 22854 28262 22866 28314
rect 22918 28262 27610 28314
rect 27662 28262 27674 28314
rect 27726 28262 27738 28314
rect 27790 28262 27802 28314
rect 27854 28262 27866 28314
rect 27918 28262 32610 28314
rect 32662 28262 32674 28314
rect 32726 28262 32738 28314
rect 32790 28262 32802 28314
rect 32854 28262 32866 28314
rect 32918 28262 37610 28314
rect 37662 28262 37674 28314
rect 37726 28262 37738 28314
rect 37790 28262 37802 28314
rect 37854 28262 37866 28314
rect 37918 28262 40848 28314
rect 1104 28240 40848 28262
rect 16942 28160 16948 28212
rect 17000 28200 17006 28212
rect 17402 28200 17408 28212
rect 17000 28172 17408 28200
rect 17000 28160 17006 28172
rect 17402 28160 17408 28172
rect 17460 28160 17466 28212
rect 24854 28160 24860 28212
rect 24912 28160 24918 28212
rect 5534 28092 5540 28144
rect 5592 28132 5598 28144
rect 5592 28104 31432 28132
rect 5592 28092 5598 28104
rect 24394 28024 24400 28076
rect 24452 28024 24458 28076
rect 24670 28024 24676 28076
rect 24728 28024 24734 28076
rect 30926 28024 30932 28076
rect 30984 28064 30990 28076
rect 31404 28073 31432 28104
rect 31021 28067 31079 28073
rect 31021 28064 31033 28067
rect 30984 28036 31033 28064
rect 30984 28024 30990 28036
rect 31021 28033 31033 28036
rect 31067 28033 31079 28067
rect 31021 28027 31079 28033
rect 31389 28067 31447 28073
rect 31389 28033 31401 28067
rect 31435 28033 31447 28067
rect 31389 28027 31447 28033
rect 11698 27956 11704 28008
rect 11756 27996 11762 28008
rect 31757 27999 31815 28005
rect 31757 27996 31769 27999
rect 11756 27968 31769 27996
rect 11756 27956 11762 27968
rect 31757 27965 31769 27968
rect 31803 27965 31815 27999
rect 31757 27959 31815 27965
rect 22370 27888 22376 27940
rect 22428 27928 22434 27940
rect 24489 27931 24547 27937
rect 24489 27928 24501 27931
rect 22428 27900 24501 27928
rect 22428 27888 22434 27900
rect 24489 27897 24501 27900
rect 24535 27897 24547 27931
rect 31021 27931 31079 27937
rect 31021 27928 31033 27931
rect 24489 27891 24547 27897
rect 26206 27900 31033 27928
rect 20806 27820 20812 27872
rect 20864 27860 20870 27872
rect 21542 27860 21548 27872
rect 20864 27832 21548 27860
rect 20864 27820 20870 27832
rect 21542 27820 21548 27832
rect 21600 27860 21606 27872
rect 26206 27860 26234 27900
rect 31021 27897 31033 27900
rect 31067 27897 31079 27931
rect 31021 27891 31079 27897
rect 21600 27832 26234 27860
rect 21600 27820 21606 27832
rect 32950 27820 32956 27872
rect 33008 27860 33014 27872
rect 35986 27860 35992 27872
rect 33008 27832 35992 27860
rect 33008 27820 33014 27832
rect 35986 27820 35992 27832
rect 36044 27820 36050 27872
rect 1104 27770 40848 27792
rect 1104 27718 1950 27770
rect 2002 27718 2014 27770
rect 2066 27718 2078 27770
rect 2130 27718 2142 27770
rect 2194 27718 2206 27770
rect 2258 27718 6950 27770
rect 7002 27718 7014 27770
rect 7066 27718 7078 27770
rect 7130 27718 7142 27770
rect 7194 27718 7206 27770
rect 7258 27718 11950 27770
rect 12002 27718 12014 27770
rect 12066 27718 12078 27770
rect 12130 27718 12142 27770
rect 12194 27718 12206 27770
rect 12258 27718 16950 27770
rect 17002 27718 17014 27770
rect 17066 27718 17078 27770
rect 17130 27718 17142 27770
rect 17194 27718 17206 27770
rect 17258 27718 21950 27770
rect 22002 27718 22014 27770
rect 22066 27718 22078 27770
rect 22130 27718 22142 27770
rect 22194 27718 22206 27770
rect 22258 27718 26950 27770
rect 27002 27718 27014 27770
rect 27066 27718 27078 27770
rect 27130 27718 27142 27770
rect 27194 27718 27206 27770
rect 27258 27718 31950 27770
rect 32002 27718 32014 27770
rect 32066 27718 32078 27770
rect 32130 27718 32142 27770
rect 32194 27718 32206 27770
rect 32258 27718 36950 27770
rect 37002 27718 37014 27770
rect 37066 27718 37078 27770
rect 37130 27718 37142 27770
rect 37194 27718 37206 27770
rect 37258 27718 40848 27770
rect 1104 27696 40848 27718
rect 17218 27616 17224 27668
rect 17276 27656 17282 27668
rect 17402 27656 17408 27668
rect 17276 27628 17408 27656
rect 17276 27616 17282 27628
rect 17402 27616 17408 27628
rect 17460 27616 17466 27668
rect 19794 27616 19800 27668
rect 19852 27656 19858 27668
rect 20622 27656 20628 27668
rect 19852 27628 20628 27656
rect 19852 27616 19858 27628
rect 20622 27616 20628 27628
rect 20680 27616 20686 27668
rect 34514 27616 34520 27668
rect 34572 27656 34578 27668
rect 34793 27659 34851 27665
rect 34793 27656 34805 27659
rect 34572 27628 34805 27656
rect 34572 27616 34578 27628
rect 34793 27625 34805 27628
rect 34839 27625 34851 27659
rect 34793 27619 34851 27625
rect 23290 27548 23296 27600
rect 23348 27588 23354 27600
rect 24210 27588 24216 27600
rect 23348 27560 24216 27588
rect 23348 27548 23354 27560
rect 24210 27548 24216 27560
rect 24268 27548 24274 27600
rect 33410 27480 33416 27532
rect 33468 27520 33474 27532
rect 33468 27492 35480 27520
rect 33468 27480 33474 27492
rect 32490 27412 32496 27464
rect 32548 27452 32554 27464
rect 35452 27461 35480 27492
rect 34701 27455 34759 27461
rect 34701 27452 34713 27455
rect 32548 27424 34713 27452
rect 32548 27412 32554 27424
rect 34701 27421 34713 27424
rect 34747 27421 34759 27455
rect 34701 27415 34759 27421
rect 35069 27455 35127 27461
rect 35069 27421 35081 27455
rect 35115 27421 35127 27455
rect 35069 27415 35127 27421
rect 35437 27455 35495 27461
rect 35437 27421 35449 27455
rect 35483 27421 35495 27455
rect 35437 27415 35495 27421
rect 30374 27344 30380 27396
rect 30432 27384 30438 27396
rect 35084 27384 35112 27415
rect 30432 27356 35112 27384
rect 30432 27344 30438 27356
rect 1104 27226 40848 27248
rect 1104 27174 2610 27226
rect 2662 27174 2674 27226
rect 2726 27174 2738 27226
rect 2790 27174 2802 27226
rect 2854 27174 2866 27226
rect 2918 27174 7610 27226
rect 7662 27174 7674 27226
rect 7726 27174 7738 27226
rect 7790 27174 7802 27226
rect 7854 27174 7866 27226
rect 7918 27174 12610 27226
rect 12662 27174 12674 27226
rect 12726 27174 12738 27226
rect 12790 27174 12802 27226
rect 12854 27174 12866 27226
rect 12918 27174 17610 27226
rect 17662 27174 17674 27226
rect 17726 27174 17738 27226
rect 17790 27174 17802 27226
rect 17854 27174 17866 27226
rect 17918 27174 22610 27226
rect 22662 27174 22674 27226
rect 22726 27174 22738 27226
rect 22790 27174 22802 27226
rect 22854 27174 22866 27226
rect 22918 27174 27610 27226
rect 27662 27174 27674 27226
rect 27726 27174 27738 27226
rect 27790 27174 27802 27226
rect 27854 27174 27866 27226
rect 27918 27174 32610 27226
rect 32662 27174 32674 27226
rect 32726 27174 32738 27226
rect 32790 27174 32802 27226
rect 32854 27174 32866 27226
rect 32918 27174 37610 27226
rect 37662 27174 37674 27226
rect 37726 27174 37738 27226
rect 37790 27174 37802 27226
rect 37854 27174 37866 27226
rect 37918 27174 40848 27226
rect 1104 27152 40848 27174
rect 16574 27004 16580 27056
rect 16632 27044 16638 27056
rect 17402 27044 17408 27056
rect 16632 27016 17408 27044
rect 16632 27004 16638 27016
rect 17402 27004 17408 27016
rect 17460 27004 17466 27056
rect 13906 26936 13912 26988
rect 13964 26976 13970 26988
rect 17957 26979 18015 26985
rect 17957 26976 17969 26979
rect 13964 26948 17969 26976
rect 13964 26936 13970 26948
rect 17957 26945 17969 26948
rect 18003 26945 18015 26979
rect 17957 26939 18015 26945
rect 18417 26979 18475 26985
rect 18417 26945 18429 26979
rect 18463 26945 18475 26979
rect 18417 26939 18475 26945
rect 18509 26979 18567 26985
rect 18509 26945 18521 26979
rect 18555 26976 18567 26979
rect 18555 26948 22094 26976
rect 18555 26945 18567 26948
rect 18509 26939 18567 26945
rect 4062 26800 4068 26852
rect 4120 26840 4126 26852
rect 17586 26840 17592 26852
rect 4120 26812 17592 26840
rect 4120 26800 4126 26812
rect 17586 26800 17592 26812
rect 17644 26800 17650 26852
rect 18432 26840 18460 26939
rect 18598 26868 18604 26920
rect 18656 26908 18662 26920
rect 18693 26911 18751 26917
rect 18693 26908 18705 26911
rect 18656 26880 18705 26908
rect 18656 26868 18662 26880
rect 18693 26877 18705 26880
rect 18739 26908 18751 26911
rect 19150 26908 19156 26920
rect 18739 26880 19156 26908
rect 18739 26877 18751 26880
rect 18693 26871 18751 26877
rect 19150 26868 19156 26880
rect 19208 26868 19214 26920
rect 22066 26908 22094 26948
rect 23106 26908 23112 26920
rect 22066 26880 23112 26908
rect 23106 26868 23112 26880
rect 23164 26908 23170 26920
rect 33410 26908 33416 26920
rect 23164 26880 33416 26908
rect 23164 26868 23170 26880
rect 33410 26868 33416 26880
rect 33468 26908 33474 26920
rect 38562 26908 38568 26920
rect 33468 26880 38568 26908
rect 33468 26868 33474 26880
rect 38562 26868 38568 26880
rect 38620 26868 38626 26920
rect 26510 26840 26516 26852
rect 18432 26812 26516 26840
rect 26510 26800 26516 26812
rect 26568 26800 26574 26852
rect 1104 26682 40848 26704
rect 1104 26630 1950 26682
rect 2002 26630 2014 26682
rect 2066 26630 2078 26682
rect 2130 26630 2142 26682
rect 2194 26630 2206 26682
rect 2258 26630 6950 26682
rect 7002 26630 7014 26682
rect 7066 26630 7078 26682
rect 7130 26630 7142 26682
rect 7194 26630 7206 26682
rect 7258 26630 11950 26682
rect 12002 26630 12014 26682
rect 12066 26630 12078 26682
rect 12130 26630 12142 26682
rect 12194 26630 12206 26682
rect 12258 26630 16950 26682
rect 17002 26630 17014 26682
rect 17066 26630 17078 26682
rect 17130 26630 17142 26682
rect 17194 26630 17206 26682
rect 17258 26630 21950 26682
rect 22002 26630 22014 26682
rect 22066 26630 22078 26682
rect 22130 26630 22142 26682
rect 22194 26630 22206 26682
rect 22258 26630 26950 26682
rect 27002 26630 27014 26682
rect 27066 26630 27078 26682
rect 27130 26630 27142 26682
rect 27194 26630 27206 26682
rect 27258 26630 31950 26682
rect 32002 26630 32014 26682
rect 32066 26630 32078 26682
rect 32130 26630 32142 26682
rect 32194 26630 32206 26682
rect 32258 26630 36950 26682
rect 37002 26630 37014 26682
rect 37066 26630 37078 26682
rect 37130 26630 37142 26682
rect 37194 26630 37206 26682
rect 37258 26630 40848 26682
rect 1104 26608 40848 26630
rect 32585 26571 32643 26577
rect 32585 26537 32597 26571
rect 32631 26568 32643 26571
rect 36630 26568 36636 26580
rect 32631 26540 36636 26568
rect 32631 26537 32643 26540
rect 32585 26531 32643 26537
rect 24946 26460 24952 26512
rect 25004 26500 25010 26512
rect 31205 26503 31263 26509
rect 31205 26500 31217 26503
rect 25004 26472 31217 26500
rect 25004 26460 25010 26472
rect 31205 26469 31217 26472
rect 31251 26500 31263 26503
rect 31251 26472 32168 26500
rect 31251 26469 31263 26472
rect 31205 26463 31263 26469
rect 9582 26432 9588 26444
rect 4080 26404 9588 26432
rect 4080 26373 4108 26404
rect 9582 26392 9588 26404
rect 9640 26392 9646 26444
rect 16390 26392 16396 26444
rect 16448 26432 16454 26444
rect 19242 26432 19248 26444
rect 16448 26404 19248 26432
rect 16448 26392 16454 26404
rect 19242 26392 19248 26404
rect 19300 26432 19306 26444
rect 32140 26441 32168 26472
rect 32125 26435 32183 26441
rect 19300 26404 30972 26432
rect 19300 26392 19306 26404
rect 4065 26367 4123 26373
rect 4065 26333 4077 26367
rect 4111 26333 4123 26367
rect 4065 26327 4123 26333
rect 4249 26367 4307 26373
rect 4249 26333 4261 26367
rect 4295 26333 4307 26367
rect 4249 26327 4307 26333
rect 4617 26367 4675 26373
rect 4617 26333 4629 26367
rect 4663 26364 4675 26367
rect 4706 26364 4712 26376
rect 4663 26336 4712 26364
rect 4663 26333 4675 26336
rect 4617 26327 4675 26333
rect 4264 26296 4292 26327
rect 4706 26324 4712 26336
rect 4764 26324 4770 26376
rect 17218 26324 17224 26376
rect 17276 26364 17282 26376
rect 17586 26364 17592 26376
rect 17276 26336 17592 26364
rect 17276 26324 17282 26336
rect 17586 26324 17592 26336
rect 17644 26364 17650 26376
rect 30944 26364 30972 26404
rect 32125 26401 32137 26435
rect 32171 26401 32183 26435
rect 32125 26395 32183 26401
rect 32217 26435 32275 26441
rect 32217 26401 32229 26435
rect 32263 26432 32275 26435
rect 32600 26432 32628 26531
rect 36630 26528 36636 26540
rect 36688 26528 36694 26580
rect 32263 26404 32628 26432
rect 32263 26401 32275 26404
rect 32217 26395 32275 26401
rect 31573 26367 31631 26373
rect 31573 26364 31585 26367
rect 17644 26336 30880 26364
rect 30944 26336 31585 26364
rect 17644 26324 17650 26336
rect 9674 26296 9680 26308
rect 4264 26268 9680 26296
rect 9674 26256 9680 26268
rect 9732 26256 9738 26308
rect 15194 26256 15200 26308
rect 15252 26296 15258 26308
rect 30852 26296 30880 26336
rect 31573 26333 31585 26336
rect 31619 26333 31631 26367
rect 31573 26327 31631 26333
rect 31754 26324 31760 26376
rect 31812 26364 31818 26376
rect 31812 26336 31857 26364
rect 31812 26324 31818 26336
rect 32232 26296 32260 26395
rect 15252 26268 28994 26296
rect 30852 26268 32260 26296
rect 15252 26256 15258 26268
rect 6270 26188 6276 26240
rect 6328 26228 6334 26240
rect 6454 26228 6460 26240
rect 6328 26200 6460 26228
rect 6328 26188 6334 26200
rect 6454 26188 6460 26200
rect 6512 26188 6518 26240
rect 28966 26228 28994 26268
rect 30837 26231 30895 26237
rect 30837 26228 30849 26231
rect 28966 26200 30849 26228
rect 30837 26197 30849 26200
rect 30883 26228 30895 26231
rect 31754 26228 31760 26240
rect 30883 26200 31760 26228
rect 30883 26197 30895 26200
rect 30837 26191 30895 26197
rect 31754 26188 31760 26200
rect 31812 26188 31818 26240
rect 37366 26188 37372 26240
rect 37424 26228 37430 26240
rect 37550 26228 37556 26240
rect 37424 26200 37556 26228
rect 37424 26188 37430 26200
rect 37550 26188 37556 26200
rect 37608 26188 37614 26240
rect 1104 26138 40848 26160
rect 1104 26086 2610 26138
rect 2662 26086 2674 26138
rect 2726 26086 2738 26138
rect 2790 26086 2802 26138
rect 2854 26086 2866 26138
rect 2918 26086 7610 26138
rect 7662 26086 7674 26138
rect 7726 26086 7738 26138
rect 7790 26086 7802 26138
rect 7854 26086 7866 26138
rect 7918 26086 12610 26138
rect 12662 26086 12674 26138
rect 12726 26086 12738 26138
rect 12790 26086 12802 26138
rect 12854 26086 12866 26138
rect 12918 26086 17610 26138
rect 17662 26086 17674 26138
rect 17726 26086 17738 26138
rect 17790 26086 17802 26138
rect 17854 26086 17866 26138
rect 17918 26086 22610 26138
rect 22662 26086 22674 26138
rect 22726 26086 22738 26138
rect 22790 26086 22802 26138
rect 22854 26086 22866 26138
rect 22918 26086 27610 26138
rect 27662 26086 27674 26138
rect 27726 26086 27738 26138
rect 27790 26086 27802 26138
rect 27854 26086 27866 26138
rect 27918 26086 32610 26138
rect 32662 26086 32674 26138
rect 32726 26086 32738 26138
rect 32790 26086 32802 26138
rect 32854 26086 32866 26138
rect 32918 26086 37610 26138
rect 37662 26086 37674 26138
rect 37726 26086 37738 26138
rect 37790 26086 37802 26138
rect 37854 26086 37866 26138
rect 37918 26086 40848 26138
rect 1104 26064 40848 26086
rect 6454 25984 6460 26036
rect 6512 26024 6518 26036
rect 6512 25996 12434 26024
rect 6512 25984 6518 25996
rect 1670 25916 1676 25968
rect 1728 25956 1734 25968
rect 2406 25956 2412 25968
rect 1728 25928 2412 25956
rect 1728 25916 1734 25928
rect 2406 25916 2412 25928
rect 2464 25956 2470 25968
rect 2464 25928 7420 25956
rect 2464 25916 2470 25928
rect 5902 25848 5908 25900
rect 5960 25888 5966 25900
rect 6638 25888 6644 25900
rect 5960 25860 6644 25888
rect 5960 25848 5966 25860
rect 6638 25848 6644 25860
rect 6696 25848 6702 25900
rect 7392 25897 7420 25928
rect 7466 25916 7472 25968
rect 7524 25956 7530 25968
rect 8386 25956 8392 25968
rect 7524 25928 8392 25956
rect 7524 25916 7530 25928
rect 7668 25897 7696 25928
rect 8386 25916 8392 25928
rect 8444 25916 8450 25968
rect 7377 25891 7435 25897
rect 7377 25857 7389 25891
rect 7423 25857 7435 25891
rect 7377 25851 7435 25857
rect 7653 25891 7711 25897
rect 7653 25857 7665 25891
rect 7699 25857 7711 25891
rect 7653 25851 7711 25857
rect 8113 25891 8171 25897
rect 8113 25857 8125 25891
rect 8159 25888 8171 25891
rect 9030 25888 9036 25900
rect 8159 25860 9036 25888
rect 8159 25857 8171 25860
rect 8113 25851 8171 25857
rect 5534 25780 5540 25832
rect 5592 25820 5598 25832
rect 6917 25823 6975 25829
rect 6917 25820 6929 25823
rect 5592 25792 6929 25820
rect 5592 25780 5598 25792
rect 6917 25789 6929 25792
rect 6963 25789 6975 25823
rect 7392 25820 7420 25851
rect 9030 25848 9036 25860
rect 9088 25848 9094 25900
rect 12406 25888 12434 25996
rect 17494 25984 17500 26036
rect 17552 26024 17558 26036
rect 17589 26027 17647 26033
rect 17589 26024 17601 26027
rect 17552 25996 17601 26024
rect 17552 25984 17558 25996
rect 17589 25993 17601 25996
rect 17635 25993 17647 26027
rect 17589 25987 17647 25993
rect 18046 25916 18052 25968
rect 18104 25916 18110 25968
rect 25225 25959 25283 25965
rect 25225 25925 25237 25959
rect 25271 25956 25283 25959
rect 25314 25956 25320 25968
rect 25271 25928 25320 25956
rect 25271 25925 25283 25928
rect 25225 25919 25283 25925
rect 25314 25916 25320 25928
rect 25372 25916 25378 25968
rect 24673 25891 24731 25897
rect 24673 25888 24685 25891
rect 12406 25860 24685 25888
rect 24673 25857 24685 25860
rect 24719 25857 24731 25891
rect 24673 25851 24731 25857
rect 24857 25891 24915 25897
rect 24857 25857 24869 25891
rect 24903 25888 24915 25891
rect 25130 25888 25136 25900
rect 24903 25860 25136 25888
rect 24903 25857 24915 25860
rect 24857 25851 24915 25857
rect 25130 25848 25136 25860
rect 25188 25848 25194 25900
rect 11054 25820 11060 25832
rect 7392 25792 11060 25820
rect 6917 25783 6975 25789
rect 11054 25780 11060 25792
rect 11112 25780 11118 25832
rect 17218 25780 17224 25832
rect 17276 25820 17282 25832
rect 17402 25820 17408 25832
rect 17276 25792 17408 25820
rect 17276 25780 17282 25792
rect 17402 25780 17408 25792
rect 17460 25780 17466 25832
rect 18966 25780 18972 25832
rect 19024 25820 19030 25832
rect 31018 25820 31024 25832
rect 19024 25792 31024 25820
rect 19024 25780 19030 25792
rect 31018 25780 31024 25792
rect 31076 25780 31082 25832
rect 16850 25712 16856 25764
rect 16908 25752 16914 25764
rect 17681 25755 17739 25761
rect 17681 25752 17693 25755
rect 16908 25724 17693 25752
rect 16908 25712 16914 25724
rect 17681 25721 17693 25724
rect 17727 25721 17739 25755
rect 17681 25715 17739 25721
rect 24302 25712 24308 25764
rect 24360 25752 24366 25764
rect 38930 25752 38936 25764
rect 24360 25724 38936 25752
rect 24360 25712 24366 25724
rect 38930 25712 38936 25724
rect 38988 25712 38994 25764
rect 15654 25644 15660 25696
rect 15712 25684 15718 25696
rect 26050 25684 26056 25696
rect 15712 25656 26056 25684
rect 15712 25644 15718 25656
rect 26050 25644 26056 25656
rect 26108 25644 26114 25696
rect 1104 25594 40848 25616
rect 1104 25542 1950 25594
rect 2002 25542 2014 25594
rect 2066 25542 2078 25594
rect 2130 25542 2142 25594
rect 2194 25542 2206 25594
rect 2258 25542 6950 25594
rect 7002 25542 7014 25594
rect 7066 25542 7078 25594
rect 7130 25542 7142 25594
rect 7194 25542 7206 25594
rect 7258 25542 11950 25594
rect 12002 25542 12014 25594
rect 12066 25542 12078 25594
rect 12130 25542 12142 25594
rect 12194 25542 12206 25594
rect 12258 25542 16950 25594
rect 17002 25542 17014 25594
rect 17066 25542 17078 25594
rect 17130 25542 17142 25594
rect 17194 25542 17206 25594
rect 17258 25542 21950 25594
rect 22002 25542 22014 25594
rect 22066 25542 22078 25594
rect 22130 25542 22142 25594
rect 22194 25542 22206 25594
rect 22258 25542 26950 25594
rect 27002 25542 27014 25594
rect 27066 25542 27078 25594
rect 27130 25542 27142 25594
rect 27194 25542 27206 25594
rect 27258 25542 31950 25594
rect 32002 25542 32014 25594
rect 32066 25542 32078 25594
rect 32130 25542 32142 25594
rect 32194 25542 32206 25594
rect 32258 25542 36950 25594
rect 37002 25542 37014 25594
rect 37066 25542 37078 25594
rect 37130 25542 37142 25594
rect 37194 25542 37206 25594
rect 37258 25542 40848 25594
rect 1104 25520 40848 25542
rect 16298 25440 16304 25492
rect 16356 25480 16362 25492
rect 16850 25480 16856 25492
rect 16356 25452 16856 25480
rect 16356 25440 16362 25452
rect 16850 25440 16856 25452
rect 16908 25440 16914 25492
rect 10689 25415 10747 25421
rect 10689 25381 10701 25415
rect 10735 25412 10747 25415
rect 15930 25412 15936 25424
rect 10735 25384 15936 25412
rect 10735 25381 10747 25384
rect 10689 25375 10747 25381
rect 15930 25372 15936 25384
rect 15988 25372 15994 25424
rect 34054 25372 34060 25424
rect 34112 25412 34118 25424
rect 34112 25384 38608 25412
rect 34112 25372 34118 25384
rect 10505 25347 10563 25353
rect 10505 25313 10517 25347
rect 10551 25344 10563 25347
rect 17310 25344 17316 25356
rect 10551 25316 17316 25344
rect 10551 25313 10563 25316
rect 10505 25307 10563 25313
rect 17310 25304 17316 25316
rect 17368 25304 17374 25356
rect 38105 25347 38163 25353
rect 38105 25313 38117 25347
rect 38151 25344 38163 25347
rect 38194 25344 38200 25356
rect 38151 25316 38200 25344
rect 38151 25313 38163 25316
rect 38105 25307 38163 25313
rect 38194 25304 38200 25316
rect 38252 25304 38258 25356
rect 38580 25353 38608 25384
rect 38565 25347 38623 25353
rect 38565 25313 38577 25347
rect 38611 25313 38623 25347
rect 38565 25307 38623 25313
rect 10686 25236 10692 25288
rect 10744 25276 10750 25288
rect 10781 25279 10839 25285
rect 10781 25276 10793 25279
rect 10744 25248 10793 25276
rect 10744 25236 10750 25248
rect 10781 25245 10793 25248
rect 10827 25245 10839 25279
rect 10781 25239 10839 25245
rect 38378 25236 38384 25288
rect 38436 25236 38442 25288
rect 17310 25168 17316 25220
rect 17368 25208 17374 25220
rect 17862 25208 17868 25220
rect 17368 25180 17868 25208
rect 17368 25168 17374 25180
rect 17862 25168 17868 25180
rect 17920 25168 17926 25220
rect 31478 25168 31484 25220
rect 31536 25208 31542 25220
rect 37553 25211 37611 25217
rect 37553 25208 37565 25211
rect 31536 25180 37565 25208
rect 31536 25168 31542 25180
rect 37553 25177 37565 25180
rect 37599 25177 37611 25211
rect 37553 25171 37611 25177
rect 10321 25143 10379 25149
rect 10321 25109 10333 25143
rect 10367 25140 10379 25143
rect 19518 25140 19524 25152
rect 10367 25112 19524 25140
rect 10367 25109 10379 25112
rect 10321 25103 10379 25109
rect 19518 25100 19524 25112
rect 19576 25100 19582 25152
rect 1104 25050 40848 25072
rect 1104 24998 2610 25050
rect 2662 24998 2674 25050
rect 2726 24998 2738 25050
rect 2790 24998 2802 25050
rect 2854 24998 2866 25050
rect 2918 24998 7610 25050
rect 7662 24998 7674 25050
rect 7726 24998 7738 25050
rect 7790 24998 7802 25050
rect 7854 24998 7866 25050
rect 7918 24998 12610 25050
rect 12662 24998 12674 25050
rect 12726 24998 12738 25050
rect 12790 24998 12802 25050
rect 12854 24998 12866 25050
rect 12918 24998 17610 25050
rect 17662 24998 17674 25050
rect 17726 24998 17738 25050
rect 17790 24998 17802 25050
rect 17854 24998 17866 25050
rect 17918 24998 22610 25050
rect 22662 24998 22674 25050
rect 22726 24998 22738 25050
rect 22790 24998 22802 25050
rect 22854 24998 22866 25050
rect 22918 24998 27610 25050
rect 27662 24998 27674 25050
rect 27726 24998 27738 25050
rect 27790 24998 27802 25050
rect 27854 24998 27866 25050
rect 27918 24998 32610 25050
rect 32662 24998 32674 25050
rect 32726 24998 32738 25050
rect 32790 24998 32802 25050
rect 32854 24998 32866 25050
rect 32918 24998 37610 25050
rect 37662 24998 37674 25050
rect 37726 24998 37738 25050
rect 37790 24998 37802 25050
rect 37854 24998 37866 25050
rect 37918 24998 40848 25050
rect 1104 24976 40848 24998
rect 27522 24896 27528 24948
rect 27580 24896 27586 24948
rect 19904 24840 20116 24868
rect 3418 24760 3424 24812
rect 3476 24800 3482 24812
rect 5166 24800 5172 24812
rect 3476 24772 5172 24800
rect 3476 24760 3482 24772
rect 5166 24760 5172 24772
rect 5224 24760 5230 24812
rect 7653 24803 7711 24809
rect 7653 24769 7665 24803
rect 7699 24800 7711 24803
rect 8018 24800 8024 24812
rect 7699 24772 8024 24800
rect 7699 24769 7711 24772
rect 7653 24763 7711 24769
rect 8018 24760 8024 24772
rect 8076 24760 8082 24812
rect 10502 24760 10508 24812
rect 10560 24760 10566 24812
rect 10965 24803 11023 24809
rect 10965 24769 10977 24803
rect 11011 24769 11023 24803
rect 10965 24763 11023 24769
rect 18325 24803 18383 24809
rect 18325 24769 18337 24803
rect 18371 24800 18383 24803
rect 18598 24800 18604 24812
rect 18371 24772 18604 24800
rect 18371 24769 18383 24772
rect 18325 24763 18383 24769
rect 7282 24692 7288 24744
rect 7340 24732 7346 24744
rect 7466 24732 7472 24744
rect 7340 24704 7472 24732
rect 7340 24692 7346 24704
rect 7466 24692 7472 24704
rect 7524 24692 7530 24744
rect 10410 24624 10416 24676
rect 10468 24624 10474 24676
rect 10980 24664 11008 24763
rect 18598 24760 18604 24772
rect 18656 24800 18662 24812
rect 19904 24800 19932 24840
rect 18656 24772 19932 24800
rect 18656 24760 18662 24772
rect 19978 24760 19984 24812
rect 20036 24760 20042 24812
rect 20088 24800 20116 24840
rect 20530 24800 20536 24812
rect 20088 24772 20536 24800
rect 20530 24760 20536 24772
rect 20588 24760 20594 24812
rect 26326 24760 26332 24812
rect 26384 24800 26390 24812
rect 27430 24800 27436 24812
rect 26384 24772 27436 24800
rect 26384 24760 26390 24772
rect 27430 24760 27436 24772
rect 27488 24760 27494 24812
rect 11241 24735 11299 24741
rect 11241 24701 11253 24735
rect 11287 24732 11299 24735
rect 20714 24732 20720 24744
rect 11287 24704 20720 24732
rect 11287 24701 11299 24704
rect 11241 24695 11299 24701
rect 20714 24692 20720 24704
rect 20772 24692 20778 24744
rect 22370 24664 22376 24676
rect 10980 24636 22376 24664
rect 19996 24608 20024 24636
rect 22370 24624 22376 24636
rect 22428 24624 22434 24676
rect 7193 24599 7251 24605
rect 7193 24565 7205 24599
rect 7239 24596 7251 24599
rect 7282 24596 7288 24608
rect 7239 24568 7288 24596
rect 7239 24565 7251 24568
rect 7193 24559 7251 24565
rect 7282 24556 7288 24568
rect 7340 24556 7346 24608
rect 19978 24556 19984 24608
rect 20036 24556 20042 24608
rect 27338 24556 27344 24608
rect 27396 24596 27402 24608
rect 27540 24596 27568 24896
rect 38562 24760 38568 24812
rect 38620 24800 38626 24812
rect 39206 24800 39212 24812
rect 38620 24772 39212 24800
rect 38620 24760 38626 24772
rect 39206 24760 39212 24772
rect 39264 24760 39270 24812
rect 27614 24692 27620 24744
rect 27672 24732 27678 24744
rect 38286 24732 38292 24744
rect 27672 24704 38292 24732
rect 27672 24692 27678 24704
rect 38286 24692 38292 24704
rect 38344 24692 38350 24744
rect 27396 24568 27568 24596
rect 27396 24556 27402 24568
rect 1104 24506 40848 24528
rect 1104 24454 1950 24506
rect 2002 24454 2014 24506
rect 2066 24454 2078 24506
rect 2130 24454 2142 24506
rect 2194 24454 2206 24506
rect 2258 24454 6950 24506
rect 7002 24454 7014 24506
rect 7066 24454 7078 24506
rect 7130 24454 7142 24506
rect 7194 24454 7206 24506
rect 7258 24454 11950 24506
rect 12002 24454 12014 24506
rect 12066 24454 12078 24506
rect 12130 24454 12142 24506
rect 12194 24454 12206 24506
rect 12258 24454 16950 24506
rect 17002 24454 17014 24506
rect 17066 24454 17078 24506
rect 17130 24454 17142 24506
rect 17194 24454 17206 24506
rect 17258 24454 21950 24506
rect 22002 24454 22014 24506
rect 22066 24454 22078 24506
rect 22130 24454 22142 24506
rect 22194 24454 22206 24506
rect 22258 24454 26950 24506
rect 27002 24454 27014 24506
rect 27066 24454 27078 24506
rect 27130 24454 27142 24506
rect 27194 24454 27206 24506
rect 27258 24454 31950 24506
rect 32002 24454 32014 24506
rect 32066 24454 32078 24506
rect 32130 24454 32142 24506
rect 32194 24454 32206 24506
rect 32258 24454 36950 24506
rect 37002 24454 37014 24506
rect 37066 24454 37078 24506
rect 37130 24454 37142 24506
rect 37194 24454 37206 24506
rect 37258 24454 40848 24506
rect 1104 24432 40848 24454
rect 8110 24352 8116 24404
rect 8168 24392 8174 24404
rect 8294 24392 8300 24404
rect 8168 24364 8300 24392
rect 8168 24352 8174 24364
rect 8294 24352 8300 24364
rect 8352 24352 8358 24404
rect 10502 24352 10508 24404
rect 10560 24392 10566 24404
rect 24670 24392 24676 24404
rect 10560 24364 24676 24392
rect 10560 24352 10566 24364
rect 24670 24352 24676 24364
rect 24728 24352 24734 24404
rect 33689 24395 33747 24401
rect 33689 24361 33701 24395
rect 33735 24392 33747 24395
rect 36354 24392 36360 24404
rect 33735 24364 36360 24392
rect 33735 24361 33747 24364
rect 33689 24355 33747 24361
rect 36354 24352 36360 24364
rect 36412 24352 36418 24404
rect 1670 24284 1676 24336
rect 1728 24324 1734 24336
rect 4982 24324 4988 24336
rect 1728 24296 4988 24324
rect 1728 24284 1734 24296
rect 4982 24284 4988 24296
rect 5040 24284 5046 24336
rect 1762 24216 1768 24268
rect 1820 24256 1826 24268
rect 10962 24256 10968 24268
rect 1820 24228 10968 24256
rect 1820 24216 1826 24228
rect 10962 24216 10968 24228
rect 11020 24216 11026 24268
rect 18966 24216 18972 24268
rect 19024 24216 19030 24268
rect 7193 24191 7251 24197
rect 7193 24157 7205 24191
rect 7239 24188 7251 24191
rect 7466 24188 7472 24200
rect 7239 24160 7472 24188
rect 7239 24157 7251 24160
rect 7193 24151 7251 24157
rect 7466 24148 7472 24160
rect 7524 24148 7530 24200
rect 12342 24148 12348 24200
rect 12400 24188 12406 24200
rect 17773 24191 17831 24197
rect 17773 24188 17785 24191
rect 12400 24160 17785 24188
rect 12400 24148 12406 24160
rect 17773 24157 17785 24160
rect 17819 24157 17831 24191
rect 17773 24151 17831 24157
rect 18138 24148 18144 24200
rect 18196 24148 18202 24200
rect 18690 24148 18696 24200
rect 18748 24148 18754 24200
rect 23290 24148 23296 24200
rect 23348 24188 23354 24200
rect 33042 24188 33048 24200
rect 23348 24160 33048 24188
rect 23348 24148 23354 24160
rect 33042 24148 33048 24160
rect 33100 24148 33106 24200
rect 33410 24148 33416 24200
rect 33468 24148 33474 24200
rect 33505 24191 33563 24197
rect 33505 24157 33517 24191
rect 33551 24188 33563 24191
rect 34238 24188 34244 24200
rect 33551 24160 34244 24188
rect 33551 24157 33563 24160
rect 33505 24151 33563 24157
rect 34238 24148 34244 24160
rect 34296 24148 34302 24200
rect 8018 24080 8024 24132
rect 8076 24080 8082 24132
rect 26050 24080 26056 24132
rect 26108 24080 26114 24132
rect 26142 24080 26148 24132
rect 26200 24120 26206 24132
rect 26421 24123 26479 24129
rect 26421 24120 26433 24123
rect 26200 24092 26433 24120
rect 26200 24080 26206 24092
rect 26421 24089 26433 24092
rect 26467 24089 26479 24123
rect 26421 24083 26479 24089
rect 29638 24080 29644 24132
rect 29696 24120 29702 24132
rect 33689 24123 33747 24129
rect 33689 24120 33701 24123
rect 29696 24092 33701 24120
rect 29696 24080 29702 24092
rect 33689 24089 33701 24092
rect 33735 24120 33747 24123
rect 36538 24120 36544 24132
rect 33735 24092 36544 24120
rect 33735 24089 33747 24092
rect 33689 24083 33747 24089
rect 36538 24080 36544 24092
rect 36596 24080 36602 24132
rect 19150 24012 19156 24064
rect 19208 24052 19214 24064
rect 26237 24055 26295 24061
rect 26237 24052 26249 24055
rect 19208 24024 26249 24052
rect 19208 24012 19214 24024
rect 26237 24021 26249 24024
rect 26283 24021 26295 24055
rect 26237 24015 26295 24021
rect 26326 24012 26332 24064
rect 26384 24012 26390 24064
rect 26510 24012 26516 24064
rect 26568 24012 26574 24064
rect 1104 23962 40848 23984
rect 1104 23910 2610 23962
rect 2662 23910 2674 23962
rect 2726 23910 2738 23962
rect 2790 23910 2802 23962
rect 2854 23910 2866 23962
rect 2918 23910 7610 23962
rect 7662 23910 7674 23962
rect 7726 23910 7738 23962
rect 7790 23910 7802 23962
rect 7854 23910 7866 23962
rect 7918 23910 12610 23962
rect 12662 23910 12674 23962
rect 12726 23910 12738 23962
rect 12790 23910 12802 23962
rect 12854 23910 12866 23962
rect 12918 23910 17610 23962
rect 17662 23910 17674 23962
rect 17726 23910 17738 23962
rect 17790 23910 17802 23962
rect 17854 23910 17866 23962
rect 17918 23910 22610 23962
rect 22662 23910 22674 23962
rect 22726 23910 22738 23962
rect 22790 23910 22802 23962
rect 22854 23910 22866 23962
rect 22918 23910 27610 23962
rect 27662 23910 27674 23962
rect 27726 23910 27738 23962
rect 27790 23910 27802 23962
rect 27854 23910 27866 23962
rect 27918 23910 32610 23962
rect 32662 23910 32674 23962
rect 32726 23910 32738 23962
rect 32790 23910 32802 23962
rect 32854 23910 32866 23962
rect 32918 23910 37610 23962
rect 37662 23910 37674 23962
rect 37726 23910 37738 23962
rect 37790 23910 37802 23962
rect 37854 23910 37866 23962
rect 37918 23910 40848 23962
rect 1104 23888 40848 23910
rect 8294 23848 8300 23860
rect 6656 23820 8300 23848
rect 6656 23721 6684 23820
rect 8294 23808 8300 23820
rect 8352 23808 8358 23860
rect 25866 23808 25872 23860
rect 25924 23848 25930 23860
rect 26142 23848 26148 23860
rect 25924 23820 26148 23848
rect 25924 23808 25930 23820
rect 26142 23808 26148 23820
rect 26200 23848 26206 23860
rect 26326 23848 26332 23860
rect 26200 23820 26332 23848
rect 26200 23808 26206 23820
rect 26326 23808 26332 23820
rect 26384 23808 26390 23860
rect 6917 23783 6975 23789
rect 6917 23749 6929 23783
rect 6963 23780 6975 23783
rect 7466 23780 7472 23792
rect 6963 23752 7472 23780
rect 6963 23749 6975 23752
rect 6917 23743 6975 23749
rect 7466 23740 7472 23752
rect 7524 23740 7530 23792
rect 8110 23780 8116 23792
rect 7576 23752 8116 23780
rect 6641 23715 6699 23721
rect 6641 23681 6653 23715
rect 6687 23681 6699 23715
rect 6641 23675 6699 23681
rect 6825 23715 6883 23721
rect 6825 23681 6837 23715
rect 6871 23681 6883 23715
rect 6825 23675 6883 23681
rect 7061 23715 7119 23721
rect 7061 23681 7073 23715
rect 7107 23712 7119 23715
rect 7576 23712 7604 23752
rect 8110 23740 8116 23752
rect 8168 23740 8174 23792
rect 34885 23783 34943 23789
rect 34885 23749 34897 23783
rect 34931 23780 34943 23783
rect 35434 23780 35440 23792
rect 34931 23752 35440 23780
rect 34931 23749 34943 23752
rect 34885 23743 34943 23749
rect 35434 23740 35440 23752
rect 35492 23740 35498 23792
rect 7107 23684 7604 23712
rect 7653 23715 7711 23721
rect 7107 23681 7119 23684
rect 7061 23675 7119 23681
rect 7653 23681 7665 23715
rect 7699 23712 7711 23715
rect 7699 23684 12434 23712
rect 7699 23681 7711 23684
rect 7653 23675 7711 23681
rect 6840 23644 6868 23675
rect 7668 23644 7696 23675
rect 6840 23616 7696 23644
rect 7745 23647 7803 23653
rect 7745 23613 7757 23647
rect 7791 23644 7803 23647
rect 8294 23644 8300 23656
rect 7791 23616 8300 23644
rect 7791 23613 7803 23616
rect 7745 23607 7803 23613
rect 8294 23604 8300 23616
rect 8352 23604 8358 23656
rect 12406 23644 12434 23684
rect 24578 23672 24584 23724
rect 24636 23712 24642 23724
rect 33873 23715 33931 23721
rect 33873 23712 33885 23715
rect 24636 23684 33885 23712
rect 24636 23672 24642 23684
rect 33873 23681 33885 23684
rect 33919 23681 33931 23715
rect 33873 23675 33931 23681
rect 34238 23672 34244 23724
rect 34296 23672 34302 23724
rect 27522 23644 27528 23656
rect 12406 23616 27528 23644
rect 27522 23604 27528 23616
rect 27580 23604 27586 23656
rect 33042 23604 33048 23656
rect 33100 23644 33106 23656
rect 33965 23647 34023 23653
rect 33965 23644 33977 23647
rect 33100 23616 33977 23644
rect 33100 23604 33106 23616
rect 33965 23613 33977 23616
rect 34011 23613 34023 23647
rect 33965 23607 34023 23613
rect 34146 23604 34152 23656
rect 34204 23604 34210 23656
rect 7193 23579 7251 23585
rect 7193 23545 7205 23579
rect 7239 23576 7251 23579
rect 26326 23576 26332 23588
rect 7239 23548 26332 23576
rect 7239 23545 7251 23548
rect 7193 23539 7251 23545
rect 26326 23536 26332 23548
rect 26384 23536 26390 23588
rect 33778 23536 33784 23588
rect 33836 23576 33842 23588
rect 34164 23576 34192 23604
rect 33836 23548 34192 23576
rect 33836 23536 33842 23548
rect 8205 23511 8263 23517
rect 8205 23477 8217 23511
rect 8251 23508 8263 23511
rect 8478 23508 8484 23520
rect 8251 23480 8484 23508
rect 8251 23477 8263 23480
rect 8205 23471 8263 23477
rect 8478 23468 8484 23480
rect 8536 23468 8542 23520
rect 1104 23418 40848 23440
rect 1104 23366 1950 23418
rect 2002 23366 2014 23418
rect 2066 23366 2078 23418
rect 2130 23366 2142 23418
rect 2194 23366 2206 23418
rect 2258 23366 6950 23418
rect 7002 23366 7014 23418
rect 7066 23366 7078 23418
rect 7130 23366 7142 23418
rect 7194 23366 7206 23418
rect 7258 23366 11950 23418
rect 12002 23366 12014 23418
rect 12066 23366 12078 23418
rect 12130 23366 12142 23418
rect 12194 23366 12206 23418
rect 12258 23366 16950 23418
rect 17002 23366 17014 23418
rect 17066 23366 17078 23418
rect 17130 23366 17142 23418
rect 17194 23366 17206 23418
rect 17258 23366 21950 23418
rect 22002 23366 22014 23418
rect 22066 23366 22078 23418
rect 22130 23366 22142 23418
rect 22194 23366 22206 23418
rect 22258 23366 26950 23418
rect 27002 23366 27014 23418
rect 27066 23366 27078 23418
rect 27130 23366 27142 23418
rect 27194 23366 27206 23418
rect 27258 23366 31950 23418
rect 32002 23366 32014 23418
rect 32066 23366 32078 23418
rect 32130 23366 32142 23418
rect 32194 23366 32206 23418
rect 32258 23366 36950 23418
rect 37002 23366 37014 23418
rect 37066 23366 37078 23418
rect 37130 23366 37142 23418
rect 37194 23366 37206 23418
rect 37258 23366 40848 23418
rect 1104 23344 40848 23366
rect 3602 23264 3608 23316
rect 3660 23304 3666 23316
rect 3970 23304 3976 23316
rect 3660 23276 3976 23304
rect 3660 23264 3666 23276
rect 3970 23264 3976 23276
rect 4028 23264 4034 23316
rect 17310 23304 17316 23316
rect 6932 23276 17316 23304
rect 6733 23239 6791 23245
rect 6733 23205 6745 23239
rect 6779 23236 6791 23239
rect 6822 23236 6828 23248
rect 6779 23208 6828 23236
rect 6779 23205 6791 23208
rect 6733 23199 6791 23205
rect 6822 23196 6828 23208
rect 6880 23196 6886 23248
rect 6932 23109 6960 23276
rect 17310 23264 17316 23276
rect 17368 23264 17374 23316
rect 18322 23264 18328 23316
rect 18380 23304 18386 23316
rect 21726 23304 21732 23316
rect 18380 23276 21732 23304
rect 18380 23264 18386 23276
rect 21726 23264 21732 23276
rect 21784 23264 21790 23316
rect 8938 23236 8944 23248
rect 7300 23208 8944 23236
rect 7300 23109 7328 23208
rect 8938 23196 8944 23208
rect 8996 23196 9002 23248
rect 11698 23196 11704 23248
rect 11756 23236 11762 23248
rect 12250 23236 12256 23248
rect 11756 23208 12256 23236
rect 11756 23196 11762 23208
rect 12250 23196 12256 23208
rect 12308 23196 12314 23248
rect 8389 23171 8447 23177
rect 8389 23137 8401 23171
rect 8435 23168 8447 23171
rect 10318 23168 10324 23180
rect 8435 23140 10324 23168
rect 8435 23137 8447 23140
rect 8389 23131 8447 23137
rect 10318 23128 10324 23140
rect 10376 23128 10382 23180
rect 15010 23128 15016 23180
rect 15068 23168 15074 23180
rect 27430 23168 27436 23180
rect 15068 23140 27436 23168
rect 15068 23128 15074 23140
rect 27430 23128 27436 23140
rect 27488 23128 27494 23180
rect 6917 23103 6975 23109
rect 6917 23069 6929 23103
rect 6963 23069 6975 23103
rect 6917 23063 6975 23069
rect 7285 23103 7343 23109
rect 7285 23069 7297 23103
rect 7331 23069 7343 23103
rect 7285 23063 7343 23069
rect 7377 23103 7435 23109
rect 7377 23069 7389 23103
rect 7423 23069 7435 23103
rect 7377 23063 7435 23069
rect 8297 23103 8355 23109
rect 8297 23069 8309 23103
rect 8343 23100 8355 23103
rect 17954 23100 17960 23112
rect 8343 23072 17960 23100
rect 8343 23069 8355 23072
rect 8297 23063 8355 23069
rect 7392 23032 7420 23063
rect 17954 23060 17960 23072
rect 18012 23100 18018 23112
rect 18230 23100 18236 23112
rect 18012 23072 18236 23100
rect 18012 23060 18018 23072
rect 18230 23060 18236 23072
rect 18288 23060 18294 23112
rect 20625 23103 20683 23109
rect 20625 23069 20637 23103
rect 20671 23069 20683 23103
rect 20625 23063 20683 23069
rect 19886 23032 19892 23044
rect 7392 23004 19892 23032
rect 19886 22992 19892 23004
rect 19944 23032 19950 23044
rect 20640 23032 20668 23063
rect 19944 23004 20668 23032
rect 21177 23035 21235 23041
rect 19944 22992 19950 23004
rect 21177 23001 21189 23035
rect 21223 23032 21235 23035
rect 30374 23032 30380 23044
rect 21223 23004 30380 23032
rect 21223 23001 21235 23004
rect 21177 22995 21235 23001
rect 30374 22992 30380 23004
rect 30432 22992 30438 23044
rect 4982 22924 4988 22976
rect 5040 22964 5046 22976
rect 7929 22967 7987 22973
rect 7929 22964 7941 22967
rect 5040 22936 7941 22964
rect 5040 22924 5046 22936
rect 7929 22933 7941 22936
rect 7975 22933 7987 22967
rect 7929 22927 7987 22933
rect 8662 22924 8668 22976
rect 8720 22964 8726 22976
rect 8938 22964 8944 22976
rect 8720 22936 8944 22964
rect 8720 22924 8726 22936
rect 8938 22924 8944 22936
rect 8996 22924 9002 22976
rect 18230 22924 18236 22976
rect 18288 22964 18294 22976
rect 37366 22964 37372 22976
rect 18288 22936 37372 22964
rect 18288 22924 18294 22936
rect 37366 22924 37372 22936
rect 37424 22924 37430 22976
rect 1104 22874 40848 22896
rect 1104 22822 2610 22874
rect 2662 22822 2674 22874
rect 2726 22822 2738 22874
rect 2790 22822 2802 22874
rect 2854 22822 2866 22874
rect 2918 22822 7610 22874
rect 7662 22822 7674 22874
rect 7726 22822 7738 22874
rect 7790 22822 7802 22874
rect 7854 22822 7866 22874
rect 7918 22822 12610 22874
rect 12662 22822 12674 22874
rect 12726 22822 12738 22874
rect 12790 22822 12802 22874
rect 12854 22822 12866 22874
rect 12918 22822 17610 22874
rect 17662 22822 17674 22874
rect 17726 22822 17738 22874
rect 17790 22822 17802 22874
rect 17854 22822 17866 22874
rect 17918 22822 22610 22874
rect 22662 22822 22674 22874
rect 22726 22822 22738 22874
rect 22790 22822 22802 22874
rect 22854 22822 22866 22874
rect 22918 22822 27610 22874
rect 27662 22822 27674 22874
rect 27726 22822 27738 22874
rect 27790 22822 27802 22874
rect 27854 22822 27866 22874
rect 27918 22822 32610 22874
rect 32662 22822 32674 22874
rect 32726 22822 32738 22874
rect 32790 22822 32802 22874
rect 32854 22822 32866 22874
rect 32918 22822 37610 22874
rect 37662 22822 37674 22874
rect 37726 22822 37738 22874
rect 37790 22822 37802 22874
rect 37854 22822 37866 22874
rect 37918 22822 40848 22874
rect 1104 22800 40848 22822
rect 11606 22720 11612 22772
rect 11664 22760 11670 22772
rect 11701 22763 11759 22769
rect 11701 22760 11713 22763
rect 11664 22732 11713 22760
rect 11664 22720 11670 22732
rect 11701 22729 11713 22732
rect 11747 22729 11759 22763
rect 11701 22723 11759 22729
rect 11793 22763 11851 22769
rect 11793 22729 11805 22763
rect 11839 22760 11851 22763
rect 11974 22760 11980 22772
rect 11839 22732 11980 22760
rect 11839 22729 11851 22732
rect 11793 22723 11851 22729
rect 11974 22720 11980 22732
rect 12032 22720 12038 22772
rect 12360 22732 15148 22760
rect 1673 22695 1731 22701
rect 1673 22661 1685 22695
rect 1719 22692 1731 22695
rect 8662 22692 8668 22704
rect 1719 22664 8668 22692
rect 1719 22661 1731 22664
rect 1673 22655 1731 22661
rect 8662 22652 8668 22664
rect 8720 22652 8726 22704
rect 11054 22652 11060 22704
rect 11112 22692 11118 22704
rect 11885 22695 11943 22701
rect 11885 22692 11897 22695
rect 11112 22664 11897 22692
rect 11112 22652 11118 22664
rect 11885 22661 11897 22664
rect 11931 22661 11943 22695
rect 11885 22655 11943 22661
rect 12250 22652 12256 22704
rect 12308 22652 12314 22704
rect 842 22584 848 22636
rect 900 22624 906 22636
rect 1397 22627 1455 22633
rect 1397 22624 1409 22627
rect 900 22596 1409 22624
rect 900 22584 906 22596
rect 1397 22593 1409 22596
rect 1443 22593 1455 22627
rect 12360 22624 12388 22732
rect 14918 22652 14924 22704
rect 14976 22652 14982 22704
rect 15010 22652 15016 22704
rect 15068 22652 15074 22704
rect 15120 22692 15148 22732
rect 17402 22720 17408 22772
rect 17460 22760 17466 22772
rect 17862 22760 17868 22772
rect 17460 22732 17868 22760
rect 17460 22720 17466 22732
rect 17862 22720 17868 22732
rect 17920 22720 17926 22772
rect 17954 22720 17960 22772
rect 18012 22760 18018 22772
rect 37366 22760 37372 22772
rect 18012 22732 37372 22760
rect 18012 22720 18018 22732
rect 37366 22720 37372 22732
rect 37424 22720 37430 22772
rect 18322 22692 18328 22704
rect 15120 22664 18328 22692
rect 18322 22652 18328 22664
rect 18380 22652 18386 22704
rect 1397 22587 1455 22593
rect 12268 22596 12388 22624
rect 6638 22516 6644 22568
rect 6696 22556 6702 22568
rect 11517 22559 11575 22565
rect 11517 22556 11529 22559
rect 6696 22528 11529 22556
rect 6696 22516 6702 22528
rect 11517 22525 11529 22528
rect 11563 22556 11575 22559
rect 12268 22556 12296 22596
rect 14642 22584 14648 22636
rect 14700 22584 14706 22636
rect 17310 22584 17316 22636
rect 17368 22584 17374 22636
rect 17586 22584 17592 22636
rect 17644 22584 17650 22636
rect 18785 22627 18843 22633
rect 18785 22624 18797 22627
rect 18524 22596 18797 22624
rect 14507 22559 14565 22565
rect 14507 22556 14519 22559
rect 11563 22528 12296 22556
rect 12406 22528 14519 22556
rect 11563 22525 11575 22528
rect 11517 22519 11575 22525
rect 7466 22448 7472 22500
rect 7524 22488 7530 22500
rect 8386 22488 8392 22500
rect 7524 22460 8392 22488
rect 7524 22448 7530 22460
rect 8386 22448 8392 22460
rect 8444 22488 8450 22500
rect 11974 22488 11980 22500
rect 8444 22460 11980 22488
rect 8444 22448 8450 22460
rect 11974 22448 11980 22460
rect 12032 22448 12038 22500
rect 3602 22380 3608 22432
rect 3660 22420 3666 22432
rect 12406 22420 12434 22528
rect 14507 22525 14519 22528
rect 14553 22525 14565 22559
rect 14507 22519 14565 22525
rect 14274 22448 14280 22500
rect 14332 22488 14338 22500
rect 16669 22491 16727 22497
rect 16669 22488 16681 22491
rect 14332 22460 16681 22488
rect 14332 22448 14338 22460
rect 16669 22457 16681 22460
rect 16715 22488 16727 22491
rect 18524 22488 18552 22596
rect 18785 22593 18797 22596
rect 18831 22593 18843 22627
rect 18785 22587 18843 22593
rect 40494 22584 40500 22636
rect 40552 22584 40558 22636
rect 19337 22559 19395 22565
rect 19337 22525 19349 22559
rect 19383 22556 19395 22559
rect 32950 22556 32956 22568
rect 19383 22528 32956 22556
rect 19383 22525 19395 22528
rect 19337 22519 19395 22525
rect 32950 22516 32956 22528
rect 33008 22516 33014 22568
rect 38838 22516 38844 22568
rect 38896 22556 38902 22568
rect 39669 22559 39727 22565
rect 39669 22556 39681 22559
rect 38896 22528 39681 22556
rect 38896 22516 38902 22528
rect 39669 22525 39681 22528
rect 39715 22525 39727 22559
rect 39669 22519 39727 22525
rect 16715 22460 18552 22488
rect 16715 22457 16727 22460
rect 16669 22451 16727 22457
rect 3660 22392 12434 22420
rect 3660 22380 3666 22392
rect 14366 22380 14372 22432
rect 14424 22380 14430 22432
rect 1104 22330 40848 22352
rect 1104 22278 1950 22330
rect 2002 22278 2014 22330
rect 2066 22278 2078 22330
rect 2130 22278 2142 22330
rect 2194 22278 2206 22330
rect 2258 22278 6950 22330
rect 7002 22278 7014 22330
rect 7066 22278 7078 22330
rect 7130 22278 7142 22330
rect 7194 22278 7206 22330
rect 7258 22278 11950 22330
rect 12002 22278 12014 22330
rect 12066 22278 12078 22330
rect 12130 22278 12142 22330
rect 12194 22278 12206 22330
rect 12258 22278 16950 22330
rect 17002 22278 17014 22330
rect 17066 22278 17078 22330
rect 17130 22278 17142 22330
rect 17194 22278 17206 22330
rect 17258 22278 21950 22330
rect 22002 22278 22014 22330
rect 22066 22278 22078 22330
rect 22130 22278 22142 22330
rect 22194 22278 22206 22330
rect 22258 22278 26950 22330
rect 27002 22278 27014 22330
rect 27066 22278 27078 22330
rect 27130 22278 27142 22330
rect 27194 22278 27206 22330
rect 27258 22278 31950 22330
rect 32002 22278 32014 22330
rect 32066 22278 32078 22330
rect 32130 22278 32142 22330
rect 32194 22278 32206 22330
rect 32258 22278 36950 22330
rect 37002 22278 37014 22330
rect 37066 22278 37078 22330
rect 37130 22278 37142 22330
rect 37194 22278 37206 22330
rect 37258 22278 40848 22330
rect 1104 22256 40848 22278
rect 17310 22176 17316 22228
rect 17368 22216 17374 22228
rect 17586 22216 17592 22228
rect 17368 22188 17592 22216
rect 17368 22176 17374 22188
rect 17586 22176 17592 22188
rect 17644 22176 17650 22228
rect 9030 22108 9036 22160
rect 9088 22148 9094 22160
rect 11606 22148 11612 22160
rect 9088 22120 11612 22148
rect 9088 22108 9094 22120
rect 11606 22108 11612 22120
rect 11664 22148 11670 22160
rect 18598 22148 18604 22160
rect 11664 22120 18604 22148
rect 11664 22108 11670 22120
rect 18598 22108 18604 22120
rect 18656 22108 18662 22160
rect 15286 22040 15292 22092
rect 15344 22040 15350 22092
rect 17218 22040 17224 22092
rect 17276 22080 17282 22092
rect 17402 22080 17408 22092
rect 17276 22052 17408 22080
rect 17276 22040 17282 22052
rect 17402 22040 17408 22052
rect 17460 22040 17466 22092
rect 25038 22040 25044 22092
rect 25096 22080 25102 22092
rect 26234 22080 26240 22092
rect 25096 22052 26240 22080
rect 25096 22040 25102 22052
rect 26234 22040 26240 22052
rect 26292 22040 26298 22092
rect 38838 22080 38844 22092
rect 35866 22052 38844 22080
rect 14826 21972 14832 22024
rect 14884 21972 14890 22024
rect 15013 22015 15071 22021
rect 15013 21981 15025 22015
rect 15059 22012 15071 22015
rect 26142 22012 26148 22024
rect 15059 21984 26148 22012
rect 15059 21981 15071 21984
rect 15013 21975 15071 21981
rect 14553 21947 14611 21953
rect 14553 21913 14565 21947
rect 14599 21944 14611 21947
rect 15028 21944 15056 21975
rect 26142 21972 26148 21984
rect 26200 22012 26206 22024
rect 35866 22012 35894 22052
rect 38838 22040 38844 22052
rect 38896 22040 38902 22092
rect 26200 21984 35894 22012
rect 26200 21972 26206 21984
rect 14599 21916 15056 21944
rect 14599 21913 14611 21916
rect 14553 21907 14611 21913
rect 17494 21836 17500 21888
rect 17552 21876 17558 21888
rect 17862 21876 17868 21888
rect 17552 21848 17868 21876
rect 17552 21836 17558 21848
rect 17862 21836 17868 21848
rect 17920 21836 17926 21888
rect 1104 21786 40848 21808
rect 1104 21734 2610 21786
rect 2662 21734 2674 21786
rect 2726 21734 2738 21786
rect 2790 21734 2802 21786
rect 2854 21734 2866 21786
rect 2918 21734 7610 21786
rect 7662 21734 7674 21786
rect 7726 21734 7738 21786
rect 7790 21734 7802 21786
rect 7854 21734 7866 21786
rect 7918 21734 12610 21786
rect 12662 21734 12674 21786
rect 12726 21734 12738 21786
rect 12790 21734 12802 21786
rect 12854 21734 12866 21786
rect 12918 21734 17610 21786
rect 17662 21734 17674 21786
rect 17726 21734 17738 21786
rect 17790 21734 17802 21786
rect 17854 21734 17866 21786
rect 17918 21734 22610 21786
rect 22662 21734 22674 21786
rect 22726 21734 22738 21786
rect 22790 21734 22802 21786
rect 22854 21734 22866 21786
rect 22918 21734 27610 21786
rect 27662 21734 27674 21786
rect 27726 21734 27738 21786
rect 27790 21734 27802 21786
rect 27854 21734 27866 21786
rect 27918 21734 32610 21786
rect 32662 21734 32674 21786
rect 32726 21734 32738 21786
rect 32790 21734 32802 21786
rect 32854 21734 32866 21786
rect 32918 21734 37610 21786
rect 37662 21734 37674 21786
rect 37726 21734 37738 21786
rect 37790 21734 37802 21786
rect 37854 21734 37866 21786
rect 37918 21734 40848 21786
rect 1104 21712 40848 21734
rect 31754 21428 31760 21480
rect 31812 21468 31818 21480
rect 39022 21468 39028 21480
rect 31812 21440 39028 21468
rect 31812 21428 31818 21440
rect 39022 21428 39028 21440
rect 39080 21428 39086 21480
rect 11698 21360 11704 21412
rect 11756 21400 11762 21412
rect 12434 21400 12440 21412
rect 11756 21372 12440 21400
rect 11756 21360 11762 21372
rect 12434 21360 12440 21372
rect 12492 21360 12498 21412
rect 17218 21360 17224 21412
rect 17276 21400 17282 21412
rect 38470 21400 38476 21412
rect 17276 21372 38476 21400
rect 17276 21360 17282 21372
rect 38470 21360 38476 21372
rect 38528 21360 38534 21412
rect 7834 21292 7840 21344
rect 7892 21332 7898 21344
rect 33226 21332 33232 21344
rect 7892 21304 33232 21332
rect 7892 21292 7898 21304
rect 33226 21292 33232 21304
rect 33284 21292 33290 21344
rect 1104 21242 40848 21264
rect 1104 21190 1950 21242
rect 2002 21190 2014 21242
rect 2066 21190 2078 21242
rect 2130 21190 2142 21242
rect 2194 21190 2206 21242
rect 2258 21190 6950 21242
rect 7002 21190 7014 21242
rect 7066 21190 7078 21242
rect 7130 21190 7142 21242
rect 7194 21190 7206 21242
rect 7258 21190 11950 21242
rect 12002 21190 12014 21242
rect 12066 21190 12078 21242
rect 12130 21190 12142 21242
rect 12194 21190 12206 21242
rect 12258 21190 16950 21242
rect 17002 21190 17014 21242
rect 17066 21190 17078 21242
rect 17130 21190 17142 21242
rect 17194 21190 17206 21242
rect 17258 21190 21950 21242
rect 22002 21190 22014 21242
rect 22066 21190 22078 21242
rect 22130 21190 22142 21242
rect 22194 21190 22206 21242
rect 22258 21190 26950 21242
rect 27002 21190 27014 21242
rect 27066 21190 27078 21242
rect 27130 21190 27142 21242
rect 27194 21190 27206 21242
rect 27258 21190 31950 21242
rect 32002 21190 32014 21242
rect 32066 21190 32078 21242
rect 32130 21190 32142 21242
rect 32194 21190 32206 21242
rect 32258 21190 36950 21242
rect 37002 21190 37014 21242
rect 37066 21190 37078 21242
rect 37130 21190 37142 21242
rect 37194 21190 37206 21242
rect 37258 21190 40848 21242
rect 1104 21168 40848 21190
rect 12986 21128 12992 21140
rect 3252 21100 12992 21128
rect 3252 20933 3280 21100
rect 12986 21088 12992 21100
rect 13044 21128 13050 21140
rect 13044 21100 16068 21128
rect 13044 21088 13050 21100
rect 15930 21060 15936 21072
rect 7116 21032 15936 21060
rect 7116 21001 7144 21032
rect 15930 21020 15936 21032
rect 15988 21020 15994 21072
rect 7101 20995 7159 21001
rect 7101 20961 7113 20995
rect 7147 20961 7159 20995
rect 10594 20992 10600 21004
rect 7101 20955 7159 20961
rect 7484 20964 10600 20992
rect 3145 20927 3203 20933
rect 3145 20893 3157 20927
rect 3191 20893 3203 20927
rect 3145 20887 3203 20893
rect 3237 20927 3295 20933
rect 3237 20893 3249 20927
rect 3283 20893 3295 20927
rect 3237 20887 3295 20893
rect 3160 20856 3188 20887
rect 3418 20884 3424 20936
rect 3476 20884 3482 20936
rect 3510 20884 3516 20936
rect 3568 20884 3574 20936
rect 7484 20933 7512 20964
rect 10594 20952 10600 20964
rect 10652 20952 10658 21004
rect 7469 20927 7527 20933
rect 7469 20893 7481 20927
rect 7515 20893 7527 20927
rect 7469 20887 7527 20893
rect 7834 20884 7840 20936
rect 7892 20884 7898 20936
rect 4982 20856 4988 20868
rect 3160 20828 4988 20856
rect 4982 20816 4988 20828
rect 5040 20816 5046 20868
rect 8021 20859 8079 20865
rect 8021 20825 8033 20859
rect 8067 20856 8079 20859
rect 9306 20856 9312 20868
rect 8067 20828 9312 20856
rect 8067 20825 8079 20828
rect 8021 20819 8079 20825
rect 9306 20816 9312 20828
rect 9364 20816 9370 20868
rect 16040 20856 16068 21100
rect 22462 21060 22468 21072
rect 22112 21032 22468 21060
rect 22112 21001 22140 21032
rect 22462 21020 22468 21032
rect 22520 21020 22526 21072
rect 22097 20995 22155 21001
rect 22097 20961 22109 20995
rect 22143 20961 22155 20995
rect 22097 20955 22155 20961
rect 22278 20952 22284 21004
rect 22336 20952 22342 21004
rect 23017 20995 23075 21001
rect 23017 20961 23029 20995
rect 23063 20992 23075 20995
rect 24026 20992 24032 21004
rect 23063 20964 24032 20992
rect 23063 20961 23075 20964
rect 23017 20955 23075 20961
rect 24026 20952 24032 20964
rect 24084 20952 24090 21004
rect 21818 20884 21824 20936
rect 21876 20924 21882 20936
rect 22005 20927 22063 20933
rect 22005 20924 22017 20927
rect 21876 20896 22017 20924
rect 21876 20884 21882 20896
rect 22005 20893 22017 20896
rect 22051 20893 22063 20927
rect 22005 20887 22063 20893
rect 22370 20884 22376 20936
rect 22428 20884 22434 20936
rect 27338 20856 27344 20868
rect 16040 20828 27344 20856
rect 27338 20816 27344 20828
rect 27396 20816 27402 20868
rect 2961 20791 3019 20797
rect 2961 20757 2973 20791
rect 3007 20788 3019 20791
rect 4798 20788 4804 20800
rect 3007 20760 4804 20788
rect 3007 20757 3019 20760
rect 2961 20751 3019 20757
rect 4798 20748 4804 20760
rect 4856 20748 4862 20800
rect 1104 20698 40848 20720
rect 1104 20646 2610 20698
rect 2662 20646 2674 20698
rect 2726 20646 2738 20698
rect 2790 20646 2802 20698
rect 2854 20646 2866 20698
rect 2918 20646 7610 20698
rect 7662 20646 7674 20698
rect 7726 20646 7738 20698
rect 7790 20646 7802 20698
rect 7854 20646 7866 20698
rect 7918 20646 12610 20698
rect 12662 20646 12674 20698
rect 12726 20646 12738 20698
rect 12790 20646 12802 20698
rect 12854 20646 12866 20698
rect 12918 20646 17610 20698
rect 17662 20646 17674 20698
rect 17726 20646 17738 20698
rect 17790 20646 17802 20698
rect 17854 20646 17866 20698
rect 17918 20646 22610 20698
rect 22662 20646 22674 20698
rect 22726 20646 22738 20698
rect 22790 20646 22802 20698
rect 22854 20646 22866 20698
rect 22918 20646 27610 20698
rect 27662 20646 27674 20698
rect 27726 20646 27738 20698
rect 27790 20646 27802 20698
rect 27854 20646 27866 20698
rect 27918 20646 32610 20698
rect 32662 20646 32674 20698
rect 32726 20646 32738 20698
rect 32790 20646 32802 20698
rect 32854 20646 32866 20698
rect 32918 20646 37610 20698
rect 37662 20646 37674 20698
rect 37726 20646 37738 20698
rect 37790 20646 37802 20698
rect 37854 20646 37866 20698
rect 37918 20646 40848 20698
rect 1104 20624 40848 20646
rect 1670 20544 1676 20596
rect 1728 20544 1734 20596
rect 20622 20544 20628 20596
rect 20680 20584 20686 20596
rect 24857 20587 24915 20593
rect 20680 20556 24808 20584
rect 20680 20544 20686 20556
rect 1578 20476 1584 20528
rect 1636 20516 1642 20528
rect 1949 20519 2007 20525
rect 1949 20516 1961 20519
rect 1636 20488 1961 20516
rect 1636 20476 1642 20488
rect 1949 20485 1961 20488
rect 1995 20485 2007 20519
rect 1949 20479 2007 20485
rect 23014 20476 23020 20528
rect 23072 20516 23078 20528
rect 24780 20516 24808 20556
rect 24857 20553 24869 20587
rect 24903 20584 24915 20587
rect 24946 20584 24952 20596
rect 24903 20556 24952 20584
rect 24903 20553 24915 20556
rect 24857 20547 24915 20553
rect 24946 20544 24952 20556
rect 25004 20544 25010 20596
rect 37458 20584 37464 20596
rect 26206 20556 37464 20584
rect 26206 20516 26234 20556
rect 37458 20544 37464 20556
rect 37516 20544 37522 20596
rect 23072 20488 24440 20516
rect 24780 20488 26234 20516
rect 33137 20519 33195 20525
rect 23072 20476 23078 20488
rect 1765 20451 1823 20457
rect 1765 20417 1777 20451
rect 1811 20448 1823 20451
rect 5074 20448 5080 20460
rect 1811 20420 5080 20448
rect 1811 20417 1823 20420
rect 1765 20411 1823 20417
rect 5074 20408 5080 20420
rect 5132 20408 5138 20460
rect 24118 20408 24124 20460
rect 24176 20408 24182 20460
rect 24305 20451 24363 20457
rect 24305 20417 24317 20451
rect 24351 20417 24363 20451
rect 24412 20448 24440 20488
rect 33137 20485 33149 20519
rect 33183 20516 33195 20519
rect 35710 20516 35716 20528
rect 33183 20488 35716 20516
rect 33183 20485 33195 20488
rect 33137 20479 33195 20485
rect 35710 20476 35716 20488
rect 35768 20476 35774 20528
rect 24765 20451 24823 20457
rect 24765 20448 24777 20451
rect 24412 20420 24777 20448
rect 24305 20411 24363 20417
rect 24765 20417 24777 20420
rect 24811 20417 24823 20451
rect 24765 20411 24823 20417
rect 25317 20451 25375 20457
rect 25317 20417 25329 20451
rect 25363 20417 25375 20451
rect 25317 20411 25375 20417
rect 22370 20340 22376 20392
rect 22428 20380 22434 20392
rect 23290 20380 23296 20392
rect 22428 20352 23296 20380
rect 22428 20340 22434 20352
rect 23290 20340 23296 20352
rect 23348 20380 23354 20392
rect 24320 20380 24348 20411
rect 23348 20352 24348 20380
rect 23348 20340 23354 20352
rect 24670 20340 24676 20392
rect 24728 20340 24734 20392
rect 24578 20272 24584 20324
rect 24636 20272 24642 20324
rect 23290 20204 23296 20256
rect 23348 20244 23354 20256
rect 25332 20244 25360 20411
rect 27338 20408 27344 20460
rect 27396 20448 27402 20460
rect 33321 20451 33379 20457
rect 33321 20448 33333 20451
rect 27396 20420 33333 20448
rect 27396 20408 27402 20420
rect 33321 20417 33333 20420
rect 33367 20417 33379 20451
rect 33321 20411 33379 20417
rect 33413 20451 33471 20457
rect 33413 20417 33425 20451
rect 33459 20448 33471 20451
rect 34974 20448 34980 20460
rect 33459 20420 34980 20448
rect 33459 20417 33471 20420
rect 33413 20411 33471 20417
rect 25777 20383 25835 20389
rect 25777 20349 25789 20383
rect 25823 20380 25835 20383
rect 33336 20380 33364 20411
rect 34974 20408 34980 20420
rect 35032 20408 35038 20460
rect 35066 20380 35072 20392
rect 25823 20352 33272 20380
rect 33336 20352 35072 20380
rect 25823 20349 25835 20352
rect 25777 20343 25835 20349
rect 23348 20216 25360 20244
rect 23348 20204 23354 20216
rect 33134 20204 33140 20256
rect 33192 20204 33198 20256
rect 33244 20244 33272 20352
rect 35066 20340 35072 20352
rect 35124 20340 35130 20392
rect 35158 20244 35164 20256
rect 33244 20216 35164 20244
rect 35158 20204 35164 20216
rect 35216 20204 35222 20256
rect 1104 20154 40848 20176
rect 1104 20102 1950 20154
rect 2002 20102 2014 20154
rect 2066 20102 2078 20154
rect 2130 20102 2142 20154
rect 2194 20102 2206 20154
rect 2258 20102 6950 20154
rect 7002 20102 7014 20154
rect 7066 20102 7078 20154
rect 7130 20102 7142 20154
rect 7194 20102 7206 20154
rect 7258 20102 11950 20154
rect 12002 20102 12014 20154
rect 12066 20102 12078 20154
rect 12130 20102 12142 20154
rect 12194 20102 12206 20154
rect 12258 20102 16950 20154
rect 17002 20102 17014 20154
rect 17066 20102 17078 20154
rect 17130 20102 17142 20154
rect 17194 20102 17206 20154
rect 17258 20102 21950 20154
rect 22002 20102 22014 20154
rect 22066 20102 22078 20154
rect 22130 20102 22142 20154
rect 22194 20102 22206 20154
rect 22258 20102 26950 20154
rect 27002 20102 27014 20154
rect 27066 20102 27078 20154
rect 27130 20102 27142 20154
rect 27194 20102 27206 20154
rect 27258 20102 31950 20154
rect 32002 20102 32014 20154
rect 32066 20102 32078 20154
rect 32130 20102 32142 20154
rect 32194 20102 32206 20154
rect 32258 20102 36950 20154
rect 37002 20102 37014 20154
rect 37066 20102 37078 20154
rect 37130 20102 37142 20154
rect 37194 20102 37206 20154
rect 37258 20102 40848 20154
rect 1104 20080 40848 20102
rect 18414 20000 18420 20052
rect 18472 20040 18478 20052
rect 27338 20040 27344 20052
rect 18472 20012 27344 20040
rect 18472 20000 18478 20012
rect 27338 20000 27344 20012
rect 27396 20000 27402 20052
rect 33226 20000 33232 20052
rect 33284 20040 33290 20052
rect 33502 20040 33508 20052
rect 33284 20012 33508 20040
rect 33284 20000 33290 20012
rect 33502 20000 33508 20012
rect 33560 20000 33566 20052
rect 4614 19972 4620 19984
rect 4080 19944 4620 19972
rect 4080 19845 4108 19944
rect 4614 19932 4620 19944
rect 4672 19932 4678 19984
rect 19518 19932 19524 19984
rect 19576 19972 19582 19984
rect 19576 19944 37964 19972
rect 19576 19932 19582 19944
rect 4157 19907 4215 19913
rect 4157 19873 4169 19907
rect 4203 19904 4215 19907
rect 7561 19907 7619 19913
rect 4203 19876 6914 19904
rect 4203 19873 4215 19876
rect 4157 19867 4215 19873
rect 4065 19839 4123 19845
rect 4065 19805 4077 19839
rect 4111 19805 4123 19839
rect 4065 19799 4123 19805
rect 4338 19796 4344 19848
rect 4396 19796 4402 19848
rect 6886 19836 6914 19876
rect 7561 19873 7573 19907
rect 7607 19904 7619 19907
rect 8018 19904 8024 19916
rect 7607 19876 8024 19904
rect 7607 19873 7619 19876
rect 7561 19867 7619 19873
rect 8018 19864 8024 19876
rect 8076 19864 8082 19916
rect 13170 19904 13176 19916
rect 12406 19876 13176 19904
rect 12406 19836 12434 19876
rect 13170 19864 13176 19876
rect 13228 19904 13234 19916
rect 18230 19904 18236 19916
rect 13228 19876 18236 19904
rect 13228 19864 13234 19876
rect 18230 19864 18236 19876
rect 18288 19864 18294 19916
rect 37458 19864 37464 19916
rect 37516 19864 37522 19916
rect 6886 19808 12434 19836
rect 15746 19796 15752 19848
rect 15804 19796 15810 19848
rect 33226 19796 33232 19848
rect 33284 19796 33290 19848
rect 33318 19796 33324 19848
rect 33376 19836 33382 19848
rect 33781 19839 33839 19845
rect 33781 19836 33793 19839
rect 33376 19808 33793 19836
rect 33376 19796 33382 19808
rect 33781 19805 33793 19808
rect 33827 19805 33839 19839
rect 33781 19799 33839 19805
rect 37366 19796 37372 19848
rect 37424 19836 37430 19848
rect 37936 19845 37964 19944
rect 38010 19932 38016 19984
rect 38068 19972 38074 19984
rect 38105 19975 38163 19981
rect 38105 19972 38117 19975
rect 38068 19944 38117 19972
rect 38068 19932 38074 19944
rect 38105 19941 38117 19944
rect 38151 19941 38163 19975
rect 38105 19935 38163 19941
rect 37553 19839 37611 19845
rect 37553 19836 37565 19839
rect 37424 19808 37565 19836
rect 37424 19796 37430 19808
rect 37553 19805 37565 19808
rect 37599 19805 37611 19839
rect 37553 19799 37611 19805
rect 37921 19839 37979 19845
rect 37921 19805 37933 19839
rect 37967 19805 37979 19839
rect 37921 19799 37979 19805
rect 16945 19771 17003 19777
rect 16945 19737 16957 19771
rect 16991 19768 17003 19771
rect 17402 19768 17408 19780
rect 16991 19740 17408 19768
rect 16991 19737 17003 19740
rect 16945 19731 17003 19737
rect 17402 19728 17408 19740
rect 17460 19728 17466 19780
rect 18506 19728 18512 19780
rect 18564 19768 18570 19780
rect 18690 19768 18696 19780
rect 18564 19740 18696 19768
rect 18564 19728 18570 19740
rect 18690 19728 18696 19740
rect 18748 19768 18754 19780
rect 18748 19740 33626 19768
rect 18748 19728 18754 19740
rect 6270 19660 6276 19712
rect 6328 19700 6334 19712
rect 7101 19703 7159 19709
rect 7101 19700 7113 19703
rect 6328 19672 7113 19700
rect 6328 19660 6334 19672
rect 7101 19669 7113 19672
rect 7147 19669 7159 19703
rect 7101 19663 7159 19669
rect 7190 19660 7196 19712
rect 7248 19700 7254 19712
rect 8110 19700 8116 19712
rect 7248 19672 8116 19700
rect 7248 19660 7254 19672
rect 8110 19660 8116 19672
rect 8168 19700 8174 19712
rect 30834 19700 30840 19712
rect 8168 19672 30840 19700
rect 8168 19660 8174 19672
rect 30834 19660 30840 19672
rect 30892 19660 30898 19712
rect 33226 19660 33232 19712
rect 33284 19700 33290 19712
rect 33778 19700 33784 19712
rect 33284 19672 33784 19700
rect 33284 19660 33290 19672
rect 33778 19660 33784 19672
rect 33836 19660 33842 19712
rect 1104 19610 40848 19632
rect 1104 19558 2610 19610
rect 2662 19558 2674 19610
rect 2726 19558 2738 19610
rect 2790 19558 2802 19610
rect 2854 19558 2866 19610
rect 2918 19558 7610 19610
rect 7662 19558 7674 19610
rect 7726 19558 7738 19610
rect 7790 19558 7802 19610
rect 7854 19558 7866 19610
rect 7918 19558 12610 19610
rect 12662 19558 12674 19610
rect 12726 19558 12738 19610
rect 12790 19558 12802 19610
rect 12854 19558 12866 19610
rect 12918 19558 17610 19610
rect 17662 19558 17674 19610
rect 17726 19558 17738 19610
rect 17790 19558 17802 19610
rect 17854 19558 17866 19610
rect 17918 19558 22610 19610
rect 22662 19558 22674 19610
rect 22726 19558 22738 19610
rect 22790 19558 22802 19610
rect 22854 19558 22866 19610
rect 22918 19558 27610 19610
rect 27662 19558 27674 19610
rect 27726 19558 27738 19610
rect 27790 19558 27802 19610
rect 27854 19558 27866 19610
rect 27918 19558 32610 19610
rect 32662 19558 32674 19610
rect 32726 19558 32738 19610
rect 32790 19558 32802 19610
rect 32854 19558 32866 19610
rect 32918 19558 37610 19610
rect 37662 19558 37674 19610
rect 37726 19558 37738 19610
rect 37790 19558 37802 19610
rect 37854 19558 37866 19610
rect 37918 19558 40848 19610
rect 1104 19536 40848 19558
rect 18966 19496 18972 19508
rect 7576 19468 18972 19496
rect 7576 19428 7604 19468
rect 18966 19456 18972 19468
rect 19024 19456 19030 19508
rect 24670 19456 24676 19508
rect 24728 19496 24734 19508
rect 33134 19496 33140 19508
rect 24728 19468 33140 19496
rect 24728 19456 24734 19468
rect 33134 19456 33140 19468
rect 33192 19456 33198 19508
rect 7484 19400 7604 19428
rect 7101 19363 7159 19369
rect 7101 19329 7113 19363
rect 7147 19360 7159 19363
rect 7190 19360 7196 19372
rect 7147 19332 7196 19360
rect 7147 19329 7159 19332
rect 7101 19323 7159 19329
rect 7190 19320 7196 19332
rect 7248 19320 7254 19372
rect 7484 19369 7512 19400
rect 8018 19388 8024 19440
rect 8076 19428 8082 19440
rect 13541 19431 13599 19437
rect 8076 19400 12434 19428
rect 8076 19388 8082 19400
rect 7469 19363 7527 19369
rect 7469 19329 7481 19363
rect 7515 19329 7527 19363
rect 7469 19323 7527 19329
rect 7837 19363 7895 19369
rect 7837 19329 7849 19363
rect 7883 19360 7895 19363
rect 9490 19360 9496 19372
rect 7883 19332 9496 19360
rect 7883 19329 7895 19332
rect 7837 19323 7895 19329
rect 9490 19320 9496 19332
rect 9548 19320 9554 19372
rect 12406 19360 12434 19400
rect 13541 19397 13553 19431
rect 13587 19428 13599 19431
rect 18414 19428 18420 19440
rect 13587 19400 18420 19428
rect 13587 19397 13599 19400
rect 13541 19391 13599 19397
rect 18414 19388 18420 19400
rect 18472 19388 18478 19440
rect 12897 19363 12955 19369
rect 12897 19360 12909 19363
rect 12406 19332 12909 19360
rect 12897 19329 12909 19332
rect 12943 19360 12955 19363
rect 18690 19360 18696 19372
rect 12943 19332 18696 19360
rect 12943 19329 12955 19332
rect 12897 19323 12955 19329
rect 18690 19320 18696 19332
rect 18748 19320 18754 19372
rect 7745 19295 7803 19301
rect 7745 19261 7757 19295
rect 7791 19292 7803 19295
rect 8018 19292 8024 19304
rect 7791 19264 8024 19292
rect 7791 19261 7803 19264
rect 7745 19255 7803 19261
rect 8018 19252 8024 19264
rect 8076 19292 8082 19304
rect 8202 19292 8208 19304
rect 8076 19264 8208 19292
rect 8076 19252 8082 19264
rect 8202 19252 8208 19264
rect 8260 19252 8266 19304
rect 17862 19116 17868 19168
rect 17920 19156 17926 19168
rect 22278 19156 22284 19168
rect 17920 19128 22284 19156
rect 17920 19116 17926 19128
rect 22278 19116 22284 19128
rect 22336 19116 22342 19168
rect 1104 19066 40848 19088
rect 1104 19014 1950 19066
rect 2002 19014 2014 19066
rect 2066 19014 2078 19066
rect 2130 19014 2142 19066
rect 2194 19014 2206 19066
rect 2258 19014 6950 19066
rect 7002 19014 7014 19066
rect 7066 19014 7078 19066
rect 7130 19014 7142 19066
rect 7194 19014 7206 19066
rect 7258 19014 11950 19066
rect 12002 19014 12014 19066
rect 12066 19014 12078 19066
rect 12130 19014 12142 19066
rect 12194 19014 12206 19066
rect 12258 19014 16950 19066
rect 17002 19014 17014 19066
rect 17066 19014 17078 19066
rect 17130 19014 17142 19066
rect 17194 19014 17206 19066
rect 17258 19014 21950 19066
rect 22002 19014 22014 19066
rect 22066 19014 22078 19066
rect 22130 19014 22142 19066
rect 22194 19014 22206 19066
rect 22258 19014 26950 19066
rect 27002 19014 27014 19066
rect 27066 19014 27078 19066
rect 27130 19014 27142 19066
rect 27194 19014 27206 19066
rect 27258 19014 31950 19066
rect 32002 19014 32014 19066
rect 32066 19014 32078 19066
rect 32130 19014 32142 19066
rect 32194 19014 32206 19066
rect 32258 19014 36950 19066
rect 37002 19014 37014 19066
rect 37066 19014 37078 19066
rect 37130 19014 37142 19066
rect 37194 19014 37206 19066
rect 37258 19014 40848 19066
rect 1104 18992 40848 19014
rect 17589 18887 17647 18893
rect 17589 18884 17601 18887
rect 12406 18856 17601 18884
rect 10962 18776 10968 18828
rect 11020 18816 11026 18828
rect 12406 18816 12434 18856
rect 17589 18853 17601 18856
rect 17635 18853 17647 18887
rect 17589 18847 17647 18853
rect 11020 18788 12434 18816
rect 11020 18776 11026 18788
rect 17604 18680 17632 18847
rect 25590 18844 25596 18896
rect 25648 18884 25654 18896
rect 25648 18856 26234 18884
rect 25648 18844 25654 18856
rect 21082 18776 21088 18828
rect 21140 18816 21146 18828
rect 25777 18819 25835 18825
rect 25777 18816 25789 18819
rect 21140 18788 25789 18816
rect 21140 18776 21146 18788
rect 25777 18785 25789 18788
rect 25823 18785 25835 18819
rect 26206 18816 26234 18856
rect 26697 18819 26755 18825
rect 26697 18816 26709 18819
rect 26206 18788 26709 18816
rect 25777 18779 25835 18785
rect 26697 18785 26709 18788
rect 26743 18785 26755 18819
rect 26697 18779 26755 18785
rect 17862 18708 17868 18760
rect 17920 18708 17926 18760
rect 18414 18708 18420 18760
rect 18472 18748 18478 18760
rect 18598 18748 18604 18760
rect 18472 18720 18604 18748
rect 18472 18708 18478 18720
rect 18598 18708 18604 18720
rect 18656 18708 18662 18760
rect 18690 18708 18696 18760
rect 18748 18748 18754 18760
rect 19245 18751 19303 18757
rect 19245 18748 19257 18751
rect 18748 18720 19257 18748
rect 18748 18708 18754 18720
rect 19245 18717 19257 18720
rect 19291 18717 19303 18751
rect 19245 18711 19303 18717
rect 26234 18708 26240 18760
rect 26292 18708 26298 18760
rect 26418 18708 26424 18760
rect 26476 18708 26482 18760
rect 26602 18708 26608 18760
rect 26660 18748 26666 18760
rect 26789 18751 26847 18757
rect 26789 18748 26801 18751
rect 26660 18720 26801 18748
rect 26660 18708 26666 18720
rect 26789 18717 26801 18720
rect 26835 18717 26847 18751
rect 26789 18711 26847 18717
rect 30926 18680 30932 18692
rect 17604 18652 30932 18680
rect 30926 18640 30932 18652
rect 30984 18640 30990 18692
rect 19429 18615 19487 18621
rect 19429 18581 19441 18615
rect 19475 18612 19487 18615
rect 19518 18612 19524 18624
rect 19475 18584 19524 18612
rect 19475 18581 19487 18584
rect 19429 18575 19487 18581
rect 19518 18572 19524 18584
rect 19576 18572 19582 18624
rect 1104 18522 40848 18544
rect 1104 18470 2610 18522
rect 2662 18470 2674 18522
rect 2726 18470 2738 18522
rect 2790 18470 2802 18522
rect 2854 18470 2866 18522
rect 2918 18470 7610 18522
rect 7662 18470 7674 18522
rect 7726 18470 7738 18522
rect 7790 18470 7802 18522
rect 7854 18470 7866 18522
rect 7918 18470 12610 18522
rect 12662 18470 12674 18522
rect 12726 18470 12738 18522
rect 12790 18470 12802 18522
rect 12854 18470 12866 18522
rect 12918 18470 17610 18522
rect 17662 18470 17674 18522
rect 17726 18470 17738 18522
rect 17790 18470 17802 18522
rect 17854 18470 17866 18522
rect 17918 18470 22610 18522
rect 22662 18470 22674 18522
rect 22726 18470 22738 18522
rect 22790 18470 22802 18522
rect 22854 18470 22866 18522
rect 22918 18470 27610 18522
rect 27662 18470 27674 18522
rect 27726 18470 27738 18522
rect 27790 18470 27802 18522
rect 27854 18470 27866 18522
rect 27918 18470 32610 18522
rect 32662 18470 32674 18522
rect 32726 18470 32738 18522
rect 32790 18470 32802 18522
rect 32854 18470 32866 18522
rect 32918 18470 37610 18522
rect 37662 18470 37674 18522
rect 37726 18470 37738 18522
rect 37790 18470 37802 18522
rect 37854 18470 37866 18522
rect 37918 18470 40848 18522
rect 1104 18448 40848 18470
rect 7466 18368 7472 18420
rect 7524 18408 7530 18420
rect 8110 18408 8116 18420
rect 7524 18380 8116 18408
rect 7524 18368 7530 18380
rect 8110 18368 8116 18380
rect 8168 18368 8174 18420
rect 29549 18411 29607 18417
rect 29549 18377 29561 18411
rect 29595 18408 29607 18411
rect 29638 18408 29644 18420
rect 29595 18380 29644 18408
rect 29595 18377 29607 18380
rect 29549 18371 29607 18377
rect 29638 18368 29644 18380
rect 29696 18408 29702 18420
rect 35618 18408 35624 18420
rect 29696 18380 35624 18408
rect 29696 18368 29702 18380
rect 35618 18368 35624 18380
rect 35676 18368 35682 18420
rect 25406 18232 25412 18284
rect 25464 18272 25470 18284
rect 29457 18275 29515 18281
rect 29457 18272 29469 18275
rect 25464 18244 29469 18272
rect 25464 18232 25470 18244
rect 29457 18241 29469 18244
rect 29503 18241 29515 18275
rect 29457 18235 29515 18241
rect 29546 18232 29552 18284
rect 29604 18272 29610 18284
rect 30009 18275 30067 18281
rect 30009 18272 30021 18275
rect 29604 18244 30021 18272
rect 29604 18232 29610 18244
rect 30009 18241 30021 18244
rect 30055 18272 30067 18275
rect 30098 18272 30104 18284
rect 30055 18244 30104 18272
rect 30055 18241 30067 18244
rect 30009 18235 30067 18241
rect 30098 18232 30104 18244
rect 30156 18232 30162 18284
rect 25682 18164 25688 18216
rect 25740 18204 25746 18216
rect 30285 18207 30343 18213
rect 30285 18204 30297 18207
rect 25740 18176 30297 18204
rect 25740 18164 25746 18176
rect 30285 18173 30297 18176
rect 30331 18173 30343 18207
rect 30285 18167 30343 18173
rect 33870 18028 33876 18080
rect 33928 18068 33934 18080
rect 37366 18068 37372 18080
rect 33928 18040 37372 18068
rect 33928 18028 33934 18040
rect 37366 18028 37372 18040
rect 37424 18028 37430 18080
rect 1104 17978 40848 18000
rect 1104 17926 1950 17978
rect 2002 17926 2014 17978
rect 2066 17926 2078 17978
rect 2130 17926 2142 17978
rect 2194 17926 2206 17978
rect 2258 17926 6950 17978
rect 7002 17926 7014 17978
rect 7066 17926 7078 17978
rect 7130 17926 7142 17978
rect 7194 17926 7206 17978
rect 7258 17926 11950 17978
rect 12002 17926 12014 17978
rect 12066 17926 12078 17978
rect 12130 17926 12142 17978
rect 12194 17926 12206 17978
rect 12258 17926 16950 17978
rect 17002 17926 17014 17978
rect 17066 17926 17078 17978
rect 17130 17926 17142 17978
rect 17194 17926 17206 17978
rect 17258 17926 21950 17978
rect 22002 17926 22014 17978
rect 22066 17926 22078 17978
rect 22130 17926 22142 17978
rect 22194 17926 22206 17978
rect 22258 17926 26950 17978
rect 27002 17926 27014 17978
rect 27066 17926 27078 17978
rect 27130 17926 27142 17978
rect 27194 17926 27206 17978
rect 27258 17926 31950 17978
rect 32002 17926 32014 17978
rect 32066 17926 32078 17978
rect 32130 17926 32142 17978
rect 32194 17926 32206 17978
rect 32258 17926 36950 17978
rect 37002 17926 37014 17978
rect 37066 17926 37078 17978
rect 37130 17926 37142 17978
rect 37194 17926 37206 17978
rect 37258 17926 40848 17978
rect 1104 17904 40848 17926
rect 34330 17824 34336 17876
rect 34388 17864 34394 17876
rect 35342 17864 35348 17876
rect 34388 17836 35348 17864
rect 34388 17824 34394 17836
rect 35342 17824 35348 17836
rect 35400 17824 35406 17876
rect 36722 17824 36728 17876
rect 36780 17864 36786 17876
rect 38657 17867 38715 17873
rect 38657 17864 38669 17867
rect 36780 17836 38669 17864
rect 36780 17824 36786 17836
rect 38657 17833 38669 17836
rect 38703 17833 38715 17867
rect 38657 17827 38715 17833
rect 24210 17688 24216 17740
rect 24268 17728 24274 17740
rect 39117 17731 39175 17737
rect 39117 17728 39129 17731
rect 24268 17700 39129 17728
rect 24268 17688 24274 17700
rect 39117 17697 39129 17700
rect 39163 17697 39175 17731
rect 39117 17691 39175 17697
rect 18874 17620 18880 17672
rect 18932 17660 18938 17672
rect 38841 17663 38899 17669
rect 38841 17660 38853 17663
rect 18932 17632 38853 17660
rect 18932 17620 18938 17632
rect 38841 17629 38853 17632
rect 38887 17629 38899 17663
rect 38841 17623 38899 17629
rect 38930 17620 38936 17672
rect 38988 17620 38994 17672
rect 39025 17663 39083 17669
rect 39025 17629 39037 17663
rect 39071 17629 39083 17663
rect 39025 17623 39083 17629
rect 35066 17552 35072 17604
rect 35124 17592 35130 17604
rect 39040 17592 39068 17623
rect 35124 17564 39068 17592
rect 35124 17552 35130 17564
rect 4522 17484 4528 17536
rect 4580 17524 4586 17536
rect 14550 17524 14556 17536
rect 4580 17496 14556 17524
rect 4580 17484 4586 17496
rect 14550 17484 14556 17496
rect 14608 17484 14614 17536
rect 1104 17434 40848 17456
rect 1104 17382 2610 17434
rect 2662 17382 2674 17434
rect 2726 17382 2738 17434
rect 2790 17382 2802 17434
rect 2854 17382 2866 17434
rect 2918 17382 7610 17434
rect 7662 17382 7674 17434
rect 7726 17382 7738 17434
rect 7790 17382 7802 17434
rect 7854 17382 7866 17434
rect 7918 17382 12610 17434
rect 12662 17382 12674 17434
rect 12726 17382 12738 17434
rect 12790 17382 12802 17434
rect 12854 17382 12866 17434
rect 12918 17382 17610 17434
rect 17662 17382 17674 17434
rect 17726 17382 17738 17434
rect 17790 17382 17802 17434
rect 17854 17382 17866 17434
rect 17918 17382 22610 17434
rect 22662 17382 22674 17434
rect 22726 17382 22738 17434
rect 22790 17382 22802 17434
rect 22854 17382 22866 17434
rect 22918 17382 27610 17434
rect 27662 17382 27674 17434
rect 27726 17382 27738 17434
rect 27790 17382 27802 17434
rect 27854 17382 27866 17434
rect 27918 17382 32610 17434
rect 32662 17382 32674 17434
rect 32726 17382 32738 17434
rect 32790 17382 32802 17434
rect 32854 17382 32866 17434
rect 32918 17382 37610 17434
rect 37662 17382 37674 17434
rect 37726 17382 37738 17434
rect 37790 17382 37802 17434
rect 37854 17382 37866 17434
rect 37918 17382 40848 17434
rect 1104 17360 40848 17382
rect 3050 17280 3056 17332
rect 3108 17320 3114 17332
rect 18138 17320 18144 17332
rect 3108 17292 18144 17320
rect 3108 17280 3114 17292
rect 18138 17280 18144 17292
rect 18196 17280 18202 17332
rect 7466 17212 7472 17264
rect 7524 17252 7530 17264
rect 30006 17252 30012 17264
rect 7524 17224 30012 17252
rect 7524 17212 7530 17224
rect 30006 17212 30012 17224
rect 30064 17212 30070 17264
rect 1104 16890 40848 16912
rect 1104 16838 1950 16890
rect 2002 16838 2014 16890
rect 2066 16838 2078 16890
rect 2130 16838 2142 16890
rect 2194 16838 2206 16890
rect 2258 16838 6950 16890
rect 7002 16838 7014 16890
rect 7066 16838 7078 16890
rect 7130 16838 7142 16890
rect 7194 16838 7206 16890
rect 7258 16838 11950 16890
rect 12002 16838 12014 16890
rect 12066 16838 12078 16890
rect 12130 16838 12142 16890
rect 12194 16838 12206 16890
rect 12258 16838 16950 16890
rect 17002 16838 17014 16890
rect 17066 16838 17078 16890
rect 17130 16838 17142 16890
rect 17194 16838 17206 16890
rect 17258 16838 21950 16890
rect 22002 16838 22014 16890
rect 22066 16838 22078 16890
rect 22130 16838 22142 16890
rect 22194 16838 22206 16890
rect 22258 16838 26950 16890
rect 27002 16838 27014 16890
rect 27066 16838 27078 16890
rect 27130 16838 27142 16890
rect 27194 16838 27206 16890
rect 27258 16838 31950 16890
rect 32002 16838 32014 16890
rect 32066 16838 32078 16890
rect 32130 16838 32142 16890
rect 32194 16838 32206 16890
rect 32258 16838 36950 16890
rect 37002 16838 37014 16890
rect 37066 16838 37078 16890
rect 37130 16838 37142 16890
rect 37194 16838 37206 16890
rect 37258 16838 40848 16890
rect 1104 16816 40848 16838
rect 22278 16736 22284 16788
rect 22336 16776 22342 16788
rect 22336 16748 25084 16776
rect 22336 16736 22342 16748
rect 22370 16708 22376 16720
rect 12406 16680 22376 16708
rect 6546 16600 6552 16652
rect 6604 16600 6610 16652
rect 7101 16643 7159 16649
rect 7101 16609 7113 16643
rect 7147 16640 7159 16643
rect 12406 16640 12434 16680
rect 22370 16668 22376 16680
rect 22428 16668 22434 16720
rect 7147 16612 12434 16640
rect 7147 16609 7159 16612
rect 7101 16603 7159 16609
rect 24486 16600 24492 16652
rect 24544 16600 24550 16652
rect 25056 16649 25084 16748
rect 25041 16643 25099 16649
rect 25041 16609 25053 16643
rect 25087 16640 25099 16643
rect 34606 16640 34612 16652
rect 25087 16612 34612 16640
rect 25087 16609 25099 16612
rect 25041 16603 25099 16609
rect 34606 16600 34612 16612
rect 34664 16600 34670 16652
rect 7009 16575 7067 16581
rect 7009 16541 7021 16575
rect 7055 16572 7067 16575
rect 7374 16572 7380 16584
rect 7055 16544 7380 16572
rect 7055 16541 7067 16544
rect 7009 16535 7067 16541
rect 7374 16532 7380 16544
rect 7432 16532 7438 16584
rect 24946 16532 24952 16584
rect 25004 16572 25010 16584
rect 25590 16572 25596 16584
rect 25004 16544 25596 16572
rect 25004 16532 25010 16544
rect 25590 16532 25596 16544
rect 25648 16532 25654 16584
rect 28442 16464 28448 16516
rect 28500 16504 28506 16516
rect 35250 16504 35256 16516
rect 28500 16476 35256 16504
rect 28500 16464 28506 16476
rect 35250 16464 35256 16476
rect 35308 16464 35314 16516
rect 1104 16346 40848 16368
rect 1104 16294 2610 16346
rect 2662 16294 2674 16346
rect 2726 16294 2738 16346
rect 2790 16294 2802 16346
rect 2854 16294 2866 16346
rect 2918 16294 7610 16346
rect 7662 16294 7674 16346
rect 7726 16294 7738 16346
rect 7790 16294 7802 16346
rect 7854 16294 7866 16346
rect 7918 16294 12610 16346
rect 12662 16294 12674 16346
rect 12726 16294 12738 16346
rect 12790 16294 12802 16346
rect 12854 16294 12866 16346
rect 12918 16294 17610 16346
rect 17662 16294 17674 16346
rect 17726 16294 17738 16346
rect 17790 16294 17802 16346
rect 17854 16294 17866 16346
rect 17918 16294 22610 16346
rect 22662 16294 22674 16346
rect 22726 16294 22738 16346
rect 22790 16294 22802 16346
rect 22854 16294 22866 16346
rect 22918 16294 27610 16346
rect 27662 16294 27674 16346
rect 27726 16294 27738 16346
rect 27790 16294 27802 16346
rect 27854 16294 27866 16346
rect 27918 16294 32610 16346
rect 32662 16294 32674 16346
rect 32726 16294 32738 16346
rect 32790 16294 32802 16346
rect 32854 16294 32866 16346
rect 32918 16294 37610 16346
rect 37662 16294 37674 16346
rect 37726 16294 37738 16346
rect 37790 16294 37802 16346
rect 37854 16294 37866 16346
rect 37918 16294 40848 16346
rect 1104 16272 40848 16294
rect 2409 16235 2467 16241
rect 2409 16201 2421 16235
rect 2455 16232 2467 16235
rect 3510 16232 3516 16244
rect 2455 16204 3516 16232
rect 2455 16201 2467 16204
rect 2409 16195 2467 16201
rect 3510 16192 3516 16204
rect 3568 16192 3574 16244
rect 1949 16099 2007 16105
rect 1949 16065 1961 16099
rect 1995 16096 2007 16099
rect 2314 16096 2320 16108
rect 1995 16068 2320 16096
rect 1995 16065 2007 16068
rect 1949 16059 2007 16065
rect 2314 16056 2320 16068
rect 2372 16056 2378 16108
rect 2468 16099 2526 16105
rect 2468 16065 2480 16099
rect 2514 16096 2526 16099
rect 6362 16096 6368 16108
rect 2514 16068 6368 16096
rect 2514 16065 2526 16068
rect 2468 16059 2526 16065
rect 6362 16056 6368 16068
rect 6420 16056 6426 16108
rect 9214 16056 9220 16108
rect 9272 16096 9278 16108
rect 9272 16068 12434 16096
rect 9272 16056 9278 16068
rect 2041 16031 2099 16037
rect 2041 15997 2053 16031
rect 2087 16028 2099 16031
rect 9398 16028 9404 16040
rect 2087 16000 9404 16028
rect 2087 15997 2099 16000
rect 2041 15991 2099 15997
rect 9398 15988 9404 16000
rect 9456 15988 9462 16040
rect 12406 16028 12434 16068
rect 24854 16028 24860 16040
rect 12406 16000 24860 16028
rect 24854 15988 24860 16000
rect 24912 15988 24918 16040
rect 6178 15920 6184 15972
rect 6236 15960 6242 15972
rect 31018 15960 31024 15972
rect 6236 15932 31024 15960
rect 6236 15920 6242 15932
rect 31018 15920 31024 15932
rect 31076 15920 31082 15972
rect 2314 15852 2320 15904
rect 2372 15892 2378 15904
rect 2593 15895 2651 15901
rect 2593 15892 2605 15895
rect 2372 15864 2605 15892
rect 2372 15852 2378 15864
rect 2593 15861 2605 15864
rect 2639 15861 2651 15895
rect 2593 15855 2651 15861
rect 11790 15852 11796 15904
rect 11848 15892 11854 15904
rect 39298 15892 39304 15904
rect 11848 15864 39304 15892
rect 11848 15852 11854 15864
rect 39298 15852 39304 15864
rect 39356 15852 39362 15904
rect 1104 15802 40848 15824
rect 1104 15750 1950 15802
rect 2002 15750 2014 15802
rect 2066 15750 2078 15802
rect 2130 15750 2142 15802
rect 2194 15750 2206 15802
rect 2258 15750 6950 15802
rect 7002 15750 7014 15802
rect 7066 15750 7078 15802
rect 7130 15750 7142 15802
rect 7194 15750 7206 15802
rect 7258 15750 11950 15802
rect 12002 15750 12014 15802
rect 12066 15750 12078 15802
rect 12130 15750 12142 15802
rect 12194 15750 12206 15802
rect 12258 15750 16950 15802
rect 17002 15750 17014 15802
rect 17066 15750 17078 15802
rect 17130 15750 17142 15802
rect 17194 15750 17206 15802
rect 17258 15750 21950 15802
rect 22002 15750 22014 15802
rect 22066 15750 22078 15802
rect 22130 15750 22142 15802
rect 22194 15750 22206 15802
rect 22258 15750 26950 15802
rect 27002 15750 27014 15802
rect 27066 15750 27078 15802
rect 27130 15750 27142 15802
rect 27194 15750 27206 15802
rect 27258 15750 31950 15802
rect 32002 15750 32014 15802
rect 32066 15750 32078 15802
rect 32130 15750 32142 15802
rect 32194 15750 32206 15802
rect 32258 15750 36950 15802
rect 37002 15750 37014 15802
rect 37066 15750 37078 15802
rect 37130 15750 37142 15802
rect 37194 15750 37206 15802
rect 37258 15750 40848 15802
rect 1104 15728 40848 15750
rect 12986 15648 12992 15700
rect 13044 15648 13050 15700
rect 13446 15648 13452 15700
rect 13504 15648 13510 15700
rect 13170 15444 13176 15496
rect 13228 15444 13234 15496
rect 34698 15444 34704 15496
rect 34756 15444 34762 15496
rect 38194 15444 38200 15496
rect 38252 15484 38258 15496
rect 38562 15484 38568 15496
rect 38252 15456 38568 15484
rect 38252 15444 38258 15456
rect 38562 15444 38568 15456
rect 38620 15444 38626 15496
rect 13078 15376 13084 15428
rect 13136 15416 13142 15428
rect 13262 15416 13268 15428
rect 13136 15388 13268 15416
rect 13136 15376 13142 15388
rect 13262 15376 13268 15388
rect 13320 15376 13326 15428
rect 35526 15376 35532 15428
rect 35584 15376 35590 15428
rect 38378 15308 38384 15360
rect 38436 15348 38442 15360
rect 38562 15348 38568 15360
rect 38436 15320 38568 15348
rect 38436 15308 38442 15320
rect 38562 15308 38568 15320
rect 38620 15308 38626 15360
rect 1104 15258 40848 15280
rect 1104 15206 2610 15258
rect 2662 15206 2674 15258
rect 2726 15206 2738 15258
rect 2790 15206 2802 15258
rect 2854 15206 2866 15258
rect 2918 15206 7610 15258
rect 7662 15206 7674 15258
rect 7726 15206 7738 15258
rect 7790 15206 7802 15258
rect 7854 15206 7866 15258
rect 7918 15206 12610 15258
rect 12662 15206 12674 15258
rect 12726 15206 12738 15258
rect 12790 15206 12802 15258
rect 12854 15206 12866 15258
rect 12918 15206 17610 15258
rect 17662 15206 17674 15258
rect 17726 15206 17738 15258
rect 17790 15206 17802 15258
rect 17854 15206 17866 15258
rect 17918 15206 22610 15258
rect 22662 15206 22674 15258
rect 22726 15206 22738 15258
rect 22790 15206 22802 15258
rect 22854 15206 22866 15258
rect 22918 15206 27610 15258
rect 27662 15206 27674 15258
rect 27726 15206 27738 15258
rect 27790 15206 27802 15258
rect 27854 15206 27866 15258
rect 27918 15206 32610 15258
rect 32662 15206 32674 15258
rect 32726 15206 32738 15258
rect 32790 15206 32802 15258
rect 32854 15206 32866 15258
rect 32918 15206 37610 15258
rect 37662 15206 37674 15258
rect 37726 15206 37738 15258
rect 37790 15206 37802 15258
rect 37854 15206 37866 15258
rect 37918 15206 40848 15258
rect 1104 15184 40848 15206
rect 17218 15144 17224 15156
rect 15304 15116 17224 15144
rect 14550 15036 14556 15088
rect 14608 15036 14614 15088
rect 15304 15017 15332 15116
rect 17218 15104 17224 15116
rect 17276 15104 17282 15156
rect 18414 15104 18420 15156
rect 18472 15144 18478 15156
rect 20070 15144 20076 15156
rect 18472 15116 20076 15144
rect 18472 15104 18478 15116
rect 20070 15104 20076 15116
rect 20128 15104 20134 15156
rect 21818 15104 21824 15156
rect 21876 15144 21882 15156
rect 21876 15116 26234 15144
rect 21876 15104 21882 15116
rect 16574 15076 16580 15088
rect 15396 15048 16580 15076
rect 15289 15011 15347 15017
rect 15289 14977 15301 15011
rect 15335 14977 15347 15011
rect 15289 14971 15347 14977
rect 15105 14943 15163 14949
rect 15105 14909 15117 14943
rect 15151 14940 15163 14943
rect 15396 14940 15424 15048
rect 16574 15036 16580 15048
rect 16632 15036 16638 15088
rect 15565 15011 15623 15017
rect 15565 14977 15577 15011
rect 15611 15004 15623 15011
rect 23566 15008 23572 15020
rect 15672 15004 23572 15008
rect 15611 14980 23572 15004
rect 15611 14977 15700 14980
rect 15565 14976 15700 14977
rect 15565 14971 15623 14976
rect 23566 14968 23572 14980
rect 23624 14968 23630 15020
rect 15151 14912 15424 14940
rect 15473 14943 15531 14949
rect 15151 14909 15163 14912
rect 15105 14903 15163 14909
rect 15473 14909 15485 14943
rect 15519 14909 15531 14943
rect 15473 14903 15531 14909
rect 15488 14872 15516 14903
rect 17218 14900 17224 14952
rect 17276 14940 17282 14952
rect 26206 14940 26234 15116
rect 31018 15036 31024 15088
rect 31076 15036 31082 15088
rect 31202 15036 31208 15088
rect 31260 15076 31266 15088
rect 31260 15048 34560 15076
rect 31260 15036 31266 15048
rect 31386 14968 31392 15020
rect 31444 14968 31450 15020
rect 33686 14968 33692 15020
rect 33744 14968 33750 15020
rect 34238 14968 34244 15020
rect 34296 14968 34302 15020
rect 34532 15017 34560 15048
rect 37366 15036 37372 15088
rect 37424 15076 37430 15088
rect 37829 15079 37887 15085
rect 37829 15076 37841 15079
rect 37424 15048 37841 15076
rect 37424 15036 37430 15048
rect 37829 15045 37841 15048
rect 37875 15045 37887 15079
rect 37829 15039 37887 15045
rect 38381 15079 38439 15085
rect 38381 15045 38393 15079
rect 38427 15076 38439 15079
rect 38654 15076 38660 15088
rect 38427 15048 38660 15076
rect 38427 15045 38439 15048
rect 38381 15039 38439 15045
rect 38654 15036 38660 15048
rect 38712 15036 38718 15088
rect 34517 15011 34575 15017
rect 34517 14977 34529 15011
rect 34563 14977 34575 15011
rect 34517 14971 34575 14977
rect 17276 14912 22094 14940
rect 26206 14912 31616 14940
rect 17276 14900 17282 14912
rect 22066 14872 22094 14912
rect 31478 14872 31484 14884
rect 15488 14844 19334 14872
rect 22066 14844 31484 14872
rect 19306 14804 19334 14844
rect 31478 14832 31484 14844
rect 31536 14832 31542 14884
rect 26602 14804 26608 14816
rect 19306 14776 26608 14804
rect 26602 14764 26608 14776
rect 26660 14764 26666 14816
rect 31588 14804 31616 14912
rect 34330 14900 34336 14952
rect 34388 14900 34394 14952
rect 31754 14832 31760 14884
rect 31812 14832 31818 14884
rect 34532 14872 34560 14971
rect 35342 14968 35348 15020
rect 35400 14968 35406 15020
rect 38286 14968 38292 15020
rect 38344 14968 38350 15020
rect 34974 14900 34980 14952
rect 35032 14900 35038 14952
rect 35250 14900 35256 14952
rect 35308 14900 35314 14952
rect 39022 14872 39028 14884
rect 34532 14844 39028 14872
rect 39022 14832 39028 14844
rect 39080 14832 39086 14884
rect 38194 14804 38200 14816
rect 31588 14776 38200 14804
rect 38194 14764 38200 14776
rect 38252 14804 38258 14816
rect 38565 14807 38623 14813
rect 38565 14804 38577 14807
rect 38252 14776 38577 14804
rect 38252 14764 38258 14776
rect 38565 14773 38577 14776
rect 38611 14773 38623 14807
rect 38565 14767 38623 14773
rect 1104 14714 40848 14736
rect 1104 14662 1950 14714
rect 2002 14662 2014 14714
rect 2066 14662 2078 14714
rect 2130 14662 2142 14714
rect 2194 14662 2206 14714
rect 2258 14662 6950 14714
rect 7002 14662 7014 14714
rect 7066 14662 7078 14714
rect 7130 14662 7142 14714
rect 7194 14662 7206 14714
rect 7258 14662 11950 14714
rect 12002 14662 12014 14714
rect 12066 14662 12078 14714
rect 12130 14662 12142 14714
rect 12194 14662 12206 14714
rect 12258 14662 16950 14714
rect 17002 14662 17014 14714
rect 17066 14662 17078 14714
rect 17130 14662 17142 14714
rect 17194 14662 17206 14714
rect 17258 14662 21950 14714
rect 22002 14662 22014 14714
rect 22066 14662 22078 14714
rect 22130 14662 22142 14714
rect 22194 14662 22206 14714
rect 22258 14662 26950 14714
rect 27002 14662 27014 14714
rect 27066 14662 27078 14714
rect 27130 14662 27142 14714
rect 27194 14662 27206 14714
rect 27258 14662 31950 14714
rect 32002 14662 32014 14714
rect 32066 14662 32078 14714
rect 32130 14662 32142 14714
rect 32194 14662 32206 14714
rect 32258 14662 36950 14714
rect 37002 14662 37014 14714
rect 37066 14662 37078 14714
rect 37130 14662 37142 14714
rect 37194 14662 37206 14714
rect 37258 14662 40848 14714
rect 1104 14640 40848 14662
rect 9122 14560 9128 14612
rect 9180 14600 9186 14612
rect 38657 14603 38715 14609
rect 38657 14600 38669 14603
rect 9180 14572 38669 14600
rect 9180 14560 9186 14572
rect 38657 14569 38669 14572
rect 38703 14569 38715 14603
rect 38657 14563 38715 14569
rect 23474 14492 23480 14544
rect 23532 14532 23538 14544
rect 29086 14532 29092 14544
rect 23532 14504 29092 14532
rect 23532 14492 23538 14504
rect 29086 14492 29092 14504
rect 29144 14492 29150 14544
rect 30098 14492 30104 14544
rect 30156 14532 30162 14544
rect 31481 14535 31539 14541
rect 31481 14532 31493 14535
rect 30156 14504 31493 14532
rect 30156 14492 30162 14504
rect 31481 14501 31493 14504
rect 31527 14501 31539 14535
rect 31481 14495 31539 14501
rect 31941 14535 31999 14541
rect 31941 14501 31953 14535
rect 31987 14532 31999 14535
rect 32306 14532 32312 14544
rect 31987 14504 32312 14532
rect 31987 14501 31999 14504
rect 31941 14495 31999 14501
rect 32306 14492 32312 14504
rect 32364 14492 32370 14544
rect 38672 14532 38700 14563
rect 38672 14504 38792 14532
rect 26510 14424 26516 14476
rect 26568 14464 26574 14476
rect 26568 14436 31708 14464
rect 26568 14424 26574 14436
rect 30742 14356 30748 14408
rect 30800 14396 30806 14408
rect 31113 14399 31171 14405
rect 31113 14396 31125 14399
rect 30800 14368 31125 14396
rect 30800 14356 30806 14368
rect 31113 14365 31125 14368
rect 31159 14365 31171 14399
rect 31113 14359 31171 14365
rect 31294 14356 31300 14408
rect 31352 14356 31358 14408
rect 31680 14405 31708 14436
rect 32398 14424 32404 14476
rect 32456 14464 32462 14476
rect 38764 14464 38792 14504
rect 39393 14467 39451 14473
rect 32456 14436 35894 14464
rect 38764 14436 39252 14464
rect 32456 14424 32462 14436
rect 31665 14399 31723 14405
rect 31665 14365 31677 14399
rect 31711 14365 31723 14399
rect 31665 14359 31723 14365
rect 32217 14399 32275 14405
rect 32217 14365 32229 14399
rect 32263 14365 32275 14399
rect 32217 14359 32275 14365
rect 32677 14399 32735 14405
rect 32677 14365 32689 14399
rect 32723 14396 32735 14399
rect 33410 14396 33416 14408
rect 32723 14368 33416 14396
rect 32723 14365 32735 14368
rect 32677 14359 32735 14365
rect 29822 14288 29828 14340
rect 29880 14328 29886 14340
rect 31021 14331 31079 14337
rect 31021 14328 31033 14331
rect 29880 14300 31033 14328
rect 29880 14288 29886 14300
rect 31021 14297 31033 14300
rect 31067 14297 31079 14331
rect 31021 14291 31079 14297
rect 31202 14288 31208 14340
rect 31260 14328 31266 14340
rect 32232 14328 32260 14359
rect 33410 14356 33416 14368
rect 33468 14356 33474 14408
rect 35866 14396 35894 14436
rect 39224 14405 39252 14436
rect 39393 14433 39405 14467
rect 39439 14433 39451 14467
rect 39393 14427 39451 14433
rect 39209 14399 39267 14405
rect 35866 14368 39160 14396
rect 39132 14328 39160 14368
rect 39209 14365 39221 14399
rect 39255 14365 39267 14399
rect 39209 14359 39267 14365
rect 39298 14356 39304 14408
rect 39356 14356 39362 14408
rect 39408 14328 39436 14427
rect 39482 14424 39488 14476
rect 39540 14424 39546 14476
rect 31260 14300 32260 14328
rect 37476 14300 39068 14328
rect 39132 14300 39436 14328
rect 31260 14288 31266 14300
rect 35710 14220 35716 14272
rect 35768 14260 35774 14272
rect 37476 14260 37504 14300
rect 39040 14269 39068 14300
rect 35768 14232 37504 14260
rect 39025 14263 39083 14269
rect 35768 14220 35774 14232
rect 39025 14229 39037 14263
rect 39071 14229 39083 14263
rect 39025 14223 39083 14229
rect 1104 14170 40848 14192
rect 1104 14118 2610 14170
rect 2662 14118 2674 14170
rect 2726 14118 2738 14170
rect 2790 14118 2802 14170
rect 2854 14118 2866 14170
rect 2918 14118 7610 14170
rect 7662 14118 7674 14170
rect 7726 14118 7738 14170
rect 7790 14118 7802 14170
rect 7854 14118 7866 14170
rect 7918 14118 12610 14170
rect 12662 14118 12674 14170
rect 12726 14118 12738 14170
rect 12790 14118 12802 14170
rect 12854 14118 12866 14170
rect 12918 14118 17610 14170
rect 17662 14118 17674 14170
rect 17726 14118 17738 14170
rect 17790 14118 17802 14170
rect 17854 14118 17866 14170
rect 17918 14118 22610 14170
rect 22662 14118 22674 14170
rect 22726 14118 22738 14170
rect 22790 14118 22802 14170
rect 22854 14118 22866 14170
rect 22918 14118 27610 14170
rect 27662 14118 27674 14170
rect 27726 14118 27738 14170
rect 27790 14118 27802 14170
rect 27854 14118 27866 14170
rect 27918 14118 32610 14170
rect 32662 14118 32674 14170
rect 32726 14118 32738 14170
rect 32790 14118 32802 14170
rect 32854 14118 32866 14170
rect 32918 14118 37610 14170
rect 37662 14118 37674 14170
rect 37726 14118 37738 14170
rect 37790 14118 37802 14170
rect 37854 14118 37866 14170
rect 37918 14118 40848 14170
rect 1104 14096 40848 14118
rect 38746 14016 38752 14068
rect 38804 14056 38810 14068
rect 39025 14059 39083 14065
rect 39025 14056 39037 14059
rect 38804 14028 39037 14056
rect 38804 14016 38810 14028
rect 39025 14025 39037 14028
rect 39071 14025 39083 14059
rect 39025 14019 39083 14025
rect 1394 13880 1400 13932
rect 1452 13880 1458 13932
rect 19150 13880 19156 13932
rect 19208 13920 19214 13932
rect 38013 13923 38071 13929
rect 38013 13920 38025 13923
rect 19208 13892 38025 13920
rect 19208 13880 19214 13892
rect 38013 13889 38025 13892
rect 38059 13889 38071 13923
rect 38013 13883 38071 13889
rect 38378 13880 38384 13932
rect 38436 13880 38442 13932
rect 38749 13923 38807 13929
rect 38749 13889 38761 13923
rect 38795 13920 38807 13923
rect 38838 13920 38844 13932
rect 38795 13892 38844 13920
rect 38795 13889 38807 13892
rect 38749 13883 38807 13889
rect 38838 13880 38844 13892
rect 38896 13880 38902 13932
rect 39942 13880 39948 13932
rect 40000 13920 40006 13932
rect 40313 13923 40371 13929
rect 40313 13920 40325 13923
rect 40000 13892 40325 13920
rect 40000 13880 40006 13892
rect 40313 13889 40325 13892
rect 40359 13889 40371 13923
rect 40313 13883 40371 13889
rect 3145 13855 3203 13861
rect 3145 13821 3157 13855
rect 3191 13852 3203 13855
rect 13538 13852 13544 13864
rect 3191 13824 13544 13852
rect 3191 13821 3203 13824
rect 3145 13815 3203 13821
rect 13538 13812 13544 13824
rect 13596 13812 13602 13864
rect 33410 13812 33416 13864
rect 33468 13852 33474 13864
rect 39669 13855 39727 13861
rect 39669 13852 39681 13855
rect 33468 13824 39681 13852
rect 33468 13812 33474 13824
rect 39669 13821 39681 13824
rect 39715 13821 39727 13855
rect 39669 13815 39727 13821
rect 1104 13626 40848 13648
rect 1104 13574 1950 13626
rect 2002 13574 2014 13626
rect 2066 13574 2078 13626
rect 2130 13574 2142 13626
rect 2194 13574 2206 13626
rect 2258 13574 6950 13626
rect 7002 13574 7014 13626
rect 7066 13574 7078 13626
rect 7130 13574 7142 13626
rect 7194 13574 7206 13626
rect 7258 13574 11950 13626
rect 12002 13574 12014 13626
rect 12066 13574 12078 13626
rect 12130 13574 12142 13626
rect 12194 13574 12206 13626
rect 12258 13574 16950 13626
rect 17002 13574 17014 13626
rect 17066 13574 17078 13626
rect 17130 13574 17142 13626
rect 17194 13574 17206 13626
rect 17258 13574 21950 13626
rect 22002 13574 22014 13626
rect 22066 13574 22078 13626
rect 22130 13574 22142 13626
rect 22194 13574 22206 13626
rect 22258 13574 26950 13626
rect 27002 13574 27014 13626
rect 27066 13574 27078 13626
rect 27130 13574 27142 13626
rect 27194 13574 27206 13626
rect 27258 13574 31950 13626
rect 32002 13574 32014 13626
rect 32066 13574 32078 13626
rect 32130 13574 32142 13626
rect 32194 13574 32206 13626
rect 32258 13574 36950 13626
rect 37002 13574 37014 13626
rect 37066 13574 37078 13626
rect 37130 13574 37142 13626
rect 37194 13574 37206 13626
rect 37258 13574 40848 13626
rect 1104 13552 40848 13574
rect 38746 13472 38752 13524
rect 38804 13512 38810 13524
rect 39577 13515 39635 13521
rect 39577 13512 39589 13515
rect 38804 13484 39589 13512
rect 38804 13472 38810 13484
rect 39577 13481 39589 13484
rect 39623 13481 39635 13515
rect 39577 13475 39635 13481
rect 34238 13336 34244 13388
rect 34296 13376 34302 13388
rect 34296 13348 39528 13376
rect 34296 13336 34302 13348
rect 39022 13268 39028 13320
rect 39080 13268 39086 13320
rect 39398 13311 39456 13317
rect 39398 13308 39410 13311
rect 39132 13280 39410 13308
rect 35526 13200 35532 13252
rect 35584 13240 35590 13252
rect 39132 13240 39160 13280
rect 39398 13277 39410 13280
rect 39444 13277 39456 13311
rect 39398 13271 39456 13277
rect 35584 13212 39160 13240
rect 39209 13243 39267 13249
rect 35584 13200 35590 13212
rect 39209 13209 39221 13243
rect 39255 13209 39267 13243
rect 39209 13203 39267 13209
rect 39301 13243 39359 13249
rect 39301 13209 39313 13243
rect 39347 13240 39359 13243
rect 39500 13240 39528 13348
rect 39347 13212 39528 13240
rect 39347 13209 39359 13212
rect 39301 13203 39359 13209
rect 7374 13132 7380 13184
rect 7432 13172 7438 13184
rect 21634 13172 21640 13184
rect 7432 13144 21640 13172
rect 7432 13132 7438 13144
rect 21634 13132 21640 13144
rect 21692 13132 21698 13184
rect 38562 13132 38568 13184
rect 38620 13172 38626 13184
rect 39224 13172 39252 13203
rect 38620 13144 39252 13172
rect 38620 13132 38626 13144
rect 1104 13082 40848 13104
rect 1104 13030 2610 13082
rect 2662 13030 2674 13082
rect 2726 13030 2738 13082
rect 2790 13030 2802 13082
rect 2854 13030 2866 13082
rect 2918 13030 7610 13082
rect 7662 13030 7674 13082
rect 7726 13030 7738 13082
rect 7790 13030 7802 13082
rect 7854 13030 7866 13082
rect 7918 13030 12610 13082
rect 12662 13030 12674 13082
rect 12726 13030 12738 13082
rect 12790 13030 12802 13082
rect 12854 13030 12866 13082
rect 12918 13030 17610 13082
rect 17662 13030 17674 13082
rect 17726 13030 17738 13082
rect 17790 13030 17802 13082
rect 17854 13030 17866 13082
rect 17918 13030 22610 13082
rect 22662 13030 22674 13082
rect 22726 13030 22738 13082
rect 22790 13030 22802 13082
rect 22854 13030 22866 13082
rect 22918 13030 27610 13082
rect 27662 13030 27674 13082
rect 27726 13030 27738 13082
rect 27790 13030 27802 13082
rect 27854 13030 27866 13082
rect 27918 13030 32610 13082
rect 32662 13030 32674 13082
rect 32726 13030 32738 13082
rect 32790 13030 32802 13082
rect 32854 13030 32866 13082
rect 32918 13030 37610 13082
rect 37662 13030 37674 13082
rect 37726 13030 37738 13082
rect 37790 13030 37802 13082
rect 37854 13030 37866 13082
rect 37918 13030 40848 13082
rect 1104 13008 40848 13030
rect 23290 12928 23296 12980
rect 23348 12928 23354 12980
rect 38746 12928 38752 12980
rect 38804 12968 38810 12980
rect 39025 12971 39083 12977
rect 39025 12968 39037 12971
rect 38804 12940 39037 12968
rect 38804 12928 38810 12940
rect 39025 12937 39037 12940
rect 39071 12937 39083 12971
rect 39025 12931 39083 12937
rect 21450 12792 21456 12844
rect 21508 12832 21514 12844
rect 23201 12835 23259 12841
rect 23201 12832 23213 12835
rect 21508 12804 23213 12832
rect 21508 12792 21514 12804
rect 23201 12801 23213 12804
rect 23247 12801 23259 12835
rect 23201 12795 23259 12801
rect 23216 12764 23244 12795
rect 23382 12792 23388 12844
rect 23440 12792 23446 12844
rect 30282 12764 30288 12776
rect 23216 12736 30288 12764
rect 30282 12724 30288 12736
rect 30340 12724 30346 12776
rect 1104 12538 40848 12560
rect 1104 12486 1950 12538
rect 2002 12486 2014 12538
rect 2066 12486 2078 12538
rect 2130 12486 2142 12538
rect 2194 12486 2206 12538
rect 2258 12486 6950 12538
rect 7002 12486 7014 12538
rect 7066 12486 7078 12538
rect 7130 12486 7142 12538
rect 7194 12486 7206 12538
rect 7258 12486 11950 12538
rect 12002 12486 12014 12538
rect 12066 12486 12078 12538
rect 12130 12486 12142 12538
rect 12194 12486 12206 12538
rect 12258 12486 16950 12538
rect 17002 12486 17014 12538
rect 17066 12486 17078 12538
rect 17130 12486 17142 12538
rect 17194 12486 17206 12538
rect 17258 12486 21950 12538
rect 22002 12486 22014 12538
rect 22066 12486 22078 12538
rect 22130 12486 22142 12538
rect 22194 12486 22206 12538
rect 22258 12486 26950 12538
rect 27002 12486 27014 12538
rect 27066 12486 27078 12538
rect 27130 12486 27142 12538
rect 27194 12486 27206 12538
rect 27258 12486 31950 12538
rect 32002 12486 32014 12538
rect 32066 12486 32078 12538
rect 32130 12486 32142 12538
rect 32194 12486 32206 12538
rect 32258 12486 36950 12538
rect 37002 12486 37014 12538
rect 37066 12486 37078 12538
rect 37130 12486 37142 12538
rect 37194 12486 37206 12538
rect 37258 12486 40848 12538
rect 1104 12464 40848 12486
rect 21542 12288 21548 12300
rect 16684 12260 21548 12288
rect 16482 12180 16488 12232
rect 16540 12180 16546 12232
rect 16684 12229 16712 12260
rect 21542 12248 21548 12260
rect 21600 12248 21606 12300
rect 16669 12223 16727 12229
rect 16669 12189 16681 12223
rect 16715 12189 16727 12223
rect 16669 12183 16727 12189
rect 16853 12223 16911 12229
rect 16853 12189 16865 12223
rect 16899 12220 16911 12223
rect 21358 12220 21364 12232
rect 16899 12192 21364 12220
rect 16899 12189 16911 12192
rect 16853 12183 16911 12189
rect 21358 12180 21364 12192
rect 21416 12180 21422 12232
rect 17313 12155 17371 12161
rect 17313 12121 17325 12155
rect 17359 12152 17371 12155
rect 31754 12152 31760 12164
rect 17359 12124 31760 12152
rect 17359 12121 17371 12124
rect 17313 12115 17371 12121
rect 31754 12112 31760 12124
rect 31812 12112 31818 12164
rect 1104 11994 40848 12016
rect 1104 11942 2610 11994
rect 2662 11942 2674 11994
rect 2726 11942 2738 11994
rect 2790 11942 2802 11994
rect 2854 11942 2866 11994
rect 2918 11942 7610 11994
rect 7662 11942 7674 11994
rect 7726 11942 7738 11994
rect 7790 11942 7802 11994
rect 7854 11942 7866 11994
rect 7918 11942 12610 11994
rect 12662 11942 12674 11994
rect 12726 11942 12738 11994
rect 12790 11942 12802 11994
rect 12854 11942 12866 11994
rect 12918 11942 17610 11994
rect 17662 11942 17674 11994
rect 17726 11942 17738 11994
rect 17790 11942 17802 11994
rect 17854 11942 17866 11994
rect 17918 11942 22610 11994
rect 22662 11942 22674 11994
rect 22726 11942 22738 11994
rect 22790 11942 22802 11994
rect 22854 11942 22866 11994
rect 22918 11942 27610 11994
rect 27662 11942 27674 11994
rect 27726 11942 27738 11994
rect 27790 11942 27802 11994
rect 27854 11942 27866 11994
rect 27918 11942 32610 11994
rect 32662 11942 32674 11994
rect 32726 11942 32738 11994
rect 32790 11942 32802 11994
rect 32854 11942 32866 11994
rect 32918 11942 37610 11994
rect 37662 11942 37674 11994
rect 37726 11942 37738 11994
rect 37790 11942 37802 11994
rect 37854 11942 37866 11994
rect 37918 11942 40848 11994
rect 1104 11920 40848 11942
rect 3142 11704 3148 11756
rect 3200 11744 3206 11756
rect 29638 11744 29644 11756
rect 3200 11716 29644 11744
rect 3200 11704 3206 11716
rect 29638 11704 29644 11716
rect 29696 11704 29702 11756
rect 1104 11450 40848 11472
rect 1104 11398 1950 11450
rect 2002 11398 2014 11450
rect 2066 11398 2078 11450
rect 2130 11398 2142 11450
rect 2194 11398 2206 11450
rect 2258 11398 6950 11450
rect 7002 11398 7014 11450
rect 7066 11398 7078 11450
rect 7130 11398 7142 11450
rect 7194 11398 7206 11450
rect 7258 11398 11950 11450
rect 12002 11398 12014 11450
rect 12066 11398 12078 11450
rect 12130 11398 12142 11450
rect 12194 11398 12206 11450
rect 12258 11398 16950 11450
rect 17002 11398 17014 11450
rect 17066 11398 17078 11450
rect 17130 11398 17142 11450
rect 17194 11398 17206 11450
rect 17258 11398 21950 11450
rect 22002 11398 22014 11450
rect 22066 11398 22078 11450
rect 22130 11398 22142 11450
rect 22194 11398 22206 11450
rect 22258 11398 26950 11450
rect 27002 11398 27014 11450
rect 27066 11398 27078 11450
rect 27130 11398 27142 11450
rect 27194 11398 27206 11450
rect 27258 11398 31950 11450
rect 32002 11398 32014 11450
rect 32066 11398 32078 11450
rect 32130 11398 32142 11450
rect 32194 11398 32206 11450
rect 32258 11398 36950 11450
rect 37002 11398 37014 11450
rect 37066 11398 37078 11450
rect 37130 11398 37142 11450
rect 37194 11398 37206 11450
rect 37258 11398 40848 11450
rect 1104 11376 40848 11398
rect 13262 11228 13268 11280
rect 13320 11268 13326 11280
rect 13320 11240 32628 11268
rect 13320 11228 13326 11240
rect 21082 11200 21088 11212
rect 14936 11172 21088 11200
rect 2406 11092 2412 11144
rect 2464 11092 2470 11144
rect 14936 11141 14964 11172
rect 21082 11160 21088 11172
rect 21140 11160 21146 11212
rect 23566 11160 23572 11212
rect 23624 11200 23630 11212
rect 23624 11172 26234 11200
rect 23624 11160 23630 11172
rect 14921 11135 14979 11141
rect 14921 11101 14933 11135
rect 14967 11101 14979 11135
rect 14921 11095 14979 11101
rect 15102 11092 15108 11144
rect 15160 11092 15166 11144
rect 15289 11135 15347 11141
rect 15289 11101 15301 11135
rect 15335 11132 15347 11135
rect 16574 11132 16580 11144
rect 15335 11104 16580 11132
rect 15335 11101 15347 11104
rect 15289 11095 15347 11101
rect 16574 11092 16580 11104
rect 16632 11092 16638 11144
rect 3421 11067 3479 11073
rect 3421 11033 3433 11067
rect 3467 11064 3479 11067
rect 6086 11064 6092 11076
rect 3467 11036 6092 11064
rect 3467 11033 3479 11036
rect 3421 11027 3479 11033
rect 6086 11024 6092 11036
rect 6144 11024 6150 11076
rect 15749 11067 15807 11073
rect 15749 11033 15761 11067
rect 15795 11064 15807 11067
rect 18414 11064 18420 11076
rect 15795 11036 18420 11064
rect 15795 11033 15807 11036
rect 15749 11027 15807 11033
rect 18414 11024 18420 11036
rect 18472 11024 18478 11076
rect 26206 11064 26234 11172
rect 32398 11092 32404 11144
rect 32456 11092 32462 11144
rect 32600 11141 32628 11240
rect 32585 11135 32643 11141
rect 32585 11101 32597 11135
rect 32631 11101 32643 11135
rect 32585 11095 32643 11101
rect 33594 11092 33600 11144
rect 33652 11092 33658 11144
rect 34606 11092 34612 11144
rect 34664 11132 34670 11144
rect 37461 11135 37519 11141
rect 37461 11132 37473 11135
rect 34664 11104 37473 11132
rect 34664 11092 34670 11104
rect 37461 11101 37473 11104
rect 37507 11101 37519 11135
rect 37461 11095 37519 11101
rect 36449 11067 36507 11073
rect 36449 11064 36461 11067
rect 26206 11036 36461 11064
rect 36449 11033 36461 11036
rect 36495 11033 36507 11067
rect 36449 11027 36507 11033
rect 21174 10956 21180 11008
rect 21232 10996 21238 11008
rect 28166 10996 28172 11008
rect 21232 10968 28172 10996
rect 21232 10956 21238 10968
rect 28166 10956 28172 10968
rect 28224 10956 28230 11008
rect 1104 10906 40848 10928
rect 1104 10854 2610 10906
rect 2662 10854 2674 10906
rect 2726 10854 2738 10906
rect 2790 10854 2802 10906
rect 2854 10854 2866 10906
rect 2918 10854 7610 10906
rect 7662 10854 7674 10906
rect 7726 10854 7738 10906
rect 7790 10854 7802 10906
rect 7854 10854 7866 10906
rect 7918 10854 12610 10906
rect 12662 10854 12674 10906
rect 12726 10854 12738 10906
rect 12790 10854 12802 10906
rect 12854 10854 12866 10906
rect 12918 10854 17610 10906
rect 17662 10854 17674 10906
rect 17726 10854 17738 10906
rect 17790 10854 17802 10906
rect 17854 10854 17866 10906
rect 17918 10854 22610 10906
rect 22662 10854 22674 10906
rect 22726 10854 22738 10906
rect 22790 10854 22802 10906
rect 22854 10854 22866 10906
rect 22918 10854 27610 10906
rect 27662 10854 27674 10906
rect 27726 10854 27738 10906
rect 27790 10854 27802 10906
rect 27854 10854 27866 10906
rect 27918 10854 32610 10906
rect 32662 10854 32674 10906
rect 32726 10854 32738 10906
rect 32790 10854 32802 10906
rect 32854 10854 32866 10906
rect 32918 10854 37610 10906
rect 37662 10854 37674 10906
rect 37726 10854 37738 10906
rect 37790 10854 37802 10906
rect 37854 10854 37866 10906
rect 37918 10854 40848 10906
rect 1104 10832 40848 10854
rect 2700 10696 6914 10724
rect 2700 10665 2728 10696
rect 2685 10659 2743 10665
rect 2685 10625 2697 10659
rect 2731 10625 2743 10659
rect 2685 10619 2743 10625
rect 3050 10616 3056 10668
rect 3108 10616 3114 10668
rect 6886 10656 6914 10696
rect 10962 10684 10968 10736
rect 11020 10724 11026 10736
rect 20438 10724 20444 10736
rect 11020 10696 20444 10724
rect 11020 10684 11026 10696
rect 20438 10684 20444 10696
rect 20496 10684 20502 10736
rect 18690 10656 18696 10668
rect 6886 10628 18696 10656
rect 18690 10616 18696 10628
rect 18748 10616 18754 10668
rect 3145 10591 3203 10597
rect 3145 10557 3157 10591
rect 3191 10588 3203 10591
rect 12342 10588 12348 10600
rect 3191 10560 12348 10588
rect 3191 10557 3203 10560
rect 3145 10551 3203 10557
rect 12342 10548 12348 10560
rect 12400 10548 12406 10600
rect 2501 10523 2559 10529
rect 2501 10489 2513 10523
rect 2547 10520 2559 10523
rect 8202 10520 8208 10532
rect 2547 10492 8208 10520
rect 2547 10489 2559 10492
rect 2501 10483 2559 10489
rect 8202 10480 8208 10492
rect 8260 10480 8266 10532
rect 17954 10480 17960 10532
rect 18012 10520 18018 10532
rect 36814 10520 36820 10532
rect 18012 10492 36820 10520
rect 18012 10480 18018 10492
rect 36814 10480 36820 10492
rect 36872 10480 36878 10532
rect 9306 10412 9312 10464
rect 9364 10452 9370 10464
rect 31202 10452 31208 10464
rect 9364 10424 31208 10452
rect 9364 10412 9370 10424
rect 31202 10412 31208 10424
rect 31260 10412 31266 10464
rect 1104 10362 40848 10384
rect 1104 10310 1950 10362
rect 2002 10310 2014 10362
rect 2066 10310 2078 10362
rect 2130 10310 2142 10362
rect 2194 10310 2206 10362
rect 2258 10310 6950 10362
rect 7002 10310 7014 10362
rect 7066 10310 7078 10362
rect 7130 10310 7142 10362
rect 7194 10310 7206 10362
rect 7258 10310 11950 10362
rect 12002 10310 12014 10362
rect 12066 10310 12078 10362
rect 12130 10310 12142 10362
rect 12194 10310 12206 10362
rect 12258 10310 16950 10362
rect 17002 10310 17014 10362
rect 17066 10310 17078 10362
rect 17130 10310 17142 10362
rect 17194 10310 17206 10362
rect 17258 10310 21950 10362
rect 22002 10310 22014 10362
rect 22066 10310 22078 10362
rect 22130 10310 22142 10362
rect 22194 10310 22206 10362
rect 22258 10310 26950 10362
rect 27002 10310 27014 10362
rect 27066 10310 27078 10362
rect 27130 10310 27142 10362
rect 27194 10310 27206 10362
rect 27258 10310 31950 10362
rect 32002 10310 32014 10362
rect 32066 10310 32078 10362
rect 32130 10310 32142 10362
rect 32194 10310 32206 10362
rect 32258 10310 36950 10362
rect 37002 10310 37014 10362
rect 37066 10310 37078 10362
rect 37130 10310 37142 10362
rect 37194 10310 37206 10362
rect 37258 10310 40848 10362
rect 1104 10288 40848 10310
rect 1104 9818 40848 9840
rect 1104 9766 2610 9818
rect 2662 9766 2674 9818
rect 2726 9766 2738 9818
rect 2790 9766 2802 9818
rect 2854 9766 2866 9818
rect 2918 9766 7610 9818
rect 7662 9766 7674 9818
rect 7726 9766 7738 9818
rect 7790 9766 7802 9818
rect 7854 9766 7866 9818
rect 7918 9766 12610 9818
rect 12662 9766 12674 9818
rect 12726 9766 12738 9818
rect 12790 9766 12802 9818
rect 12854 9766 12866 9818
rect 12918 9766 17610 9818
rect 17662 9766 17674 9818
rect 17726 9766 17738 9818
rect 17790 9766 17802 9818
rect 17854 9766 17866 9818
rect 17918 9766 22610 9818
rect 22662 9766 22674 9818
rect 22726 9766 22738 9818
rect 22790 9766 22802 9818
rect 22854 9766 22866 9818
rect 22918 9766 27610 9818
rect 27662 9766 27674 9818
rect 27726 9766 27738 9818
rect 27790 9766 27802 9818
rect 27854 9766 27866 9818
rect 27918 9766 32610 9818
rect 32662 9766 32674 9818
rect 32726 9766 32738 9818
rect 32790 9766 32802 9818
rect 32854 9766 32866 9818
rect 32918 9766 37610 9818
rect 37662 9766 37674 9818
rect 37726 9766 37738 9818
rect 37790 9766 37802 9818
rect 37854 9766 37866 9818
rect 37918 9766 40848 9818
rect 1104 9744 40848 9766
rect 14108 9676 14320 9704
rect 12986 9596 12992 9648
rect 13044 9636 13050 9648
rect 14108 9636 14136 9676
rect 13044 9608 14136 9636
rect 13044 9596 13050 9608
rect 14182 9596 14188 9648
rect 14240 9596 14246 9648
rect 13630 9528 13636 9580
rect 13688 9528 13694 9580
rect 13814 9528 13820 9580
rect 13872 9528 13878 9580
rect 14292 9577 14320 9676
rect 16669 9639 16727 9645
rect 16669 9605 16681 9639
rect 16715 9605 16727 9639
rect 16669 9599 16727 9605
rect 14001 9571 14059 9577
rect 14001 9537 14013 9571
rect 14047 9568 14059 9571
rect 14277 9571 14335 9577
rect 14047 9540 14228 9568
rect 14047 9537 14059 9540
rect 14001 9531 14059 9537
rect 2498 9460 2504 9512
rect 2556 9500 2562 9512
rect 14200 9500 14228 9540
rect 14277 9537 14289 9571
rect 14323 9568 14335 9571
rect 14323 9540 16160 9568
rect 14323 9537 14335 9540
rect 14277 9531 14335 9537
rect 15654 9500 15660 9512
rect 2556 9472 14044 9500
rect 14200 9472 15660 9500
rect 2556 9460 2562 9472
rect 14016 9432 14044 9472
rect 15654 9460 15660 9472
rect 15712 9500 15718 9512
rect 16022 9500 16028 9512
rect 15712 9472 16028 9500
rect 15712 9460 15718 9472
rect 16022 9460 16028 9472
rect 16080 9460 16086 9512
rect 16132 9500 16160 9540
rect 16574 9528 16580 9580
rect 16632 9568 16638 9580
rect 16684 9568 16712 9599
rect 16850 9596 16856 9648
rect 16908 9596 16914 9648
rect 32398 9636 32404 9648
rect 16960 9608 32404 9636
rect 16960 9568 16988 9608
rect 32398 9596 32404 9608
rect 32456 9596 32462 9648
rect 16632 9540 16988 9568
rect 17129 9571 17187 9577
rect 16632 9528 16638 9540
rect 17129 9537 17141 9571
rect 17175 9568 17187 9571
rect 17954 9568 17960 9580
rect 17175 9540 17960 9568
rect 17175 9537 17187 9540
rect 17129 9531 17187 9537
rect 17954 9528 17960 9540
rect 18012 9528 18018 9580
rect 23474 9500 23480 9512
rect 16132 9472 23480 9500
rect 23474 9460 23480 9472
rect 23532 9460 23538 9512
rect 17402 9432 17408 9444
rect 14016 9404 17408 9432
rect 17402 9392 17408 9404
rect 17460 9392 17466 9444
rect 16666 9324 16672 9376
rect 16724 9364 16730 9376
rect 16853 9367 16911 9373
rect 16853 9364 16865 9367
rect 16724 9336 16865 9364
rect 16724 9324 16730 9336
rect 16853 9333 16865 9336
rect 16899 9333 16911 9367
rect 16853 9327 16911 9333
rect 1104 9274 40848 9296
rect 1104 9222 1950 9274
rect 2002 9222 2014 9274
rect 2066 9222 2078 9274
rect 2130 9222 2142 9274
rect 2194 9222 2206 9274
rect 2258 9222 6950 9274
rect 7002 9222 7014 9274
rect 7066 9222 7078 9274
rect 7130 9222 7142 9274
rect 7194 9222 7206 9274
rect 7258 9222 11950 9274
rect 12002 9222 12014 9274
rect 12066 9222 12078 9274
rect 12130 9222 12142 9274
rect 12194 9222 12206 9274
rect 12258 9222 16950 9274
rect 17002 9222 17014 9274
rect 17066 9222 17078 9274
rect 17130 9222 17142 9274
rect 17194 9222 17206 9274
rect 17258 9222 21950 9274
rect 22002 9222 22014 9274
rect 22066 9222 22078 9274
rect 22130 9222 22142 9274
rect 22194 9222 22206 9274
rect 22258 9222 26950 9274
rect 27002 9222 27014 9274
rect 27066 9222 27078 9274
rect 27130 9222 27142 9274
rect 27194 9222 27206 9274
rect 27258 9222 31950 9274
rect 32002 9222 32014 9274
rect 32066 9222 32078 9274
rect 32130 9222 32142 9274
rect 32194 9222 32206 9274
rect 32258 9222 36950 9274
rect 37002 9222 37014 9274
rect 37066 9222 37078 9274
rect 37130 9222 37142 9274
rect 37194 9222 37206 9274
rect 37258 9222 40848 9274
rect 1104 9200 40848 9222
rect 35158 9120 35164 9172
rect 35216 9120 35222 9172
rect 3602 9092 3608 9104
rect 2332 9064 3608 9092
rect 1854 8984 1860 9036
rect 1912 8984 1918 9036
rect 2332 9033 2360 9064
rect 3602 9052 3608 9064
rect 3660 9052 3666 9104
rect 8202 9052 8208 9104
rect 8260 9092 8266 9104
rect 19150 9092 19156 9104
rect 8260 9064 19156 9092
rect 8260 9052 8266 9064
rect 19150 9052 19156 9064
rect 19208 9052 19214 9104
rect 23382 9052 23388 9104
rect 23440 9092 23446 9104
rect 34793 9095 34851 9101
rect 34793 9092 34805 9095
rect 23440 9064 34805 9092
rect 23440 9052 23446 9064
rect 34793 9061 34805 9064
rect 34839 9061 34851 9095
rect 34793 9055 34851 9061
rect 2317 9027 2375 9033
rect 2317 8993 2329 9027
rect 2363 8993 2375 9027
rect 4890 9024 4896 9036
rect 2317 8987 2375 8993
rect 2608 8996 4896 9024
rect 2225 8959 2283 8965
rect 2225 8925 2237 8959
rect 2271 8956 2283 8959
rect 2498 8956 2504 8968
rect 2271 8928 2504 8956
rect 2271 8925 2283 8928
rect 2225 8919 2283 8925
rect 2498 8916 2504 8928
rect 2556 8916 2562 8968
rect 2608 8965 2636 8996
rect 4890 8984 4896 8996
rect 4948 8984 4954 9036
rect 30282 8984 30288 9036
rect 30340 9024 30346 9036
rect 34701 9027 34759 9033
rect 34701 9024 34713 9027
rect 30340 8996 34713 9024
rect 30340 8984 30346 8996
rect 34701 8993 34713 8996
rect 34747 8993 34759 9027
rect 34701 8987 34759 8993
rect 2593 8959 2651 8965
rect 2593 8925 2605 8959
rect 2639 8925 2651 8959
rect 2593 8919 2651 8925
rect 2777 8959 2835 8965
rect 2777 8925 2789 8959
rect 2823 8956 2835 8959
rect 2823 8928 6914 8956
rect 2823 8925 2835 8928
rect 2777 8919 2835 8925
rect 6886 8888 6914 8928
rect 26694 8916 26700 8968
rect 26752 8956 26758 8968
rect 27065 8959 27123 8965
rect 27065 8956 27077 8959
rect 26752 8928 27077 8956
rect 26752 8916 26758 8928
rect 27065 8925 27077 8928
rect 27111 8925 27123 8959
rect 27065 8919 27123 8925
rect 27338 8916 27344 8968
rect 27396 8956 27402 8968
rect 27522 8956 27528 8968
rect 27396 8928 27528 8956
rect 27396 8916 27402 8928
rect 27522 8916 27528 8928
rect 27580 8916 27586 8968
rect 34977 8959 35035 8965
rect 34977 8925 34989 8959
rect 35023 8956 35035 8959
rect 35066 8956 35072 8968
rect 35023 8928 35072 8956
rect 35023 8925 35035 8928
rect 34977 8919 35035 8925
rect 35066 8916 35072 8928
rect 35124 8916 35130 8968
rect 26424 8900 26476 8906
rect 16574 8888 16580 8900
rect 6886 8860 16580 8888
rect 16574 8848 16580 8860
rect 16632 8848 16638 8900
rect 20254 8848 20260 8900
rect 20312 8888 20318 8900
rect 20312 8860 26424 8888
rect 20312 8848 20318 8860
rect 26424 8842 26476 8848
rect 1104 8730 40848 8752
rect 1104 8678 2610 8730
rect 2662 8678 2674 8730
rect 2726 8678 2738 8730
rect 2790 8678 2802 8730
rect 2854 8678 2866 8730
rect 2918 8678 7610 8730
rect 7662 8678 7674 8730
rect 7726 8678 7738 8730
rect 7790 8678 7802 8730
rect 7854 8678 7866 8730
rect 7918 8678 12610 8730
rect 12662 8678 12674 8730
rect 12726 8678 12738 8730
rect 12790 8678 12802 8730
rect 12854 8678 12866 8730
rect 12918 8678 17610 8730
rect 17662 8678 17674 8730
rect 17726 8678 17738 8730
rect 17790 8678 17802 8730
rect 17854 8678 17866 8730
rect 17918 8678 22610 8730
rect 22662 8678 22674 8730
rect 22726 8678 22738 8730
rect 22790 8678 22802 8730
rect 22854 8678 22866 8730
rect 22918 8678 27610 8730
rect 27662 8678 27674 8730
rect 27726 8678 27738 8730
rect 27790 8678 27802 8730
rect 27854 8678 27866 8730
rect 27918 8678 32610 8730
rect 32662 8678 32674 8730
rect 32726 8678 32738 8730
rect 32790 8678 32802 8730
rect 32854 8678 32866 8730
rect 32918 8678 37610 8730
rect 37662 8678 37674 8730
rect 37726 8678 37738 8730
rect 37790 8678 37802 8730
rect 37854 8678 37866 8730
rect 37918 8678 40848 8730
rect 1104 8656 40848 8678
rect 16206 8304 16212 8356
rect 16264 8344 16270 8356
rect 16666 8344 16672 8356
rect 16264 8316 16672 8344
rect 16264 8304 16270 8316
rect 16666 8304 16672 8316
rect 16724 8304 16730 8356
rect 34606 8304 34612 8356
rect 34664 8344 34670 8356
rect 36262 8344 36268 8356
rect 34664 8316 36268 8344
rect 34664 8304 34670 8316
rect 36262 8304 36268 8316
rect 36320 8304 36326 8356
rect 1104 8186 40848 8208
rect 1104 8134 1950 8186
rect 2002 8134 2014 8186
rect 2066 8134 2078 8186
rect 2130 8134 2142 8186
rect 2194 8134 2206 8186
rect 2258 8134 6950 8186
rect 7002 8134 7014 8186
rect 7066 8134 7078 8186
rect 7130 8134 7142 8186
rect 7194 8134 7206 8186
rect 7258 8134 11950 8186
rect 12002 8134 12014 8186
rect 12066 8134 12078 8186
rect 12130 8134 12142 8186
rect 12194 8134 12206 8186
rect 12258 8134 16950 8186
rect 17002 8134 17014 8186
rect 17066 8134 17078 8186
rect 17130 8134 17142 8186
rect 17194 8134 17206 8186
rect 17258 8134 21950 8186
rect 22002 8134 22014 8186
rect 22066 8134 22078 8186
rect 22130 8134 22142 8186
rect 22194 8134 22206 8186
rect 22258 8134 26950 8186
rect 27002 8134 27014 8186
rect 27066 8134 27078 8186
rect 27130 8134 27142 8186
rect 27194 8134 27206 8186
rect 27258 8134 31950 8186
rect 32002 8134 32014 8186
rect 32066 8134 32078 8186
rect 32130 8134 32142 8186
rect 32194 8134 32206 8186
rect 32258 8134 36950 8186
rect 37002 8134 37014 8186
rect 37066 8134 37078 8186
rect 37130 8134 37142 8186
rect 37194 8134 37206 8186
rect 37258 8134 40848 8186
rect 1104 8112 40848 8134
rect 26786 8032 26792 8084
rect 26844 8072 26850 8084
rect 27157 8075 27215 8081
rect 27157 8072 27169 8075
rect 26844 8044 27169 8072
rect 26844 8032 26850 8044
rect 27157 8041 27169 8044
rect 27203 8041 27215 8075
rect 27157 8035 27215 8041
rect 14642 7964 14648 8016
rect 14700 8004 14706 8016
rect 14700 7976 16574 8004
rect 14700 7964 14706 7976
rect 16390 7936 16396 7948
rect 15856 7908 16396 7936
rect 15654 7828 15660 7880
rect 15712 7828 15718 7880
rect 15856 7877 15884 7908
rect 16390 7896 16396 7908
rect 16448 7896 16454 7948
rect 15841 7871 15899 7877
rect 15841 7837 15853 7871
rect 15887 7837 15899 7871
rect 15841 7831 15899 7837
rect 16025 7871 16083 7877
rect 16025 7837 16037 7871
rect 16071 7837 16083 7871
rect 16546 7868 16574 7976
rect 30926 7964 30932 8016
rect 30984 8004 30990 8016
rect 37737 8007 37795 8013
rect 37737 8004 37749 8007
rect 30984 7976 37749 8004
rect 30984 7964 30990 7976
rect 37737 7973 37749 7976
rect 37783 7973 37795 8007
rect 37737 7967 37795 7973
rect 22462 7896 22468 7948
rect 22520 7936 22526 7948
rect 22520 7908 27844 7936
rect 22520 7896 22526 7908
rect 27709 7871 27767 7877
rect 27709 7868 27721 7871
rect 16546 7840 27721 7868
rect 16025 7831 16083 7837
rect 27709 7837 27721 7840
rect 27755 7837 27767 7871
rect 27816 7868 27844 7908
rect 36538 7896 36544 7948
rect 36596 7936 36602 7948
rect 37461 7939 37519 7945
rect 37461 7936 37473 7939
rect 36596 7908 37473 7936
rect 36596 7896 36602 7908
rect 37461 7905 37473 7908
rect 37507 7905 37519 7939
rect 37461 7899 37519 7905
rect 28077 7871 28135 7877
rect 28077 7868 28089 7871
rect 27816 7840 28089 7868
rect 27709 7831 27767 7837
rect 28077 7837 28089 7840
rect 28123 7837 28135 7871
rect 28077 7831 28135 7837
rect 13630 7760 13636 7812
rect 13688 7800 13694 7812
rect 16040 7800 16068 7831
rect 13688 7772 16068 7800
rect 16485 7803 16543 7809
rect 13688 7760 13694 7772
rect 16485 7769 16497 7803
rect 16531 7800 16543 7803
rect 22370 7800 22376 7812
rect 16531 7772 22376 7800
rect 16531 7769 16543 7772
rect 16485 7763 16543 7769
rect 22370 7760 22376 7772
rect 22428 7760 22434 7812
rect 24854 7692 24860 7744
rect 24912 7732 24918 7744
rect 37921 7735 37979 7741
rect 37921 7732 37933 7735
rect 24912 7704 37933 7732
rect 24912 7692 24918 7704
rect 37921 7701 37933 7704
rect 37967 7701 37979 7735
rect 37921 7695 37979 7701
rect 1104 7642 40848 7664
rect 1104 7590 2610 7642
rect 2662 7590 2674 7642
rect 2726 7590 2738 7642
rect 2790 7590 2802 7642
rect 2854 7590 2866 7642
rect 2918 7590 7610 7642
rect 7662 7590 7674 7642
rect 7726 7590 7738 7642
rect 7790 7590 7802 7642
rect 7854 7590 7866 7642
rect 7918 7590 12610 7642
rect 12662 7590 12674 7642
rect 12726 7590 12738 7642
rect 12790 7590 12802 7642
rect 12854 7590 12866 7642
rect 12918 7590 17610 7642
rect 17662 7590 17674 7642
rect 17726 7590 17738 7642
rect 17790 7590 17802 7642
rect 17854 7590 17866 7642
rect 17918 7590 22610 7642
rect 22662 7590 22674 7642
rect 22726 7590 22738 7642
rect 22790 7590 22802 7642
rect 22854 7590 22866 7642
rect 22918 7590 27610 7642
rect 27662 7590 27674 7642
rect 27726 7590 27738 7642
rect 27790 7590 27802 7642
rect 27854 7590 27866 7642
rect 27918 7590 32610 7642
rect 32662 7590 32674 7642
rect 32726 7590 32738 7642
rect 32790 7590 32802 7642
rect 32854 7590 32866 7642
rect 32918 7590 37610 7642
rect 37662 7590 37674 7642
rect 37726 7590 37738 7642
rect 37790 7590 37802 7642
rect 37854 7590 37866 7642
rect 37918 7590 40848 7642
rect 1104 7568 40848 7590
rect 8938 7488 8944 7540
rect 8996 7528 9002 7540
rect 8996 7500 21036 7528
rect 8996 7488 9002 7500
rect 18248 7432 20300 7460
rect 15746 7352 15752 7404
rect 15804 7392 15810 7404
rect 18248 7392 18276 7432
rect 15804 7364 18276 7392
rect 15804 7352 15810 7364
rect 19794 7352 19800 7404
rect 19852 7392 19858 7404
rect 20070 7392 20076 7404
rect 19852 7364 20076 7392
rect 19852 7352 19858 7364
rect 20070 7352 20076 7364
rect 20128 7352 20134 7404
rect 20272 7401 20300 7432
rect 21008 7401 21036 7500
rect 20257 7395 20315 7401
rect 20257 7361 20269 7395
rect 20303 7361 20315 7395
rect 20717 7395 20775 7401
rect 20717 7392 20729 7395
rect 20257 7355 20315 7361
rect 20548 7364 20729 7392
rect 6086 7284 6092 7336
rect 6144 7324 6150 7336
rect 6144 7296 6914 7324
rect 6144 7284 6150 7296
rect 6886 7256 6914 7296
rect 19886 7284 19892 7336
rect 19944 7284 19950 7336
rect 20548 7324 20576 7364
rect 20717 7361 20729 7364
rect 20763 7361 20775 7395
rect 20717 7355 20775 7361
rect 20993 7395 21051 7401
rect 20993 7361 21005 7395
rect 21039 7361 21051 7395
rect 20993 7355 21051 7361
rect 24946 7324 24952 7336
rect 20548 7296 24952 7324
rect 20548 7256 20576 7296
rect 24946 7284 24952 7296
rect 25004 7284 25010 7336
rect 6886 7228 20576 7256
rect 1104 7098 40848 7120
rect 1104 7046 1950 7098
rect 2002 7046 2014 7098
rect 2066 7046 2078 7098
rect 2130 7046 2142 7098
rect 2194 7046 2206 7098
rect 2258 7046 6950 7098
rect 7002 7046 7014 7098
rect 7066 7046 7078 7098
rect 7130 7046 7142 7098
rect 7194 7046 7206 7098
rect 7258 7046 11950 7098
rect 12002 7046 12014 7098
rect 12066 7046 12078 7098
rect 12130 7046 12142 7098
rect 12194 7046 12206 7098
rect 12258 7046 16950 7098
rect 17002 7046 17014 7098
rect 17066 7046 17078 7098
rect 17130 7046 17142 7098
rect 17194 7046 17206 7098
rect 17258 7046 21950 7098
rect 22002 7046 22014 7098
rect 22066 7046 22078 7098
rect 22130 7046 22142 7098
rect 22194 7046 22206 7098
rect 22258 7046 26950 7098
rect 27002 7046 27014 7098
rect 27066 7046 27078 7098
rect 27130 7046 27142 7098
rect 27194 7046 27206 7098
rect 27258 7046 31950 7098
rect 32002 7046 32014 7098
rect 32066 7046 32078 7098
rect 32130 7046 32142 7098
rect 32194 7046 32206 7098
rect 32258 7046 36950 7098
rect 37002 7046 37014 7098
rect 37066 7046 37078 7098
rect 37130 7046 37142 7098
rect 37194 7046 37206 7098
rect 37258 7046 40848 7098
rect 1104 7024 40848 7046
rect 34514 6808 34520 6860
rect 34572 6848 34578 6860
rect 34572 6820 35572 6848
rect 34572 6808 34578 6820
rect 35544 6792 35572 6820
rect 6822 6740 6828 6792
rect 6880 6780 6886 6792
rect 34885 6783 34943 6789
rect 34885 6780 34897 6783
rect 6880 6752 34897 6780
rect 6880 6740 6886 6752
rect 34885 6749 34897 6752
rect 34931 6749 34943 6783
rect 34885 6743 34943 6749
rect 16942 6672 16948 6724
rect 17000 6712 17006 6724
rect 21726 6712 21732 6724
rect 17000 6684 21732 6712
rect 17000 6672 17006 6684
rect 21726 6672 21732 6684
rect 21784 6672 21790 6724
rect 29638 6672 29644 6724
rect 29696 6712 29702 6724
rect 29696 6684 34652 6712
rect 29696 6672 29702 6684
rect 6178 6604 6184 6656
rect 6236 6644 6242 6656
rect 30190 6644 30196 6656
rect 6236 6616 30196 6644
rect 6236 6604 6242 6616
rect 30190 6604 30196 6616
rect 30248 6604 30254 6656
rect 34624 6644 34652 6684
rect 34698 6672 34704 6724
rect 34756 6672 34762 6724
rect 34900 6712 34928 6743
rect 35526 6740 35532 6792
rect 35584 6740 35590 6792
rect 35618 6740 35624 6792
rect 35676 6740 35682 6792
rect 37274 6712 37280 6724
rect 34900 6684 37280 6712
rect 37274 6672 37280 6684
rect 37332 6672 37338 6724
rect 35618 6644 35624 6656
rect 34624 6616 35624 6644
rect 35618 6604 35624 6616
rect 35676 6604 35682 6656
rect 1104 6554 40848 6576
rect 1104 6502 2610 6554
rect 2662 6502 2674 6554
rect 2726 6502 2738 6554
rect 2790 6502 2802 6554
rect 2854 6502 2866 6554
rect 2918 6502 7610 6554
rect 7662 6502 7674 6554
rect 7726 6502 7738 6554
rect 7790 6502 7802 6554
rect 7854 6502 7866 6554
rect 7918 6502 12610 6554
rect 12662 6502 12674 6554
rect 12726 6502 12738 6554
rect 12790 6502 12802 6554
rect 12854 6502 12866 6554
rect 12918 6502 17610 6554
rect 17662 6502 17674 6554
rect 17726 6502 17738 6554
rect 17790 6502 17802 6554
rect 17854 6502 17866 6554
rect 17918 6502 22610 6554
rect 22662 6502 22674 6554
rect 22726 6502 22738 6554
rect 22790 6502 22802 6554
rect 22854 6502 22866 6554
rect 22918 6502 27610 6554
rect 27662 6502 27674 6554
rect 27726 6502 27738 6554
rect 27790 6502 27802 6554
rect 27854 6502 27866 6554
rect 27918 6502 32610 6554
rect 32662 6502 32674 6554
rect 32726 6502 32738 6554
rect 32790 6502 32802 6554
rect 32854 6502 32866 6554
rect 32918 6502 37610 6554
rect 37662 6502 37674 6554
rect 37726 6502 37738 6554
rect 37790 6502 37802 6554
rect 37854 6502 37866 6554
rect 37918 6502 40848 6554
rect 1104 6480 40848 6502
rect 5718 6400 5724 6452
rect 5776 6400 5782 6452
rect 37366 6440 37372 6452
rect 5828 6412 37372 6440
rect 1394 6332 1400 6384
rect 1452 6372 1458 6384
rect 5828 6372 5856 6412
rect 37366 6400 37372 6412
rect 37424 6400 37430 6452
rect 17405 6375 17463 6381
rect 1452 6344 5856 6372
rect 5920 6344 6914 6372
rect 1452 6332 1458 6344
rect 5920 6313 5948 6344
rect 5905 6307 5963 6313
rect 5905 6273 5917 6307
rect 5951 6273 5963 6307
rect 5905 6267 5963 6273
rect 6178 6264 6184 6316
rect 6236 6264 6242 6316
rect 5169 6239 5227 6245
rect 5169 6205 5181 6239
rect 5215 6236 5227 6239
rect 6196 6236 6224 6264
rect 5215 6208 6224 6236
rect 6886 6236 6914 6344
rect 17405 6341 17417 6375
rect 17451 6372 17463 6375
rect 17494 6372 17500 6384
rect 17451 6344 17500 6372
rect 17451 6341 17463 6344
rect 17405 6335 17463 6341
rect 17494 6332 17500 6344
rect 17552 6332 17558 6384
rect 16666 6264 16672 6316
rect 16724 6264 16730 6316
rect 16758 6264 16764 6316
rect 16816 6264 16822 6316
rect 16942 6264 16948 6316
rect 17000 6264 17006 6316
rect 25222 6304 25228 6316
rect 17880 6276 25228 6304
rect 17880 6236 17908 6276
rect 25222 6264 25228 6276
rect 25280 6264 25286 6316
rect 31202 6264 31208 6316
rect 31260 6264 31266 6316
rect 31573 6307 31631 6313
rect 31573 6273 31585 6307
rect 31619 6304 31631 6307
rect 31662 6304 31668 6316
rect 31619 6276 31668 6304
rect 31619 6273 31631 6276
rect 31573 6267 31631 6273
rect 31662 6264 31668 6276
rect 31720 6264 31726 6316
rect 31846 6264 31852 6316
rect 31904 6264 31910 6316
rect 6886 6208 17908 6236
rect 5215 6205 5227 6208
rect 5169 6199 5227 6205
rect 18782 6196 18788 6248
rect 18840 6236 18846 6248
rect 34146 6236 34152 6248
rect 18840 6208 34152 6236
rect 18840 6196 18846 6208
rect 34146 6196 34152 6208
rect 34204 6196 34210 6248
rect 6089 6171 6147 6177
rect 6089 6137 6101 6171
rect 6135 6168 6147 6171
rect 29546 6168 29552 6180
rect 6135 6140 29552 6168
rect 6135 6137 6147 6140
rect 6089 6131 6147 6137
rect 29546 6128 29552 6140
rect 29604 6128 29610 6180
rect 1104 6010 40848 6032
rect 1104 5958 1950 6010
rect 2002 5958 2014 6010
rect 2066 5958 2078 6010
rect 2130 5958 2142 6010
rect 2194 5958 2206 6010
rect 2258 5958 6950 6010
rect 7002 5958 7014 6010
rect 7066 5958 7078 6010
rect 7130 5958 7142 6010
rect 7194 5958 7206 6010
rect 7258 5958 11950 6010
rect 12002 5958 12014 6010
rect 12066 5958 12078 6010
rect 12130 5958 12142 6010
rect 12194 5958 12206 6010
rect 12258 5958 16950 6010
rect 17002 5958 17014 6010
rect 17066 5958 17078 6010
rect 17130 5958 17142 6010
rect 17194 5958 17206 6010
rect 17258 5958 21950 6010
rect 22002 5958 22014 6010
rect 22066 5958 22078 6010
rect 22130 5958 22142 6010
rect 22194 5958 22206 6010
rect 22258 5958 26950 6010
rect 27002 5958 27014 6010
rect 27066 5958 27078 6010
rect 27130 5958 27142 6010
rect 27194 5958 27206 6010
rect 27258 5958 31950 6010
rect 32002 5958 32014 6010
rect 32066 5958 32078 6010
rect 32130 5958 32142 6010
rect 32194 5958 32206 6010
rect 32258 5958 36950 6010
rect 37002 5958 37014 6010
rect 37066 5958 37078 6010
rect 37130 5958 37142 6010
rect 37194 5958 37206 6010
rect 37258 5958 40848 6010
rect 1104 5936 40848 5958
rect 1104 5466 40848 5488
rect 1104 5414 2610 5466
rect 2662 5414 2674 5466
rect 2726 5414 2738 5466
rect 2790 5414 2802 5466
rect 2854 5414 2866 5466
rect 2918 5414 7610 5466
rect 7662 5414 7674 5466
rect 7726 5414 7738 5466
rect 7790 5414 7802 5466
rect 7854 5414 7866 5466
rect 7918 5414 12610 5466
rect 12662 5414 12674 5466
rect 12726 5414 12738 5466
rect 12790 5414 12802 5466
rect 12854 5414 12866 5466
rect 12918 5414 17610 5466
rect 17662 5414 17674 5466
rect 17726 5414 17738 5466
rect 17790 5414 17802 5466
rect 17854 5414 17866 5466
rect 17918 5414 22610 5466
rect 22662 5414 22674 5466
rect 22726 5414 22738 5466
rect 22790 5414 22802 5466
rect 22854 5414 22866 5466
rect 22918 5414 27610 5466
rect 27662 5414 27674 5466
rect 27726 5414 27738 5466
rect 27790 5414 27802 5466
rect 27854 5414 27866 5466
rect 27918 5414 32610 5466
rect 32662 5414 32674 5466
rect 32726 5414 32738 5466
rect 32790 5414 32802 5466
rect 32854 5414 32866 5466
rect 32918 5414 37610 5466
rect 37662 5414 37674 5466
rect 37726 5414 37738 5466
rect 37790 5414 37802 5466
rect 37854 5414 37866 5466
rect 37918 5414 40848 5466
rect 1104 5392 40848 5414
rect 3694 5312 3700 5364
rect 3752 5352 3758 5364
rect 12526 5352 12532 5364
rect 3752 5324 12532 5352
rect 3752 5312 3758 5324
rect 12526 5312 12532 5324
rect 12584 5352 12590 5364
rect 12986 5352 12992 5364
rect 12584 5324 12992 5352
rect 12584 5312 12590 5324
rect 12986 5312 12992 5324
rect 13044 5312 13050 5364
rect 8386 5244 8392 5296
rect 8444 5284 8450 5296
rect 8444 5256 16574 5284
rect 8444 5244 8450 5256
rect 8202 5176 8208 5228
rect 8260 5176 8266 5228
rect 8478 5176 8484 5228
rect 8536 5176 8542 5228
rect 8578 5219 8636 5225
rect 8578 5185 8590 5219
rect 8624 5185 8636 5219
rect 16546 5216 16574 5256
rect 22462 5216 22468 5228
rect 16546 5188 22468 5216
rect 8578 5179 8636 5185
rect 7282 5108 7288 5160
rect 7340 5148 7346 5160
rect 8588 5148 8616 5179
rect 22462 5176 22468 5188
rect 22520 5176 22526 5228
rect 7340 5120 8616 5148
rect 7340 5108 7346 5120
rect 8754 5040 8760 5092
rect 8812 5040 8818 5092
rect 19610 5080 19616 5092
rect 16546 5052 19616 5080
rect 4338 4972 4344 5024
rect 4396 5012 4402 5024
rect 8110 5012 8116 5024
rect 4396 4984 8116 5012
rect 4396 4972 4402 4984
rect 8110 4972 8116 4984
rect 8168 5012 8174 5024
rect 16546 5012 16574 5052
rect 19610 5040 19616 5052
rect 19668 5040 19674 5092
rect 8168 4984 16574 5012
rect 8168 4972 8174 4984
rect 31018 4972 31024 5024
rect 31076 5012 31082 5024
rect 37458 5012 37464 5024
rect 31076 4984 37464 5012
rect 31076 4972 31082 4984
rect 37458 4972 37464 4984
rect 37516 5012 37522 5024
rect 38562 5012 38568 5024
rect 37516 4984 38568 5012
rect 37516 4972 37522 4984
rect 38562 4972 38568 4984
rect 38620 4972 38626 5024
rect 1104 4922 40848 4944
rect 1104 4870 1950 4922
rect 2002 4870 2014 4922
rect 2066 4870 2078 4922
rect 2130 4870 2142 4922
rect 2194 4870 2206 4922
rect 2258 4870 6950 4922
rect 7002 4870 7014 4922
rect 7066 4870 7078 4922
rect 7130 4870 7142 4922
rect 7194 4870 7206 4922
rect 7258 4870 11950 4922
rect 12002 4870 12014 4922
rect 12066 4870 12078 4922
rect 12130 4870 12142 4922
rect 12194 4870 12206 4922
rect 12258 4870 16950 4922
rect 17002 4870 17014 4922
rect 17066 4870 17078 4922
rect 17130 4870 17142 4922
rect 17194 4870 17206 4922
rect 17258 4870 21950 4922
rect 22002 4870 22014 4922
rect 22066 4870 22078 4922
rect 22130 4870 22142 4922
rect 22194 4870 22206 4922
rect 22258 4870 26950 4922
rect 27002 4870 27014 4922
rect 27066 4870 27078 4922
rect 27130 4870 27142 4922
rect 27194 4870 27206 4922
rect 27258 4870 31950 4922
rect 32002 4870 32014 4922
rect 32066 4870 32078 4922
rect 32130 4870 32142 4922
rect 32194 4870 32206 4922
rect 32258 4870 36950 4922
rect 37002 4870 37014 4922
rect 37066 4870 37078 4922
rect 37130 4870 37142 4922
rect 37194 4870 37206 4922
rect 37258 4870 40848 4922
rect 1104 4848 40848 4870
rect 7193 4811 7251 4817
rect 7193 4777 7205 4811
rect 7239 4808 7251 4811
rect 7374 4808 7380 4820
rect 7239 4780 7380 4808
rect 7239 4777 7251 4780
rect 7193 4771 7251 4777
rect 7374 4768 7380 4780
rect 7432 4768 7438 4820
rect 31018 4808 31024 4820
rect 16546 4780 31024 4808
rect 8386 4740 8392 4752
rect 6748 4712 8392 4740
rect 2225 4675 2283 4681
rect 2225 4641 2237 4675
rect 2271 4672 2283 4675
rect 3694 4672 3700 4684
rect 2271 4644 3700 4672
rect 2271 4641 2283 4644
rect 2225 4635 2283 4641
rect 3694 4632 3700 4644
rect 3752 4632 3758 4684
rect 3786 4632 3792 4684
rect 3844 4632 3850 4684
rect 6748 4681 6776 4712
rect 8386 4700 8392 4712
rect 8444 4700 8450 4752
rect 16546 4740 16574 4780
rect 31018 4768 31024 4780
rect 31076 4768 31082 4820
rect 35618 4768 35624 4820
rect 35676 4808 35682 4820
rect 35676 4780 38424 4808
rect 35676 4768 35682 4780
rect 15764 4712 16574 4740
rect 6733 4675 6791 4681
rect 6733 4672 6745 4675
rect 4172 4644 6745 4672
rect 842 4564 848 4616
rect 900 4604 906 4616
rect 1397 4607 1455 4613
rect 1397 4604 1409 4607
rect 900 4576 1409 4604
rect 900 4564 906 4576
rect 1397 4573 1409 4576
rect 1443 4573 1455 4607
rect 1397 4567 1455 4573
rect 4172 4545 4200 4644
rect 6733 4641 6745 4644
rect 6779 4641 6791 4675
rect 7466 4672 7472 4684
rect 6733 4635 6791 4641
rect 6932 4644 7472 4672
rect 4338 4564 4344 4616
rect 4396 4564 4402 4616
rect 6086 4564 6092 4616
rect 6144 4604 6150 4616
rect 6932 4613 6960 4644
rect 7466 4632 7472 4644
rect 7524 4632 7530 4684
rect 14090 4632 14096 4684
rect 14148 4632 14154 4684
rect 6641 4607 6699 4613
rect 6641 4604 6653 4607
rect 6144 4576 6653 4604
rect 6144 4564 6150 4576
rect 6641 4573 6653 4576
rect 6687 4573 6699 4607
rect 6641 4567 6699 4573
rect 6917 4607 6975 4613
rect 6917 4573 6929 4607
rect 6963 4573 6975 4607
rect 6917 4567 6975 4573
rect 7006 4564 7012 4616
rect 7064 4604 7070 4616
rect 8202 4604 8208 4616
rect 7064 4576 8208 4604
rect 7064 4564 7070 4576
rect 8202 4564 8208 4576
rect 8260 4564 8266 4616
rect 14274 4564 14280 4616
rect 14332 4564 14338 4616
rect 14921 4607 14979 4613
rect 14921 4573 14933 4607
rect 14967 4573 14979 4607
rect 14921 4567 14979 4573
rect 15289 4607 15347 4613
rect 15289 4573 15301 4607
rect 15335 4604 15347 4607
rect 15764 4604 15792 4712
rect 15335 4576 15792 4604
rect 16546 4644 19932 4672
rect 15335 4573 15347 4576
rect 15289 4567 15347 4573
rect 4157 4539 4215 4545
rect 4157 4505 4169 4539
rect 4203 4505 4215 4539
rect 4157 4499 4215 4505
rect 4249 4539 4307 4545
rect 4249 4505 4261 4539
rect 4295 4536 4307 4539
rect 4525 4539 4583 4545
rect 4295 4508 4476 4536
rect 4295 4505 4307 4508
rect 4249 4499 4307 4505
rect 4448 4468 4476 4508
rect 4525 4505 4537 4539
rect 4571 4536 4583 4539
rect 6270 4536 6276 4548
rect 4571 4508 6276 4536
rect 4571 4505 4583 4508
rect 4525 4499 4583 4505
rect 6270 4496 6276 4508
rect 6328 4496 6334 4548
rect 14936 4536 14964 4567
rect 16546 4536 16574 4644
rect 18598 4564 18604 4616
rect 18656 4604 18662 4616
rect 19429 4607 19487 4613
rect 19429 4604 19441 4607
rect 18656 4576 19441 4604
rect 18656 4564 18662 4576
rect 19429 4573 19441 4576
rect 19475 4573 19487 4607
rect 19429 4567 19487 4573
rect 19518 4564 19524 4616
rect 19576 4564 19582 4616
rect 19904 4604 19932 4644
rect 19978 4632 19984 4684
rect 20036 4632 20042 4684
rect 26418 4632 26424 4684
rect 26476 4672 26482 4684
rect 26476 4644 35894 4672
rect 26476 4632 26482 4644
rect 34698 4604 34704 4616
rect 19904 4576 34704 4604
rect 34698 4564 34704 4576
rect 34756 4564 34762 4616
rect 35866 4604 35894 4644
rect 37366 4632 37372 4684
rect 37424 4632 37430 4684
rect 38102 4672 38108 4684
rect 37752 4644 38108 4672
rect 37752 4613 37780 4644
rect 38102 4632 38108 4644
rect 38160 4632 38166 4684
rect 38396 4613 38424 4780
rect 38562 4700 38568 4752
rect 38620 4700 38626 4752
rect 37461 4607 37519 4613
rect 37461 4604 37473 4607
rect 35866 4576 37473 4604
rect 37461 4573 37473 4576
rect 37507 4573 37519 4607
rect 37461 4567 37519 4573
rect 37737 4607 37795 4613
rect 37737 4573 37749 4607
rect 37783 4573 37795 4607
rect 37737 4567 37795 4573
rect 37921 4607 37979 4613
rect 37921 4573 37933 4607
rect 37967 4573 37979 4607
rect 37921 4567 37979 4573
rect 38013 4607 38071 4613
rect 38013 4573 38025 4607
rect 38059 4573 38071 4607
rect 38013 4567 38071 4573
rect 38381 4607 38439 4613
rect 38381 4573 38393 4607
rect 38427 4573 38439 4607
rect 38381 4567 38439 4573
rect 14936 4508 16574 4536
rect 18230 4496 18236 4548
rect 18288 4536 18294 4548
rect 19245 4539 19303 4545
rect 19245 4536 19257 4539
rect 18288 4508 19257 4536
rect 18288 4496 18294 4508
rect 19245 4505 19257 4508
rect 19291 4505 19303 4539
rect 19245 4499 19303 4505
rect 19610 4496 19616 4548
rect 19668 4496 19674 4548
rect 37274 4496 37280 4548
rect 37332 4536 37338 4548
rect 37936 4536 37964 4567
rect 37332 4508 37964 4536
rect 37332 4496 37338 4508
rect 7282 4468 7288 4480
rect 4448 4440 7288 4468
rect 7282 4428 7288 4440
rect 7340 4428 7346 4480
rect 35526 4428 35532 4480
rect 35584 4468 35590 4480
rect 38028 4468 38056 4567
rect 35584 4440 38056 4468
rect 35584 4428 35590 4440
rect 1104 4378 40848 4400
rect 1104 4326 2610 4378
rect 2662 4326 2674 4378
rect 2726 4326 2738 4378
rect 2790 4326 2802 4378
rect 2854 4326 2866 4378
rect 2918 4326 7610 4378
rect 7662 4326 7674 4378
rect 7726 4326 7738 4378
rect 7790 4326 7802 4378
rect 7854 4326 7866 4378
rect 7918 4326 12610 4378
rect 12662 4326 12674 4378
rect 12726 4326 12738 4378
rect 12790 4326 12802 4378
rect 12854 4326 12866 4378
rect 12918 4326 17610 4378
rect 17662 4326 17674 4378
rect 17726 4326 17738 4378
rect 17790 4326 17802 4378
rect 17854 4326 17866 4378
rect 17918 4326 22610 4378
rect 22662 4326 22674 4378
rect 22726 4326 22738 4378
rect 22790 4326 22802 4378
rect 22854 4326 22866 4378
rect 22918 4326 27610 4378
rect 27662 4326 27674 4378
rect 27726 4326 27738 4378
rect 27790 4326 27802 4378
rect 27854 4326 27866 4378
rect 27918 4326 32610 4378
rect 32662 4326 32674 4378
rect 32726 4326 32738 4378
rect 32790 4326 32802 4378
rect 32854 4326 32866 4378
rect 32918 4326 37610 4378
rect 37662 4326 37674 4378
rect 37726 4326 37738 4378
rect 37790 4326 37802 4378
rect 37854 4326 37866 4378
rect 37918 4326 40848 4378
rect 1104 4304 40848 4326
rect 40494 4156 40500 4208
rect 40552 4156 40558 4208
rect 6454 4088 6460 4140
rect 6512 4088 6518 4140
rect 7561 4131 7619 4137
rect 7561 4097 7573 4131
rect 7607 4128 7619 4131
rect 9214 4128 9220 4140
rect 7607 4100 9220 4128
rect 7607 4097 7619 4100
rect 7561 4091 7619 4097
rect 9214 4088 9220 4100
rect 9272 4088 9278 4140
rect 34146 4088 34152 4140
rect 34204 4088 34210 4140
rect 7469 4063 7527 4069
rect 7469 4029 7481 4063
rect 7515 4060 7527 4063
rect 8846 4060 8852 4072
rect 7515 4032 8852 4060
rect 7515 4029 7527 4032
rect 7469 4023 7527 4029
rect 8846 4020 8852 4032
rect 8904 4020 8910 4072
rect 36814 4020 36820 4072
rect 36872 4060 36878 4072
rect 39669 4063 39727 4069
rect 39669 4060 39681 4063
rect 36872 4032 39681 4060
rect 36872 4020 36878 4032
rect 39669 4029 39681 4032
rect 39715 4029 39727 4063
rect 39669 4023 39727 4029
rect 1104 3834 40848 3856
rect 1104 3782 1950 3834
rect 2002 3782 2014 3834
rect 2066 3782 2078 3834
rect 2130 3782 2142 3834
rect 2194 3782 2206 3834
rect 2258 3782 6950 3834
rect 7002 3782 7014 3834
rect 7066 3782 7078 3834
rect 7130 3782 7142 3834
rect 7194 3782 7206 3834
rect 7258 3782 11950 3834
rect 12002 3782 12014 3834
rect 12066 3782 12078 3834
rect 12130 3782 12142 3834
rect 12194 3782 12206 3834
rect 12258 3782 16950 3834
rect 17002 3782 17014 3834
rect 17066 3782 17078 3834
rect 17130 3782 17142 3834
rect 17194 3782 17206 3834
rect 17258 3782 21950 3834
rect 22002 3782 22014 3834
rect 22066 3782 22078 3834
rect 22130 3782 22142 3834
rect 22194 3782 22206 3834
rect 22258 3782 26950 3834
rect 27002 3782 27014 3834
rect 27066 3782 27078 3834
rect 27130 3782 27142 3834
rect 27194 3782 27206 3834
rect 27258 3782 31950 3834
rect 32002 3782 32014 3834
rect 32066 3782 32078 3834
rect 32130 3782 32142 3834
rect 32194 3782 32206 3834
rect 32258 3782 36950 3834
rect 37002 3782 37014 3834
rect 37066 3782 37078 3834
rect 37130 3782 37142 3834
rect 37194 3782 37206 3834
rect 37258 3782 40848 3834
rect 1104 3760 40848 3782
rect 8220 3692 16574 3720
rect 4798 3476 4804 3528
rect 4856 3516 4862 3528
rect 8220 3525 8248 3692
rect 10962 3612 10968 3664
rect 11020 3612 11026 3664
rect 16546 3652 16574 3692
rect 34146 3680 34152 3732
rect 34204 3680 34210 3732
rect 33686 3652 33692 3664
rect 16546 3624 33692 3652
rect 33686 3612 33692 3624
rect 33744 3612 33750 3664
rect 10321 3587 10379 3593
rect 10321 3553 10333 3587
rect 10367 3584 10379 3587
rect 10870 3584 10876 3596
rect 10367 3556 10876 3584
rect 10367 3553 10379 3556
rect 10321 3547 10379 3553
rect 10870 3544 10876 3556
rect 10928 3544 10934 3596
rect 35894 3584 35900 3596
rect 13372 3556 35900 3584
rect 7193 3519 7251 3525
rect 7193 3516 7205 3519
rect 4856 3488 7205 3516
rect 4856 3476 4862 3488
rect 7193 3485 7205 3488
rect 7239 3485 7251 3519
rect 7193 3479 7251 3485
rect 8205 3519 8263 3525
rect 8205 3485 8217 3519
rect 8251 3485 8263 3519
rect 8205 3479 8263 3485
rect 10413 3519 10471 3525
rect 10413 3485 10425 3519
rect 10459 3485 10471 3519
rect 10413 3479 10471 3485
rect 8018 3408 8024 3460
rect 8076 3448 8082 3460
rect 10428 3448 10456 3479
rect 11146 3476 11152 3528
rect 11204 3476 11210 3528
rect 12526 3476 12532 3528
rect 12584 3516 12590 3528
rect 13372 3525 13400 3556
rect 35894 3544 35900 3556
rect 35952 3584 35958 3596
rect 36814 3584 36820 3596
rect 35952 3556 36820 3584
rect 35952 3544 35958 3556
rect 36814 3544 36820 3556
rect 36872 3544 36878 3596
rect 12805 3519 12863 3525
rect 12805 3516 12817 3519
rect 12584 3488 12817 3516
rect 12584 3476 12590 3488
rect 12805 3485 12817 3488
rect 12851 3485 12863 3519
rect 12805 3479 12863 3485
rect 13357 3519 13415 3525
rect 13357 3485 13369 3519
rect 13403 3485 13415 3519
rect 13357 3479 13415 3485
rect 13633 3519 13691 3525
rect 13633 3485 13645 3519
rect 13679 3485 13691 3519
rect 13633 3479 13691 3485
rect 13909 3519 13967 3525
rect 13909 3485 13921 3519
rect 13955 3516 13967 3519
rect 14458 3516 14464 3528
rect 13955 3488 14464 3516
rect 13955 3485 13967 3488
rect 13909 3479 13967 3485
rect 8076 3420 10456 3448
rect 8076 3408 8082 3420
rect 8202 3340 8208 3392
rect 8260 3380 8266 3392
rect 13648 3380 13676 3479
rect 14458 3476 14464 3488
rect 14516 3476 14522 3528
rect 8260 3352 13676 3380
rect 8260 3340 8266 3352
rect 26050 3340 26056 3392
rect 26108 3380 26114 3392
rect 29638 3380 29644 3392
rect 26108 3352 29644 3380
rect 26108 3340 26114 3352
rect 29638 3340 29644 3352
rect 29696 3340 29702 3392
rect 1104 3290 40848 3312
rect 1104 3238 2610 3290
rect 2662 3238 2674 3290
rect 2726 3238 2738 3290
rect 2790 3238 2802 3290
rect 2854 3238 2866 3290
rect 2918 3238 7610 3290
rect 7662 3238 7674 3290
rect 7726 3238 7738 3290
rect 7790 3238 7802 3290
rect 7854 3238 7866 3290
rect 7918 3238 12610 3290
rect 12662 3238 12674 3290
rect 12726 3238 12738 3290
rect 12790 3238 12802 3290
rect 12854 3238 12866 3290
rect 12918 3238 17610 3290
rect 17662 3238 17674 3290
rect 17726 3238 17738 3290
rect 17790 3238 17802 3290
rect 17854 3238 17866 3290
rect 17918 3238 22610 3290
rect 22662 3238 22674 3290
rect 22726 3238 22738 3290
rect 22790 3238 22802 3290
rect 22854 3238 22866 3290
rect 22918 3238 27610 3290
rect 27662 3238 27674 3290
rect 27726 3238 27738 3290
rect 27790 3238 27802 3290
rect 27854 3238 27866 3290
rect 27918 3238 32610 3290
rect 32662 3238 32674 3290
rect 32726 3238 32738 3290
rect 32790 3238 32802 3290
rect 32854 3238 32866 3290
rect 32918 3238 37610 3290
rect 37662 3238 37674 3290
rect 37726 3238 37738 3290
rect 37790 3238 37802 3290
rect 37854 3238 37866 3290
rect 37918 3238 40848 3290
rect 1104 3216 40848 3238
rect 8478 3136 8484 3188
rect 8536 3176 8542 3188
rect 8536 3148 26234 3176
rect 8536 3136 8542 3148
rect 26206 3108 26234 3148
rect 27522 3136 27528 3188
rect 27580 3176 27586 3188
rect 27580 3148 28580 3176
rect 27580 3136 27586 3148
rect 28552 3117 28580 3148
rect 34146 3136 34152 3188
rect 34204 3136 34210 3188
rect 28537 3111 28595 3117
rect 26206 3080 28396 3108
rect 28166 3000 28172 3052
rect 28224 3000 28230 3052
rect 20070 2932 20076 2984
rect 20128 2972 20134 2984
rect 27982 2972 27988 2984
rect 20128 2944 27988 2972
rect 20128 2932 20134 2944
rect 27982 2932 27988 2944
rect 28040 2932 28046 2984
rect 28368 2972 28396 3080
rect 28537 3077 28549 3111
rect 28583 3077 28595 3111
rect 28537 3071 28595 3077
rect 29638 3068 29644 3120
rect 29696 3068 29702 3120
rect 28626 3000 28632 3052
rect 28684 3000 28690 3052
rect 28721 3043 28779 3049
rect 28721 3009 28733 3043
rect 28767 3009 28779 3043
rect 28721 3003 28779 3009
rect 28905 3043 28963 3049
rect 28905 3009 28917 3043
rect 28951 3040 28963 3043
rect 33226 3040 33232 3052
rect 28951 3012 33232 3040
rect 28951 3009 28963 3012
rect 28905 3003 28963 3009
rect 28736 2972 28764 3003
rect 33226 3000 33232 3012
rect 33284 3000 33290 3052
rect 28368 2944 28764 2972
rect 26326 2864 26332 2916
rect 26384 2904 26390 2916
rect 29917 2907 29975 2913
rect 29917 2904 29929 2907
rect 26384 2876 29929 2904
rect 26384 2864 26390 2876
rect 29917 2873 29929 2876
rect 29963 2873 29975 2907
rect 29917 2867 29975 2873
rect 17310 2796 17316 2848
rect 17368 2836 17374 2848
rect 30101 2839 30159 2845
rect 30101 2836 30113 2839
rect 17368 2808 30113 2836
rect 17368 2796 17374 2808
rect 30101 2805 30113 2808
rect 30147 2805 30159 2839
rect 30101 2799 30159 2805
rect 1104 2746 40848 2768
rect 1104 2694 1950 2746
rect 2002 2694 2014 2746
rect 2066 2694 2078 2746
rect 2130 2694 2142 2746
rect 2194 2694 2206 2746
rect 2258 2694 6950 2746
rect 7002 2694 7014 2746
rect 7066 2694 7078 2746
rect 7130 2694 7142 2746
rect 7194 2694 7206 2746
rect 7258 2694 11950 2746
rect 12002 2694 12014 2746
rect 12066 2694 12078 2746
rect 12130 2694 12142 2746
rect 12194 2694 12206 2746
rect 12258 2694 16950 2746
rect 17002 2694 17014 2746
rect 17066 2694 17078 2746
rect 17130 2694 17142 2746
rect 17194 2694 17206 2746
rect 17258 2694 21950 2746
rect 22002 2694 22014 2746
rect 22066 2694 22078 2746
rect 22130 2694 22142 2746
rect 22194 2694 22206 2746
rect 22258 2694 26950 2746
rect 27002 2694 27014 2746
rect 27066 2694 27078 2746
rect 27130 2694 27142 2746
rect 27194 2694 27206 2746
rect 27258 2694 31950 2746
rect 32002 2694 32014 2746
rect 32066 2694 32078 2746
rect 32130 2694 32142 2746
rect 32194 2694 32206 2746
rect 32258 2694 36950 2746
rect 37002 2694 37014 2746
rect 37066 2694 37078 2746
rect 37130 2694 37142 2746
rect 37194 2694 37206 2746
rect 37258 2694 40848 2746
rect 1104 2672 40848 2694
rect 24578 2632 24584 2644
rect 13464 2604 24584 2632
rect 2498 2456 2504 2508
rect 2556 2456 2562 2508
rect 11698 2496 11704 2508
rect 2976 2468 11704 2496
rect 2976 2437 3004 2468
rect 11698 2456 11704 2468
rect 11756 2456 11762 2508
rect 2961 2431 3019 2437
rect 2961 2397 2973 2431
rect 3007 2397 3019 2431
rect 2961 2391 3019 2397
rect 8113 2431 8171 2437
rect 8113 2397 8125 2431
rect 8159 2428 8171 2431
rect 10134 2428 10140 2440
rect 8159 2400 10140 2428
rect 8159 2397 8171 2400
rect 8113 2391 8171 2397
rect 10134 2388 10140 2400
rect 10192 2388 10198 2440
rect 13464 2437 13492 2604
rect 24578 2592 24584 2604
rect 24636 2592 24642 2644
rect 14366 2524 14372 2576
rect 14424 2564 14430 2576
rect 39025 2567 39083 2573
rect 39025 2564 39037 2567
rect 14424 2536 39037 2564
rect 14424 2524 14430 2536
rect 39025 2533 39037 2536
rect 39071 2533 39083 2567
rect 39025 2527 39083 2533
rect 34606 2496 34612 2508
rect 18708 2468 34612 2496
rect 18708 2437 18736 2468
rect 34606 2456 34612 2468
rect 34664 2456 34670 2508
rect 13449 2431 13507 2437
rect 13449 2397 13461 2431
rect 13495 2397 13507 2431
rect 13449 2391 13507 2397
rect 18141 2431 18199 2437
rect 18141 2397 18153 2431
rect 18187 2428 18199 2431
rect 18693 2431 18751 2437
rect 18693 2428 18705 2431
rect 18187 2400 18705 2428
rect 18187 2397 18199 2400
rect 18141 2391 18199 2397
rect 18693 2397 18705 2400
rect 18739 2397 18751 2431
rect 23661 2431 23719 2437
rect 23661 2428 23673 2431
rect 18693 2391 18751 2397
rect 23308 2400 23673 2428
rect 7745 2363 7803 2369
rect 7745 2329 7757 2363
rect 7791 2360 7803 2363
rect 8018 2360 8024 2372
rect 7791 2332 8024 2360
rect 7791 2329 7803 2332
rect 7745 2323 7803 2329
rect 8018 2320 8024 2332
rect 8076 2320 8082 2372
rect 23308 2369 23336 2400
rect 23661 2397 23673 2400
rect 23707 2397 23719 2431
rect 28997 2431 29055 2437
rect 28997 2428 29009 2431
rect 23661 2391 23719 2397
rect 28644 2400 29009 2428
rect 28644 2372 28672 2400
rect 28997 2397 29009 2400
rect 29043 2397 29055 2431
rect 28997 2391 29055 2397
rect 34146 2388 34152 2440
rect 34204 2388 34210 2440
rect 39040 2428 39068 2527
rect 39393 2431 39451 2437
rect 39393 2428 39405 2431
rect 39040 2400 39405 2428
rect 39393 2397 39405 2400
rect 39439 2397 39451 2431
rect 39393 2391 39451 2397
rect 23293 2363 23351 2369
rect 23293 2360 23305 2363
rect 11716 2332 23305 2360
rect 2314 2252 2320 2304
rect 2372 2292 2378 2304
rect 11716 2292 11744 2332
rect 23293 2329 23305 2332
rect 23339 2329 23351 2363
rect 23293 2323 23351 2329
rect 28626 2320 28632 2372
rect 28684 2320 28690 2372
rect 2372 2264 11744 2292
rect 2372 2252 2378 2264
rect 13078 2252 13084 2304
rect 13136 2292 13142 2304
rect 13265 2295 13323 2301
rect 13265 2292 13277 2295
rect 13136 2264 13277 2292
rect 13136 2252 13142 2264
rect 13265 2261 13277 2264
rect 13311 2261 13323 2295
rect 13265 2255 13323 2261
rect 18322 2252 18328 2304
rect 18380 2292 18386 2304
rect 18509 2295 18567 2301
rect 18509 2292 18521 2295
rect 18380 2264 18521 2292
rect 18380 2252 18386 2264
rect 18509 2261 18521 2264
rect 18555 2261 18567 2295
rect 18509 2255 18567 2261
rect 23566 2252 23572 2304
rect 23624 2292 23630 2304
rect 23845 2295 23903 2301
rect 23845 2292 23857 2295
rect 23624 2264 23857 2292
rect 23624 2252 23630 2264
rect 23845 2261 23857 2264
rect 23891 2261 23903 2295
rect 23845 2255 23903 2261
rect 28810 2252 28816 2304
rect 28868 2292 28874 2304
rect 29181 2295 29239 2301
rect 29181 2292 29193 2295
rect 28868 2264 29193 2292
rect 28868 2252 28874 2264
rect 29181 2261 29193 2264
rect 29227 2261 29239 2295
rect 29181 2255 29239 2261
rect 34054 2252 34060 2304
rect 34112 2292 34118 2304
rect 34333 2295 34391 2301
rect 34333 2292 34345 2295
rect 34112 2264 34345 2292
rect 34112 2252 34118 2264
rect 34333 2261 34345 2264
rect 34379 2261 34391 2295
rect 34333 2255 34391 2261
rect 39298 2252 39304 2304
rect 39356 2292 39362 2304
rect 39577 2295 39635 2301
rect 39577 2292 39589 2295
rect 39356 2264 39589 2292
rect 39356 2252 39362 2264
rect 39577 2261 39589 2264
rect 39623 2261 39635 2295
rect 39577 2255 39635 2261
rect 1104 2202 40848 2224
rect 1104 2150 2610 2202
rect 2662 2150 2674 2202
rect 2726 2150 2738 2202
rect 2790 2150 2802 2202
rect 2854 2150 2866 2202
rect 2918 2150 7610 2202
rect 7662 2150 7674 2202
rect 7726 2150 7738 2202
rect 7790 2150 7802 2202
rect 7854 2150 7866 2202
rect 7918 2150 12610 2202
rect 12662 2150 12674 2202
rect 12726 2150 12738 2202
rect 12790 2150 12802 2202
rect 12854 2150 12866 2202
rect 12918 2150 17610 2202
rect 17662 2150 17674 2202
rect 17726 2150 17738 2202
rect 17790 2150 17802 2202
rect 17854 2150 17866 2202
rect 17918 2150 22610 2202
rect 22662 2150 22674 2202
rect 22726 2150 22738 2202
rect 22790 2150 22802 2202
rect 22854 2150 22866 2202
rect 22918 2150 27610 2202
rect 27662 2150 27674 2202
rect 27726 2150 27738 2202
rect 27790 2150 27802 2202
rect 27854 2150 27866 2202
rect 27918 2150 32610 2202
rect 32662 2150 32674 2202
rect 32726 2150 32738 2202
rect 32790 2150 32802 2202
rect 32854 2150 32866 2202
rect 32918 2150 37610 2202
rect 37662 2150 37674 2202
rect 37726 2150 37738 2202
rect 37790 2150 37802 2202
rect 37854 2150 37866 2202
rect 37918 2150 40848 2202
rect 1104 2128 40848 2150
<< via1 >>
rect 2610 69606 2662 69658
rect 2674 69606 2726 69658
rect 2738 69606 2790 69658
rect 2802 69606 2854 69658
rect 2866 69606 2918 69658
rect 7610 69606 7662 69658
rect 7674 69606 7726 69658
rect 7738 69606 7790 69658
rect 7802 69606 7854 69658
rect 7866 69606 7918 69658
rect 12610 69606 12662 69658
rect 12674 69606 12726 69658
rect 12738 69606 12790 69658
rect 12802 69606 12854 69658
rect 12866 69606 12918 69658
rect 17610 69606 17662 69658
rect 17674 69606 17726 69658
rect 17738 69606 17790 69658
rect 17802 69606 17854 69658
rect 17866 69606 17918 69658
rect 22610 69606 22662 69658
rect 22674 69606 22726 69658
rect 22738 69606 22790 69658
rect 22802 69606 22854 69658
rect 22866 69606 22918 69658
rect 27610 69606 27662 69658
rect 27674 69606 27726 69658
rect 27738 69606 27790 69658
rect 27802 69606 27854 69658
rect 27866 69606 27918 69658
rect 32610 69606 32662 69658
rect 32674 69606 32726 69658
rect 32738 69606 32790 69658
rect 32802 69606 32854 69658
rect 32866 69606 32918 69658
rect 37610 69606 37662 69658
rect 37674 69606 37726 69658
rect 37738 69606 37790 69658
rect 37802 69606 37854 69658
rect 37866 69606 37918 69658
rect 34980 69479 35032 69488
rect 34980 69445 34989 69479
rect 34989 69445 35023 69479
rect 35023 69445 35032 69479
rect 34980 69436 35032 69445
rect 7104 69411 7156 69420
rect 7104 69377 7113 69411
rect 7113 69377 7147 69411
rect 7147 69377 7156 69411
rect 7104 69368 7156 69377
rect 20904 69368 20956 69420
rect 9588 69300 9640 69352
rect 22376 69343 22428 69352
rect 22376 69309 22385 69343
rect 22385 69309 22419 69343
rect 22419 69309 22428 69343
rect 22376 69300 22428 69309
rect 35440 69300 35492 69352
rect 1950 69062 2002 69114
rect 2014 69062 2066 69114
rect 2078 69062 2130 69114
rect 2142 69062 2194 69114
rect 2206 69062 2258 69114
rect 6950 69062 7002 69114
rect 7014 69062 7066 69114
rect 7078 69062 7130 69114
rect 7142 69062 7194 69114
rect 7206 69062 7258 69114
rect 11950 69062 12002 69114
rect 12014 69062 12066 69114
rect 12078 69062 12130 69114
rect 12142 69062 12194 69114
rect 12206 69062 12258 69114
rect 16950 69062 17002 69114
rect 17014 69062 17066 69114
rect 17078 69062 17130 69114
rect 17142 69062 17194 69114
rect 17206 69062 17258 69114
rect 21950 69062 22002 69114
rect 22014 69062 22066 69114
rect 22078 69062 22130 69114
rect 22142 69062 22194 69114
rect 22206 69062 22258 69114
rect 26950 69062 27002 69114
rect 27014 69062 27066 69114
rect 27078 69062 27130 69114
rect 27142 69062 27194 69114
rect 27206 69062 27258 69114
rect 31950 69062 32002 69114
rect 32014 69062 32066 69114
rect 32078 69062 32130 69114
rect 32142 69062 32194 69114
rect 32206 69062 32258 69114
rect 36950 69062 37002 69114
rect 37014 69062 37066 69114
rect 37078 69062 37130 69114
rect 37142 69062 37194 69114
rect 37206 69062 37258 69114
rect 11428 68756 11480 68808
rect 11520 68688 11572 68740
rect 13176 68756 13228 68808
rect 15568 68756 15620 68808
rect 28724 68756 28776 68808
rect 31484 68799 31536 68808
rect 31484 68765 31493 68799
rect 31493 68765 31527 68799
rect 31527 68765 31536 68799
rect 31484 68756 31536 68765
rect 13268 68688 13320 68740
rect 20168 68620 20220 68672
rect 31116 68663 31168 68672
rect 31116 68629 31125 68663
rect 31125 68629 31159 68663
rect 31159 68629 31168 68663
rect 31116 68620 31168 68629
rect 2610 68518 2662 68570
rect 2674 68518 2726 68570
rect 2738 68518 2790 68570
rect 2802 68518 2854 68570
rect 2866 68518 2918 68570
rect 7610 68518 7662 68570
rect 7674 68518 7726 68570
rect 7738 68518 7790 68570
rect 7802 68518 7854 68570
rect 7866 68518 7918 68570
rect 12610 68518 12662 68570
rect 12674 68518 12726 68570
rect 12738 68518 12790 68570
rect 12802 68518 12854 68570
rect 12866 68518 12918 68570
rect 17610 68518 17662 68570
rect 17674 68518 17726 68570
rect 17738 68518 17790 68570
rect 17802 68518 17854 68570
rect 17866 68518 17918 68570
rect 22610 68518 22662 68570
rect 22674 68518 22726 68570
rect 22738 68518 22790 68570
rect 22802 68518 22854 68570
rect 22866 68518 22918 68570
rect 27610 68518 27662 68570
rect 27674 68518 27726 68570
rect 27738 68518 27790 68570
rect 27802 68518 27854 68570
rect 27866 68518 27918 68570
rect 32610 68518 32662 68570
rect 32674 68518 32726 68570
rect 32738 68518 32790 68570
rect 32802 68518 32854 68570
rect 32866 68518 32918 68570
rect 37610 68518 37662 68570
rect 37674 68518 37726 68570
rect 37738 68518 37790 68570
rect 37802 68518 37854 68570
rect 37866 68518 37918 68570
rect 23848 68348 23900 68400
rect 19800 68280 19852 68332
rect 23112 68280 23164 68332
rect 1950 67974 2002 68026
rect 2014 67974 2066 68026
rect 2078 67974 2130 68026
rect 2142 67974 2194 68026
rect 2206 67974 2258 68026
rect 6950 67974 7002 68026
rect 7014 67974 7066 68026
rect 7078 67974 7130 68026
rect 7142 67974 7194 68026
rect 7206 67974 7258 68026
rect 11950 67974 12002 68026
rect 12014 67974 12066 68026
rect 12078 67974 12130 68026
rect 12142 67974 12194 68026
rect 12206 67974 12258 68026
rect 16950 67974 17002 68026
rect 17014 67974 17066 68026
rect 17078 67974 17130 68026
rect 17142 67974 17194 68026
rect 17206 67974 17258 68026
rect 21950 67974 22002 68026
rect 22014 67974 22066 68026
rect 22078 67974 22130 68026
rect 22142 67974 22194 68026
rect 22206 67974 22258 68026
rect 26950 67974 27002 68026
rect 27014 67974 27066 68026
rect 27078 67974 27130 68026
rect 27142 67974 27194 68026
rect 27206 67974 27258 68026
rect 31950 67974 32002 68026
rect 32014 67974 32066 68026
rect 32078 67974 32130 68026
rect 32142 67974 32194 68026
rect 32206 67974 32258 68026
rect 36950 67974 37002 68026
rect 37014 67974 37066 68026
rect 37078 67974 37130 68026
rect 37142 67974 37194 68026
rect 37206 67974 37258 68026
rect 8944 67872 8996 67924
rect 35348 67872 35400 67924
rect 13636 67804 13688 67856
rect 1400 67711 1452 67720
rect 1400 67677 1409 67711
rect 1409 67677 1443 67711
rect 1443 67677 1452 67711
rect 1400 67668 1452 67677
rect 26148 67736 26200 67788
rect 6552 67600 6604 67652
rect 13084 67668 13136 67720
rect 13452 67711 13504 67720
rect 13452 67677 13461 67711
rect 13461 67677 13495 67711
rect 13495 67677 13504 67711
rect 13452 67668 13504 67677
rect 13544 67711 13596 67720
rect 13544 67677 13553 67711
rect 13553 67677 13587 67711
rect 13587 67677 13596 67711
rect 13544 67668 13596 67677
rect 35256 67711 35308 67720
rect 35256 67677 35265 67711
rect 35265 67677 35299 67711
rect 35299 67677 35308 67711
rect 35256 67668 35308 67677
rect 38016 67847 38068 67856
rect 38016 67813 38025 67847
rect 38025 67813 38059 67847
rect 38059 67813 38068 67847
rect 38016 67804 38068 67813
rect 38108 67736 38160 67788
rect 12992 67600 13044 67652
rect 33140 67600 33192 67652
rect 37096 67711 37148 67720
rect 37096 67677 37105 67711
rect 37105 67677 37139 67711
rect 37139 67677 37148 67711
rect 37096 67668 37148 67677
rect 36360 67600 36412 67652
rect 20536 67532 20588 67584
rect 38384 67600 38436 67652
rect 2610 67430 2662 67482
rect 2674 67430 2726 67482
rect 2738 67430 2790 67482
rect 2802 67430 2854 67482
rect 2866 67430 2918 67482
rect 7610 67430 7662 67482
rect 7674 67430 7726 67482
rect 7738 67430 7790 67482
rect 7802 67430 7854 67482
rect 7866 67430 7918 67482
rect 12610 67430 12662 67482
rect 12674 67430 12726 67482
rect 12738 67430 12790 67482
rect 12802 67430 12854 67482
rect 12866 67430 12918 67482
rect 17610 67430 17662 67482
rect 17674 67430 17726 67482
rect 17738 67430 17790 67482
rect 17802 67430 17854 67482
rect 17866 67430 17918 67482
rect 22610 67430 22662 67482
rect 22674 67430 22726 67482
rect 22738 67430 22790 67482
rect 22802 67430 22854 67482
rect 22866 67430 22918 67482
rect 27610 67430 27662 67482
rect 27674 67430 27726 67482
rect 27738 67430 27790 67482
rect 27802 67430 27854 67482
rect 27866 67430 27918 67482
rect 32610 67430 32662 67482
rect 32674 67430 32726 67482
rect 32738 67430 32790 67482
rect 32802 67430 32854 67482
rect 32866 67430 32918 67482
rect 37610 67430 37662 67482
rect 37674 67430 37726 67482
rect 37738 67430 37790 67482
rect 37802 67430 37854 67482
rect 37866 67430 37918 67482
rect 18144 67260 18196 67312
rect 37280 67260 37332 67312
rect 38844 67260 38896 67312
rect 10508 67099 10560 67108
rect 10508 67065 10517 67099
rect 10517 67065 10551 67099
rect 10551 67065 10560 67099
rect 10508 67056 10560 67065
rect 13176 67192 13228 67244
rect 18604 67235 18656 67244
rect 18604 67201 18613 67235
rect 18613 67201 18647 67235
rect 18647 67201 18656 67235
rect 18604 67192 18656 67201
rect 23296 67192 23348 67244
rect 24124 67192 24176 67244
rect 18236 67124 18288 67176
rect 18328 67056 18380 67108
rect 38016 67235 38068 67244
rect 38016 67201 38025 67235
rect 38025 67201 38059 67235
rect 38059 67201 38068 67235
rect 38016 67192 38068 67201
rect 38292 67235 38344 67244
rect 38292 67201 38301 67235
rect 38301 67201 38335 67235
rect 38335 67201 38344 67235
rect 38292 67192 38344 67201
rect 40500 67235 40552 67244
rect 40500 67201 40509 67235
rect 40509 67201 40543 67235
rect 40543 67201 40552 67235
rect 40500 67192 40552 67201
rect 38292 67056 38344 67108
rect 20076 66988 20128 67040
rect 1950 66886 2002 66938
rect 2014 66886 2066 66938
rect 2078 66886 2130 66938
rect 2142 66886 2194 66938
rect 2206 66886 2258 66938
rect 6950 66886 7002 66938
rect 7014 66886 7066 66938
rect 7078 66886 7130 66938
rect 7142 66886 7194 66938
rect 7206 66886 7258 66938
rect 11950 66886 12002 66938
rect 12014 66886 12066 66938
rect 12078 66886 12130 66938
rect 12142 66886 12194 66938
rect 12206 66886 12258 66938
rect 16950 66886 17002 66938
rect 17014 66886 17066 66938
rect 17078 66886 17130 66938
rect 17142 66886 17194 66938
rect 17206 66886 17258 66938
rect 21950 66886 22002 66938
rect 22014 66886 22066 66938
rect 22078 66886 22130 66938
rect 22142 66886 22194 66938
rect 22206 66886 22258 66938
rect 26950 66886 27002 66938
rect 27014 66886 27066 66938
rect 27078 66886 27130 66938
rect 27142 66886 27194 66938
rect 27206 66886 27258 66938
rect 31950 66886 32002 66938
rect 32014 66886 32066 66938
rect 32078 66886 32130 66938
rect 32142 66886 32194 66938
rect 32206 66886 32258 66938
rect 36950 66886 37002 66938
rect 37014 66886 37066 66938
rect 37078 66886 37130 66938
rect 37142 66886 37194 66938
rect 37206 66886 37258 66938
rect 8116 66759 8168 66768
rect 8116 66725 8125 66759
rect 8125 66725 8159 66759
rect 8159 66725 8168 66759
rect 8116 66716 8168 66725
rect 7472 66623 7524 66632
rect 7472 66589 7481 66623
rect 7481 66589 7515 66623
rect 7515 66589 7524 66623
rect 7472 66580 7524 66589
rect 10416 66580 10468 66632
rect 26148 66623 26200 66632
rect 26148 66589 26157 66623
rect 26157 66589 26191 66623
rect 26191 66589 26200 66623
rect 26148 66580 26200 66589
rect 26332 66623 26384 66632
rect 26332 66589 26341 66623
rect 26341 66589 26375 66623
rect 26375 66589 26384 66623
rect 26332 66580 26384 66589
rect 26424 66623 26476 66632
rect 26424 66589 26433 66623
rect 26433 66589 26467 66623
rect 26467 66589 26476 66623
rect 26424 66580 26476 66589
rect 18972 66512 19024 66564
rect 29644 66623 29696 66632
rect 29644 66589 29653 66623
rect 29653 66589 29687 66623
rect 29687 66589 29696 66623
rect 29644 66580 29696 66589
rect 30104 66623 30156 66632
rect 30104 66589 30113 66623
rect 30113 66589 30147 66623
rect 30147 66589 30156 66623
rect 30104 66580 30156 66589
rect 30288 66580 30340 66632
rect 34704 66512 34756 66564
rect 20628 66444 20680 66496
rect 29368 66444 29420 66496
rect 2610 66342 2662 66394
rect 2674 66342 2726 66394
rect 2738 66342 2790 66394
rect 2802 66342 2854 66394
rect 2866 66342 2918 66394
rect 7610 66342 7662 66394
rect 7674 66342 7726 66394
rect 7738 66342 7790 66394
rect 7802 66342 7854 66394
rect 7866 66342 7918 66394
rect 12610 66342 12662 66394
rect 12674 66342 12726 66394
rect 12738 66342 12790 66394
rect 12802 66342 12854 66394
rect 12866 66342 12918 66394
rect 17610 66342 17662 66394
rect 17674 66342 17726 66394
rect 17738 66342 17790 66394
rect 17802 66342 17854 66394
rect 17866 66342 17918 66394
rect 22610 66342 22662 66394
rect 22674 66342 22726 66394
rect 22738 66342 22790 66394
rect 22802 66342 22854 66394
rect 22866 66342 22918 66394
rect 27610 66342 27662 66394
rect 27674 66342 27726 66394
rect 27738 66342 27790 66394
rect 27802 66342 27854 66394
rect 27866 66342 27918 66394
rect 32610 66342 32662 66394
rect 32674 66342 32726 66394
rect 32738 66342 32790 66394
rect 32802 66342 32854 66394
rect 32866 66342 32918 66394
rect 37610 66342 37662 66394
rect 37674 66342 37726 66394
rect 37738 66342 37790 66394
rect 37802 66342 37854 66394
rect 37866 66342 37918 66394
rect 4528 66147 4580 66156
rect 4528 66113 4537 66147
rect 4537 66113 4571 66147
rect 4571 66113 4580 66147
rect 4528 66104 4580 66113
rect 6460 66104 6512 66156
rect 23388 66104 23440 66156
rect 39580 66172 39632 66224
rect 13176 66036 13228 66088
rect 31024 66036 31076 66088
rect 35992 66036 36044 66088
rect 4988 65968 5040 66020
rect 18880 65968 18932 66020
rect 26424 65968 26476 66020
rect 24676 65900 24728 65952
rect 1950 65798 2002 65850
rect 2014 65798 2066 65850
rect 2078 65798 2130 65850
rect 2142 65798 2194 65850
rect 2206 65798 2258 65850
rect 6950 65798 7002 65850
rect 7014 65798 7066 65850
rect 7078 65798 7130 65850
rect 7142 65798 7194 65850
rect 7206 65798 7258 65850
rect 11950 65798 12002 65850
rect 12014 65798 12066 65850
rect 12078 65798 12130 65850
rect 12142 65798 12194 65850
rect 12206 65798 12258 65850
rect 16950 65798 17002 65850
rect 17014 65798 17066 65850
rect 17078 65798 17130 65850
rect 17142 65798 17194 65850
rect 17206 65798 17258 65850
rect 21950 65798 22002 65850
rect 22014 65798 22066 65850
rect 22078 65798 22130 65850
rect 22142 65798 22194 65850
rect 22206 65798 22258 65850
rect 26950 65798 27002 65850
rect 27014 65798 27066 65850
rect 27078 65798 27130 65850
rect 27142 65798 27194 65850
rect 27206 65798 27258 65850
rect 31950 65798 32002 65850
rect 32014 65798 32066 65850
rect 32078 65798 32130 65850
rect 32142 65798 32194 65850
rect 32206 65798 32258 65850
rect 36950 65798 37002 65850
rect 37014 65798 37066 65850
rect 37078 65798 37130 65850
rect 37142 65798 37194 65850
rect 37206 65798 37258 65850
rect 14556 65696 14608 65748
rect 26332 65696 26384 65748
rect 30564 65696 30616 65748
rect 33140 65696 33192 65748
rect 2964 65560 3016 65612
rect 1584 65424 1636 65476
rect 13084 65628 13136 65680
rect 25504 65628 25556 65680
rect 25596 65628 25648 65680
rect 30104 65628 30156 65680
rect 6368 65560 6420 65612
rect 20536 65560 20588 65612
rect 21732 65560 21784 65612
rect 37280 65560 37332 65612
rect 9588 65492 9640 65544
rect 11888 65535 11940 65544
rect 11888 65501 11897 65535
rect 11897 65501 11931 65535
rect 11931 65501 11940 65535
rect 11888 65492 11940 65501
rect 12348 65424 12400 65476
rect 30472 65424 30524 65476
rect 19616 65356 19668 65408
rect 2610 65254 2662 65306
rect 2674 65254 2726 65306
rect 2738 65254 2790 65306
rect 2802 65254 2854 65306
rect 2866 65254 2918 65306
rect 7610 65254 7662 65306
rect 7674 65254 7726 65306
rect 7738 65254 7790 65306
rect 7802 65254 7854 65306
rect 7866 65254 7918 65306
rect 12610 65254 12662 65306
rect 12674 65254 12726 65306
rect 12738 65254 12790 65306
rect 12802 65254 12854 65306
rect 12866 65254 12918 65306
rect 17610 65254 17662 65306
rect 17674 65254 17726 65306
rect 17738 65254 17790 65306
rect 17802 65254 17854 65306
rect 17866 65254 17918 65306
rect 22610 65254 22662 65306
rect 22674 65254 22726 65306
rect 22738 65254 22790 65306
rect 22802 65254 22854 65306
rect 22866 65254 22918 65306
rect 27610 65254 27662 65306
rect 27674 65254 27726 65306
rect 27738 65254 27790 65306
rect 27802 65254 27854 65306
rect 27866 65254 27918 65306
rect 32610 65254 32662 65306
rect 32674 65254 32726 65306
rect 32738 65254 32790 65306
rect 32802 65254 32854 65306
rect 32866 65254 32918 65306
rect 37610 65254 37662 65306
rect 37674 65254 37726 65306
rect 37738 65254 37790 65306
rect 37802 65254 37854 65306
rect 37866 65254 37918 65306
rect 11888 65152 11940 65204
rect 16396 65152 16448 65204
rect 7840 64812 7892 64864
rect 31116 64812 31168 64864
rect 1950 64710 2002 64762
rect 2014 64710 2066 64762
rect 2078 64710 2130 64762
rect 2142 64710 2194 64762
rect 2206 64710 2258 64762
rect 6950 64710 7002 64762
rect 7014 64710 7066 64762
rect 7078 64710 7130 64762
rect 7142 64710 7194 64762
rect 7206 64710 7258 64762
rect 11950 64710 12002 64762
rect 12014 64710 12066 64762
rect 12078 64710 12130 64762
rect 12142 64710 12194 64762
rect 12206 64710 12258 64762
rect 16950 64710 17002 64762
rect 17014 64710 17066 64762
rect 17078 64710 17130 64762
rect 17142 64710 17194 64762
rect 17206 64710 17258 64762
rect 21950 64710 22002 64762
rect 22014 64710 22066 64762
rect 22078 64710 22130 64762
rect 22142 64710 22194 64762
rect 22206 64710 22258 64762
rect 26950 64710 27002 64762
rect 27014 64710 27066 64762
rect 27078 64710 27130 64762
rect 27142 64710 27194 64762
rect 27206 64710 27258 64762
rect 31950 64710 32002 64762
rect 32014 64710 32066 64762
rect 32078 64710 32130 64762
rect 32142 64710 32194 64762
rect 32206 64710 32258 64762
rect 36950 64710 37002 64762
rect 37014 64710 37066 64762
rect 37078 64710 37130 64762
rect 37142 64710 37194 64762
rect 37206 64710 37258 64762
rect 14004 64608 14056 64660
rect 20628 64608 20680 64660
rect 20812 64651 20864 64660
rect 20812 64617 20821 64651
rect 20821 64617 20855 64651
rect 20855 64617 20864 64651
rect 20812 64608 20864 64617
rect 8116 64540 8168 64592
rect 13452 64472 13504 64524
rect 32404 64540 32456 64592
rect 20168 64515 20220 64524
rect 20168 64481 20177 64515
rect 20177 64481 20211 64515
rect 20211 64481 20220 64515
rect 20168 64472 20220 64481
rect 7840 64447 7892 64456
rect 7840 64413 7849 64447
rect 7849 64413 7883 64447
rect 7883 64413 7892 64447
rect 7840 64404 7892 64413
rect 13544 64404 13596 64456
rect 19248 64404 19300 64456
rect 31484 64472 31536 64524
rect 20352 64447 20404 64456
rect 20352 64413 20361 64447
rect 20361 64413 20395 64447
rect 20395 64413 20404 64447
rect 20352 64404 20404 64413
rect 17316 64336 17368 64388
rect 20720 64447 20772 64456
rect 20720 64413 20729 64447
rect 20729 64413 20763 64447
rect 20763 64413 20772 64447
rect 20720 64404 20772 64413
rect 21088 64447 21140 64456
rect 21088 64413 21097 64447
rect 21097 64413 21131 64447
rect 21131 64413 21140 64447
rect 21088 64404 21140 64413
rect 21732 64447 21784 64456
rect 21732 64413 21741 64447
rect 21741 64413 21775 64447
rect 21775 64413 21784 64447
rect 21732 64404 21784 64413
rect 33692 64447 33744 64456
rect 33692 64413 33701 64447
rect 33701 64413 33735 64447
rect 33735 64413 33744 64447
rect 33692 64404 33744 64413
rect 36728 64404 36780 64456
rect 33600 64379 33652 64388
rect 33600 64345 33609 64379
rect 33609 64345 33643 64379
rect 33643 64345 33652 64379
rect 33600 64336 33652 64345
rect 20260 64268 20312 64320
rect 24400 64268 24452 64320
rect 2610 64166 2662 64218
rect 2674 64166 2726 64218
rect 2738 64166 2790 64218
rect 2802 64166 2854 64218
rect 2866 64166 2918 64218
rect 7610 64166 7662 64218
rect 7674 64166 7726 64218
rect 7738 64166 7790 64218
rect 7802 64166 7854 64218
rect 7866 64166 7918 64218
rect 12610 64166 12662 64218
rect 12674 64166 12726 64218
rect 12738 64166 12790 64218
rect 12802 64166 12854 64218
rect 12866 64166 12918 64218
rect 17610 64166 17662 64218
rect 17674 64166 17726 64218
rect 17738 64166 17790 64218
rect 17802 64166 17854 64218
rect 17866 64166 17918 64218
rect 22610 64166 22662 64218
rect 22674 64166 22726 64218
rect 22738 64166 22790 64218
rect 22802 64166 22854 64218
rect 22866 64166 22918 64218
rect 27610 64166 27662 64218
rect 27674 64166 27726 64218
rect 27738 64166 27790 64218
rect 27802 64166 27854 64218
rect 27866 64166 27918 64218
rect 32610 64166 32662 64218
rect 32674 64166 32726 64218
rect 32738 64166 32790 64218
rect 32802 64166 32854 64218
rect 32866 64166 32918 64218
rect 37610 64166 37662 64218
rect 37674 64166 37726 64218
rect 37738 64166 37790 64218
rect 37802 64166 37854 64218
rect 37866 64166 37918 64218
rect 15108 63996 15160 64048
rect 20720 63996 20772 64048
rect 35256 63996 35308 64048
rect 36360 63928 36412 63980
rect 38108 63971 38160 63980
rect 38108 63937 38117 63971
rect 38117 63937 38151 63971
rect 38151 63937 38160 63971
rect 38108 63928 38160 63937
rect 30196 63792 30248 63844
rect 37372 63860 37424 63912
rect 1950 63622 2002 63674
rect 2014 63622 2066 63674
rect 2078 63622 2130 63674
rect 2142 63622 2194 63674
rect 2206 63622 2258 63674
rect 6950 63622 7002 63674
rect 7014 63622 7066 63674
rect 7078 63622 7130 63674
rect 7142 63622 7194 63674
rect 7206 63622 7258 63674
rect 11950 63622 12002 63674
rect 12014 63622 12066 63674
rect 12078 63622 12130 63674
rect 12142 63622 12194 63674
rect 12206 63622 12258 63674
rect 16950 63622 17002 63674
rect 17014 63622 17066 63674
rect 17078 63622 17130 63674
rect 17142 63622 17194 63674
rect 17206 63622 17258 63674
rect 21950 63622 22002 63674
rect 22014 63622 22066 63674
rect 22078 63622 22130 63674
rect 22142 63622 22194 63674
rect 22206 63622 22258 63674
rect 26950 63622 27002 63674
rect 27014 63622 27066 63674
rect 27078 63622 27130 63674
rect 27142 63622 27194 63674
rect 27206 63622 27258 63674
rect 31950 63622 32002 63674
rect 32014 63622 32066 63674
rect 32078 63622 32130 63674
rect 32142 63622 32194 63674
rect 32206 63622 32258 63674
rect 36950 63622 37002 63674
rect 37014 63622 37066 63674
rect 37078 63622 37130 63674
rect 37142 63622 37194 63674
rect 37206 63622 37258 63674
rect 16396 63520 16448 63572
rect 34796 63520 34848 63572
rect 35256 63520 35308 63572
rect 22376 63384 22428 63436
rect 26700 63291 26752 63300
rect 26700 63257 26709 63291
rect 26709 63257 26743 63291
rect 26743 63257 26752 63291
rect 29736 63316 29788 63368
rect 26700 63248 26752 63257
rect 35440 63248 35492 63300
rect 17960 63180 18012 63232
rect 27988 63180 28040 63232
rect 2610 63078 2662 63130
rect 2674 63078 2726 63130
rect 2738 63078 2790 63130
rect 2802 63078 2854 63130
rect 2866 63078 2918 63130
rect 7610 63078 7662 63130
rect 7674 63078 7726 63130
rect 7738 63078 7790 63130
rect 7802 63078 7854 63130
rect 7866 63078 7918 63130
rect 12610 63078 12662 63130
rect 12674 63078 12726 63130
rect 12738 63078 12790 63130
rect 12802 63078 12854 63130
rect 12866 63078 12918 63130
rect 17610 63078 17662 63130
rect 17674 63078 17726 63130
rect 17738 63078 17790 63130
rect 17802 63078 17854 63130
rect 17866 63078 17918 63130
rect 22610 63078 22662 63130
rect 22674 63078 22726 63130
rect 22738 63078 22790 63130
rect 22802 63078 22854 63130
rect 22866 63078 22918 63130
rect 27610 63078 27662 63130
rect 27674 63078 27726 63130
rect 27738 63078 27790 63130
rect 27802 63078 27854 63130
rect 27866 63078 27918 63130
rect 32610 63078 32662 63130
rect 32674 63078 32726 63130
rect 32738 63078 32790 63130
rect 32802 63078 32854 63130
rect 32866 63078 32918 63130
rect 37610 63078 37662 63130
rect 37674 63078 37726 63130
rect 37738 63078 37790 63130
rect 37802 63078 37854 63130
rect 37866 63078 37918 63130
rect 16304 62976 16356 63028
rect 14648 62908 14700 62960
rect 30288 62908 30340 62960
rect 6828 62840 6880 62892
rect 10876 62840 10928 62892
rect 19984 62840 20036 62892
rect 1860 62772 1912 62824
rect 8944 62772 8996 62824
rect 16580 62772 16632 62824
rect 4896 62704 4948 62756
rect 9588 62636 9640 62688
rect 13360 62704 13412 62756
rect 25044 62704 25096 62756
rect 17960 62636 18012 62688
rect 1950 62534 2002 62586
rect 2014 62534 2066 62586
rect 2078 62534 2130 62586
rect 2142 62534 2194 62586
rect 2206 62534 2258 62586
rect 6950 62534 7002 62586
rect 7014 62534 7066 62586
rect 7078 62534 7130 62586
rect 7142 62534 7194 62586
rect 7206 62534 7258 62586
rect 11950 62534 12002 62586
rect 12014 62534 12066 62586
rect 12078 62534 12130 62586
rect 12142 62534 12194 62586
rect 12206 62534 12258 62586
rect 16950 62534 17002 62586
rect 17014 62534 17066 62586
rect 17078 62534 17130 62586
rect 17142 62534 17194 62586
rect 17206 62534 17258 62586
rect 21950 62534 22002 62586
rect 22014 62534 22066 62586
rect 22078 62534 22130 62586
rect 22142 62534 22194 62586
rect 22206 62534 22258 62586
rect 26950 62534 27002 62586
rect 27014 62534 27066 62586
rect 27078 62534 27130 62586
rect 27142 62534 27194 62586
rect 27206 62534 27258 62586
rect 31950 62534 32002 62586
rect 32014 62534 32066 62586
rect 32078 62534 32130 62586
rect 32142 62534 32194 62586
rect 32206 62534 32258 62586
rect 36950 62534 37002 62586
rect 37014 62534 37066 62586
rect 37078 62534 37130 62586
rect 37142 62534 37194 62586
rect 37206 62534 37258 62586
rect 12900 62432 12952 62484
rect 27436 62432 27488 62484
rect 7380 62271 7432 62280
rect 7380 62237 7389 62271
rect 7389 62237 7423 62271
rect 7423 62237 7432 62271
rect 7380 62228 7432 62237
rect 15108 62296 15160 62348
rect 4436 62092 4488 62144
rect 12532 62271 12584 62280
rect 12532 62237 12541 62271
rect 12541 62237 12575 62271
rect 12575 62237 12584 62271
rect 12532 62228 12584 62237
rect 12900 62271 12952 62280
rect 12900 62237 12909 62271
rect 12909 62237 12943 62271
rect 12943 62237 12952 62271
rect 12900 62228 12952 62237
rect 13360 62271 13412 62280
rect 13360 62237 13369 62271
rect 13369 62237 13403 62271
rect 13403 62237 13412 62271
rect 13360 62228 13412 62237
rect 13268 62092 13320 62144
rect 13912 62092 13964 62144
rect 17960 62092 18012 62144
rect 18144 62364 18196 62416
rect 29000 62364 29052 62416
rect 30196 62364 30248 62416
rect 18236 62296 18288 62348
rect 30288 62296 30340 62348
rect 28264 62228 28316 62280
rect 30656 62228 30708 62280
rect 35256 62271 35308 62280
rect 35256 62237 35265 62271
rect 35265 62237 35299 62271
rect 35299 62237 35308 62271
rect 35256 62228 35308 62237
rect 35624 62271 35676 62280
rect 35624 62237 35633 62271
rect 35633 62237 35667 62271
rect 35667 62237 35676 62271
rect 35624 62228 35676 62237
rect 20076 62160 20128 62212
rect 20352 62203 20404 62212
rect 20352 62169 20361 62203
rect 20361 62169 20395 62203
rect 20395 62169 20404 62203
rect 20352 62160 20404 62169
rect 20904 62203 20956 62212
rect 20904 62169 20913 62203
rect 20913 62169 20947 62203
rect 20947 62169 20956 62203
rect 20904 62160 20956 62169
rect 23204 62092 23256 62144
rect 23388 62092 23440 62144
rect 2610 61990 2662 62042
rect 2674 61990 2726 62042
rect 2738 61990 2790 62042
rect 2802 61990 2854 62042
rect 2866 61990 2918 62042
rect 7610 61990 7662 62042
rect 7674 61990 7726 62042
rect 7738 61990 7790 62042
rect 7802 61990 7854 62042
rect 7866 61990 7918 62042
rect 12610 61990 12662 62042
rect 12674 61990 12726 62042
rect 12738 61990 12790 62042
rect 12802 61990 12854 62042
rect 12866 61990 12918 62042
rect 17610 61990 17662 62042
rect 17674 61990 17726 62042
rect 17738 61990 17790 62042
rect 17802 61990 17854 62042
rect 17866 61990 17918 62042
rect 22610 61990 22662 62042
rect 22674 61990 22726 62042
rect 22738 61990 22790 62042
rect 22802 61990 22854 62042
rect 22866 61990 22918 62042
rect 27610 61990 27662 62042
rect 27674 61990 27726 62042
rect 27738 61990 27790 62042
rect 27802 61990 27854 62042
rect 27866 61990 27918 62042
rect 32610 61990 32662 62042
rect 32674 61990 32726 62042
rect 32738 61990 32790 62042
rect 32802 61990 32854 62042
rect 32866 61990 32918 62042
rect 37610 61990 37662 62042
rect 37674 61990 37726 62042
rect 37738 61990 37790 62042
rect 37802 61990 37854 62042
rect 37866 61990 37918 62042
rect 13820 61752 13872 61804
rect 11796 61684 11848 61736
rect 13728 61727 13780 61736
rect 13728 61693 13737 61727
rect 13737 61693 13771 61727
rect 13771 61693 13780 61727
rect 13728 61684 13780 61693
rect 17960 61548 18012 61600
rect 18788 61548 18840 61600
rect 1950 61446 2002 61498
rect 2014 61446 2066 61498
rect 2078 61446 2130 61498
rect 2142 61446 2194 61498
rect 2206 61446 2258 61498
rect 6950 61446 7002 61498
rect 7014 61446 7066 61498
rect 7078 61446 7130 61498
rect 7142 61446 7194 61498
rect 7206 61446 7258 61498
rect 11950 61446 12002 61498
rect 12014 61446 12066 61498
rect 12078 61446 12130 61498
rect 12142 61446 12194 61498
rect 12206 61446 12258 61498
rect 16950 61446 17002 61498
rect 17014 61446 17066 61498
rect 17078 61446 17130 61498
rect 17142 61446 17194 61498
rect 17206 61446 17258 61498
rect 21950 61446 22002 61498
rect 22014 61446 22066 61498
rect 22078 61446 22130 61498
rect 22142 61446 22194 61498
rect 22206 61446 22258 61498
rect 26950 61446 27002 61498
rect 27014 61446 27066 61498
rect 27078 61446 27130 61498
rect 27142 61446 27194 61498
rect 27206 61446 27258 61498
rect 31950 61446 32002 61498
rect 32014 61446 32066 61498
rect 32078 61446 32130 61498
rect 32142 61446 32194 61498
rect 32206 61446 32258 61498
rect 36950 61446 37002 61498
rect 37014 61446 37066 61498
rect 37078 61446 37130 61498
rect 37142 61446 37194 61498
rect 37206 61446 37258 61498
rect 13912 61344 13964 61396
rect 36544 61344 36596 61396
rect 2504 61140 2556 61192
rect 5540 61140 5592 61192
rect 8944 61183 8996 61192
rect 8944 61149 8953 61183
rect 8953 61149 8987 61183
rect 8987 61149 8996 61183
rect 8944 61140 8996 61149
rect 9220 61183 9272 61192
rect 9220 61149 9229 61183
rect 9229 61149 9263 61183
rect 9263 61149 9272 61183
rect 9220 61140 9272 61149
rect 17960 61208 18012 61260
rect 19248 61208 19300 61260
rect 33876 61140 33928 61192
rect 2320 61115 2372 61124
rect 2320 61081 2329 61115
rect 2329 61081 2363 61115
rect 2363 61081 2372 61115
rect 2320 61072 2372 61081
rect 3700 61072 3752 61124
rect 3884 61047 3936 61056
rect 3884 61013 3893 61047
rect 3893 61013 3927 61047
rect 3927 61013 3936 61047
rect 3884 61004 3936 61013
rect 4712 61072 4764 61124
rect 8024 61072 8076 61124
rect 10324 61072 10376 61124
rect 4804 61047 4856 61056
rect 4804 61013 4813 61047
rect 4813 61013 4847 61047
rect 4847 61013 4856 61047
rect 4804 61004 4856 61013
rect 2610 60902 2662 60954
rect 2674 60902 2726 60954
rect 2738 60902 2790 60954
rect 2802 60902 2854 60954
rect 2866 60902 2918 60954
rect 7610 60902 7662 60954
rect 7674 60902 7726 60954
rect 7738 60902 7790 60954
rect 7802 60902 7854 60954
rect 7866 60902 7918 60954
rect 12610 60902 12662 60954
rect 12674 60902 12726 60954
rect 12738 60902 12790 60954
rect 12802 60902 12854 60954
rect 12866 60902 12918 60954
rect 17610 60902 17662 60954
rect 17674 60902 17726 60954
rect 17738 60902 17790 60954
rect 17802 60902 17854 60954
rect 17866 60902 17918 60954
rect 22610 60902 22662 60954
rect 22674 60902 22726 60954
rect 22738 60902 22790 60954
rect 22802 60902 22854 60954
rect 22866 60902 22918 60954
rect 27610 60902 27662 60954
rect 27674 60902 27726 60954
rect 27738 60902 27790 60954
rect 27802 60902 27854 60954
rect 27866 60902 27918 60954
rect 32610 60902 32662 60954
rect 32674 60902 32726 60954
rect 32738 60902 32790 60954
rect 32802 60902 32854 60954
rect 32866 60902 32918 60954
rect 37610 60902 37662 60954
rect 37674 60902 37726 60954
rect 37738 60902 37790 60954
rect 37802 60902 37854 60954
rect 37866 60902 37918 60954
rect 4804 60732 4856 60784
rect 10692 60732 10744 60784
rect 1676 60664 1728 60716
rect 8484 60707 8536 60716
rect 8484 60673 8493 60707
rect 8493 60673 8527 60707
rect 8527 60673 8536 60707
rect 8484 60664 8536 60673
rect 5540 60596 5592 60648
rect 9036 60664 9088 60716
rect 18604 60664 18656 60716
rect 29552 60707 29604 60716
rect 29552 60673 29561 60707
rect 29561 60673 29595 60707
rect 29595 60673 29604 60707
rect 29552 60664 29604 60673
rect 38660 60707 38712 60716
rect 38660 60673 38669 60707
rect 38669 60673 38703 60707
rect 38703 60673 38712 60707
rect 38660 60664 38712 60673
rect 38752 60707 38804 60716
rect 38752 60673 38761 60707
rect 38761 60673 38795 60707
rect 38795 60673 38804 60707
rect 38752 60664 38804 60673
rect 38844 60596 38896 60648
rect 5540 60460 5592 60512
rect 8116 60460 8168 60512
rect 8852 60503 8904 60512
rect 8852 60469 8861 60503
rect 8861 60469 8895 60503
rect 8895 60469 8904 60503
rect 8852 60460 8904 60469
rect 19708 60460 19760 60512
rect 29092 60503 29144 60512
rect 29092 60469 29101 60503
rect 29101 60469 29135 60503
rect 29135 60469 29144 60503
rect 29092 60460 29144 60469
rect 39120 60503 39172 60512
rect 39120 60469 39129 60503
rect 39129 60469 39163 60503
rect 39163 60469 39172 60503
rect 39120 60460 39172 60469
rect 1950 60358 2002 60410
rect 2014 60358 2066 60410
rect 2078 60358 2130 60410
rect 2142 60358 2194 60410
rect 2206 60358 2258 60410
rect 6950 60358 7002 60410
rect 7014 60358 7066 60410
rect 7078 60358 7130 60410
rect 7142 60358 7194 60410
rect 7206 60358 7258 60410
rect 11950 60358 12002 60410
rect 12014 60358 12066 60410
rect 12078 60358 12130 60410
rect 12142 60358 12194 60410
rect 12206 60358 12258 60410
rect 16950 60358 17002 60410
rect 17014 60358 17066 60410
rect 17078 60358 17130 60410
rect 17142 60358 17194 60410
rect 17206 60358 17258 60410
rect 21950 60358 22002 60410
rect 22014 60358 22066 60410
rect 22078 60358 22130 60410
rect 22142 60358 22194 60410
rect 22206 60358 22258 60410
rect 26950 60358 27002 60410
rect 27014 60358 27066 60410
rect 27078 60358 27130 60410
rect 27142 60358 27194 60410
rect 27206 60358 27258 60410
rect 31950 60358 32002 60410
rect 32014 60358 32066 60410
rect 32078 60358 32130 60410
rect 32142 60358 32194 60410
rect 32206 60358 32258 60410
rect 36950 60358 37002 60410
rect 37014 60358 37066 60410
rect 37078 60358 37130 60410
rect 37142 60358 37194 60410
rect 37206 60358 37258 60410
rect 19616 60299 19668 60308
rect 19616 60265 19625 60299
rect 19625 60265 19659 60299
rect 19659 60265 19668 60299
rect 19616 60256 19668 60265
rect 34704 60299 34756 60308
rect 34704 60265 34713 60299
rect 34713 60265 34747 60299
rect 34747 60265 34756 60299
rect 34704 60256 34756 60265
rect 6000 60052 6052 60104
rect 19248 60095 19300 60104
rect 19248 60061 19257 60095
rect 19257 60061 19291 60095
rect 19291 60061 19300 60095
rect 19248 60052 19300 60061
rect 23848 60120 23900 60172
rect 29644 60163 29696 60172
rect 29644 60129 29653 60163
rect 29653 60129 29687 60163
rect 29687 60129 29696 60163
rect 29644 60120 29696 60129
rect 22100 60095 22152 60104
rect 22100 60061 22109 60095
rect 22109 60061 22143 60095
rect 22143 60061 22152 60095
rect 22100 60052 22152 60061
rect 23112 60052 23164 60104
rect 28908 60052 28960 60104
rect 21272 60027 21324 60036
rect 21272 59993 21281 60027
rect 21281 59993 21315 60027
rect 21315 59993 21324 60027
rect 21272 59984 21324 59993
rect 30932 60052 30984 60104
rect 33140 60095 33192 60104
rect 33140 60061 33149 60095
rect 33149 60061 33183 60095
rect 33183 60061 33192 60095
rect 33140 60052 33192 60061
rect 33416 60095 33468 60104
rect 33416 60061 33425 60095
rect 33425 60061 33459 60095
rect 33459 60061 33468 60095
rect 33416 60052 33468 60061
rect 33784 60095 33836 60104
rect 33784 60061 33793 60095
rect 33793 60061 33827 60095
rect 33827 60061 33836 60095
rect 33784 60052 33836 60061
rect 34152 60095 34204 60104
rect 34152 60061 34161 60095
rect 34161 60061 34195 60095
rect 34195 60061 34204 60095
rect 34152 60052 34204 60061
rect 34704 60027 34756 60036
rect 34704 59993 34713 60027
rect 34713 59993 34747 60027
rect 34747 59993 34756 60027
rect 34704 59984 34756 59993
rect 39120 60256 39172 60308
rect 19708 59916 19760 59968
rect 22468 59916 22520 59968
rect 27528 59916 27580 59968
rect 34888 59959 34940 59968
rect 34888 59925 34897 59959
rect 34897 59925 34931 59959
rect 34931 59925 34940 59959
rect 34888 59916 34940 59925
rect 2610 59814 2662 59866
rect 2674 59814 2726 59866
rect 2738 59814 2790 59866
rect 2802 59814 2854 59866
rect 2866 59814 2918 59866
rect 7610 59814 7662 59866
rect 7674 59814 7726 59866
rect 7738 59814 7790 59866
rect 7802 59814 7854 59866
rect 7866 59814 7918 59866
rect 12610 59814 12662 59866
rect 12674 59814 12726 59866
rect 12738 59814 12790 59866
rect 12802 59814 12854 59866
rect 12866 59814 12918 59866
rect 17610 59814 17662 59866
rect 17674 59814 17726 59866
rect 17738 59814 17790 59866
rect 17802 59814 17854 59866
rect 17866 59814 17918 59866
rect 22610 59814 22662 59866
rect 22674 59814 22726 59866
rect 22738 59814 22790 59866
rect 22802 59814 22854 59866
rect 22866 59814 22918 59866
rect 27610 59814 27662 59866
rect 27674 59814 27726 59866
rect 27738 59814 27790 59866
rect 27802 59814 27854 59866
rect 27866 59814 27918 59866
rect 32610 59814 32662 59866
rect 32674 59814 32726 59866
rect 32738 59814 32790 59866
rect 32802 59814 32854 59866
rect 32866 59814 32918 59866
rect 37610 59814 37662 59866
rect 37674 59814 37726 59866
rect 37738 59814 37790 59866
rect 37802 59814 37854 59866
rect 37866 59814 37918 59866
rect 21272 59644 21324 59696
rect 34888 59644 34940 59696
rect 39948 59576 40000 59628
rect 39672 59551 39724 59560
rect 39672 59517 39681 59551
rect 39681 59517 39715 59551
rect 39715 59517 39724 59551
rect 39672 59508 39724 59517
rect 12532 59440 12584 59492
rect 18512 59440 18564 59492
rect 18604 59372 18656 59424
rect 19064 59372 19116 59424
rect 19708 59372 19760 59424
rect 21364 59372 21416 59424
rect 1950 59270 2002 59322
rect 2014 59270 2066 59322
rect 2078 59270 2130 59322
rect 2142 59270 2194 59322
rect 2206 59270 2258 59322
rect 6950 59270 7002 59322
rect 7014 59270 7066 59322
rect 7078 59270 7130 59322
rect 7142 59270 7194 59322
rect 7206 59270 7258 59322
rect 11950 59270 12002 59322
rect 12014 59270 12066 59322
rect 12078 59270 12130 59322
rect 12142 59270 12194 59322
rect 12206 59270 12258 59322
rect 16950 59270 17002 59322
rect 17014 59270 17066 59322
rect 17078 59270 17130 59322
rect 17142 59270 17194 59322
rect 17206 59270 17258 59322
rect 21950 59270 22002 59322
rect 22014 59270 22066 59322
rect 22078 59270 22130 59322
rect 22142 59270 22194 59322
rect 22206 59270 22258 59322
rect 26950 59270 27002 59322
rect 27014 59270 27066 59322
rect 27078 59270 27130 59322
rect 27142 59270 27194 59322
rect 27206 59270 27258 59322
rect 31950 59270 32002 59322
rect 32014 59270 32066 59322
rect 32078 59270 32130 59322
rect 32142 59270 32194 59322
rect 32206 59270 32258 59322
rect 36950 59270 37002 59322
rect 37014 59270 37066 59322
rect 37078 59270 37130 59322
rect 37142 59270 37194 59322
rect 37206 59270 37258 59322
rect 26700 59168 26752 59220
rect 7472 59100 7524 59152
rect 6368 59032 6420 59084
rect 4344 59007 4396 59016
rect 4344 58973 4353 59007
rect 4353 58973 4387 59007
rect 4387 58973 4396 59007
rect 4344 58964 4396 58973
rect 6736 59007 6788 59016
rect 6736 58973 6745 59007
rect 6745 58973 6779 59007
rect 6779 58973 6788 59007
rect 6736 58964 6788 58973
rect 4620 58896 4672 58948
rect 22376 59032 22428 59084
rect 22284 58964 22336 59016
rect 23388 58964 23440 59016
rect 20812 58896 20864 58948
rect 23664 58939 23716 58948
rect 23664 58905 23673 58939
rect 23673 58905 23707 58939
rect 23707 58905 23716 58939
rect 23664 58896 23716 58905
rect 25688 58896 25740 58948
rect 31024 59032 31076 59084
rect 38016 59032 38068 59084
rect 29920 59007 29972 59016
rect 29920 58973 29929 59007
rect 29929 58973 29963 59007
rect 29963 58973 29972 59007
rect 29920 58964 29972 58973
rect 27436 58896 27488 58948
rect 31484 58964 31536 59016
rect 35164 58896 35216 58948
rect 30012 58871 30064 58880
rect 30012 58837 30021 58871
rect 30021 58837 30055 58871
rect 30055 58837 30064 58871
rect 30012 58828 30064 58837
rect 2610 58726 2662 58778
rect 2674 58726 2726 58778
rect 2738 58726 2790 58778
rect 2802 58726 2854 58778
rect 2866 58726 2918 58778
rect 7610 58726 7662 58778
rect 7674 58726 7726 58778
rect 7738 58726 7790 58778
rect 7802 58726 7854 58778
rect 7866 58726 7918 58778
rect 12610 58726 12662 58778
rect 12674 58726 12726 58778
rect 12738 58726 12790 58778
rect 12802 58726 12854 58778
rect 12866 58726 12918 58778
rect 17610 58726 17662 58778
rect 17674 58726 17726 58778
rect 17738 58726 17790 58778
rect 17802 58726 17854 58778
rect 17866 58726 17918 58778
rect 22610 58726 22662 58778
rect 22674 58726 22726 58778
rect 22738 58726 22790 58778
rect 22802 58726 22854 58778
rect 22866 58726 22918 58778
rect 27610 58726 27662 58778
rect 27674 58726 27726 58778
rect 27738 58726 27790 58778
rect 27802 58726 27854 58778
rect 27866 58726 27918 58778
rect 32610 58726 32662 58778
rect 32674 58726 32726 58778
rect 32738 58726 32790 58778
rect 32802 58726 32854 58778
rect 32866 58726 32918 58778
rect 37610 58726 37662 58778
rect 37674 58726 37726 58778
rect 37738 58726 37790 58778
rect 37802 58726 37854 58778
rect 37866 58726 37918 58778
rect 19248 58624 19300 58676
rect 30104 58624 30156 58676
rect 6736 58556 6788 58608
rect 39304 58556 39356 58608
rect 848 58488 900 58540
rect 14372 58531 14424 58540
rect 14372 58497 14381 58531
rect 14381 58497 14415 58531
rect 14415 58497 14424 58531
rect 14372 58488 14424 58497
rect 19892 58488 19944 58540
rect 14004 58463 14056 58472
rect 14004 58429 14013 58463
rect 14013 58429 14047 58463
rect 14047 58429 14056 58463
rect 14004 58420 14056 58429
rect 38016 58420 38068 58472
rect 39120 58488 39172 58540
rect 14188 58352 14240 58404
rect 1950 58182 2002 58234
rect 2014 58182 2066 58234
rect 2078 58182 2130 58234
rect 2142 58182 2194 58234
rect 2206 58182 2258 58234
rect 6950 58182 7002 58234
rect 7014 58182 7066 58234
rect 7078 58182 7130 58234
rect 7142 58182 7194 58234
rect 7206 58182 7258 58234
rect 11950 58182 12002 58234
rect 12014 58182 12066 58234
rect 12078 58182 12130 58234
rect 12142 58182 12194 58234
rect 12206 58182 12258 58234
rect 16950 58182 17002 58234
rect 17014 58182 17066 58234
rect 17078 58182 17130 58234
rect 17142 58182 17194 58234
rect 17206 58182 17258 58234
rect 21950 58182 22002 58234
rect 22014 58182 22066 58234
rect 22078 58182 22130 58234
rect 22142 58182 22194 58234
rect 22206 58182 22258 58234
rect 26950 58182 27002 58234
rect 27014 58182 27066 58234
rect 27078 58182 27130 58234
rect 27142 58182 27194 58234
rect 27206 58182 27258 58234
rect 31950 58182 32002 58234
rect 32014 58182 32066 58234
rect 32078 58182 32130 58234
rect 32142 58182 32194 58234
rect 32206 58182 32258 58234
rect 36950 58182 37002 58234
rect 37014 58182 37066 58234
rect 37078 58182 37130 58234
rect 37142 58182 37194 58234
rect 37206 58182 37258 58234
rect 27528 58123 27580 58132
rect 27528 58089 27537 58123
rect 27537 58089 27571 58123
rect 27571 58089 27580 58123
rect 27528 58080 27580 58089
rect 19892 57987 19944 57996
rect 19892 57953 19901 57987
rect 19901 57953 19935 57987
rect 19935 57953 19944 57987
rect 19892 57944 19944 57953
rect 10968 57876 11020 57928
rect 20076 57919 20128 57928
rect 20076 57885 20085 57919
rect 20085 57885 20119 57919
rect 20119 57885 20128 57919
rect 20076 57876 20128 57885
rect 20720 57876 20772 57928
rect 20996 57919 21048 57928
rect 20996 57885 21005 57919
rect 21005 57885 21039 57919
rect 21039 57885 21048 57919
rect 20996 57876 21048 57885
rect 28080 57876 28132 57928
rect 28908 57808 28960 57860
rect 12440 57740 12492 57792
rect 26148 57740 26200 57792
rect 27528 57783 27580 57792
rect 27528 57749 27546 57783
rect 27546 57749 27580 57783
rect 27528 57740 27580 57749
rect 2610 57638 2662 57690
rect 2674 57638 2726 57690
rect 2738 57638 2790 57690
rect 2802 57638 2854 57690
rect 2866 57638 2918 57690
rect 7610 57638 7662 57690
rect 7674 57638 7726 57690
rect 7738 57638 7790 57690
rect 7802 57638 7854 57690
rect 7866 57638 7918 57690
rect 12610 57638 12662 57690
rect 12674 57638 12726 57690
rect 12738 57638 12790 57690
rect 12802 57638 12854 57690
rect 12866 57638 12918 57690
rect 17610 57638 17662 57690
rect 17674 57638 17726 57690
rect 17738 57638 17790 57690
rect 17802 57638 17854 57690
rect 17866 57638 17918 57690
rect 22610 57638 22662 57690
rect 22674 57638 22726 57690
rect 22738 57638 22790 57690
rect 22802 57638 22854 57690
rect 22866 57638 22918 57690
rect 27610 57638 27662 57690
rect 27674 57638 27726 57690
rect 27738 57638 27790 57690
rect 27802 57638 27854 57690
rect 27866 57638 27918 57690
rect 32610 57638 32662 57690
rect 32674 57638 32726 57690
rect 32738 57638 32790 57690
rect 32802 57638 32854 57690
rect 32866 57638 32918 57690
rect 37610 57638 37662 57690
rect 37674 57638 37726 57690
rect 37738 57638 37790 57690
rect 37802 57638 37854 57690
rect 37866 57638 37918 57690
rect 20720 57536 20772 57588
rect 24860 57536 24912 57588
rect 31668 57536 31720 57588
rect 33416 57536 33468 57588
rect 16856 57400 16908 57452
rect 21548 57400 21600 57452
rect 16672 57375 16724 57384
rect 16672 57341 16681 57375
rect 16681 57341 16715 57375
rect 16715 57341 16724 57375
rect 16672 57332 16724 57341
rect 22376 57332 22428 57384
rect 38936 57400 38988 57452
rect 39212 57400 39264 57452
rect 39580 57443 39632 57452
rect 39580 57409 39589 57443
rect 39589 57409 39623 57443
rect 39623 57409 39632 57443
rect 39580 57400 39632 57409
rect 39856 57443 39908 57452
rect 39856 57409 39865 57443
rect 39865 57409 39899 57443
rect 39899 57409 39908 57443
rect 39856 57400 39908 57409
rect 16120 57264 16172 57316
rect 22284 57264 22336 57316
rect 23664 57264 23716 57316
rect 31208 57264 31260 57316
rect 31300 57264 31352 57316
rect 2320 57196 2372 57248
rect 33508 57196 33560 57248
rect 1950 57094 2002 57146
rect 2014 57094 2066 57146
rect 2078 57094 2130 57146
rect 2142 57094 2194 57146
rect 2206 57094 2258 57146
rect 6950 57094 7002 57146
rect 7014 57094 7066 57146
rect 7078 57094 7130 57146
rect 7142 57094 7194 57146
rect 7206 57094 7258 57146
rect 11950 57094 12002 57146
rect 12014 57094 12066 57146
rect 12078 57094 12130 57146
rect 12142 57094 12194 57146
rect 12206 57094 12258 57146
rect 16950 57094 17002 57146
rect 17014 57094 17066 57146
rect 17078 57094 17130 57146
rect 17142 57094 17194 57146
rect 17206 57094 17258 57146
rect 21950 57094 22002 57146
rect 22014 57094 22066 57146
rect 22078 57094 22130 57146
rect 22142 57094 22194 57146
rect 22206 57094 22258 57146
rect 26950 57094 27002 57146
rect 27014 57094 27066 57146
rect 27078 57094 27130 57146
rect 27142 57094 27194 57146
rect 27206 57094 27258 57146
rect 31950 57094 32002 57146
rect 32014 57094 32066 57146
rect 32078 57094 32130 57146
rect 32142 57094 32194 57146
rect 32206 57094 32258 57146
rect 36950 57094 37002 57146
rect 37014 57094 37066 57146
rect 37078 57094 37130 57146
rect 37142 57094 37194 57146
rect 37206 57094 37258 57146
rect 26240 56992 26292 57044
rect 35164 56992 35216 57044
rect 9036 56924 9088 56976
rect 39856 56924 39908 56976
rect 10140 56899 10192 56908
rect 10140 56865 10149 56899
rect 10149 56865 10183 56899
rect 10183 56865 10192 56899
rect 10140 56856 10192 56865
rect 10692 56856 10744 56908
rect 5080 56788 5132 56840
rect 10784 56831 10836 56840
rect 10784 56797 10793 56831
rect 10793 56797 10827 56831
rect 10827 56797 10836 56831
rect 10784 56788 10836 56797
rect 19800 56856 19852 56908
rect 31116 56856 31168 56908
rect 16304 56788 16356 56840
rect 26148 56788 26200 56840
rect 26240 56788 26292 56840
rect 19984 56652 20036 56704
rect 2610 56550 2662 56602
rect 2674 56550 2726 56602
rect 2738 56550 2790 56602
rect 2802 56550 2854 56602
rect 2866 56550 2918 56602
rect 7610 56550 7662 56602
rect 7674 56550 7726 56602
rect 7738 56550 7790 56602
rect 7802 56550 7854 56602
rect 7866 56550 7918 56602
rect 12610 56550 12662 56602
rect 12674 56550 12726 56602
rect 12738 56550 12790 56602
rect 12802 56550 12854 56602
rect 12866 56550 12918 56602
rect 17610 56550 17662 56602
rect 17674 56550 17726 56602
rect 17738 56550 17790 56602
rect 17802 56550 17854 56602
rect 17866 56550 17918 56602
rect 22610 56550 22662 56602
rect 22674 56550 22726 56602
rect 22738 56550 22790 56602
rect 22802 56550 22854 56602
rect 22866 56550 22918 56602
rect 27610 56550 27662 56602
rect 27674 56550 27726 56602
rect 27738 56550 27790 56602
rect 27802 56550 27854 56602
rect 27866 56550 27918 56602
rect 32610 56550 32662 56602
rect 32674 56550 32726 56602
rect 32738 56550 32790 56602
rect 32802 56550 32854 56602
rect 32866 56550 32918 56602
rect 37610 56550 37662 56602
rect 37674 56550 37726 56602
rect 37738 56550 37790 56602
rect 37802 56550 37854 56602
rect 37866 56550 37918 56602
rect 24216 56176 24268 56228
rect 29092 56176 29144 56228
rect 13820 56108 13872 56160
rect 33968 56108 34020 56160
rect 1950 56006 2002 56058
rect 2014 56006 2066 56058
rect 2078 56006 2130 56058
rect 2142 56006 2194 56058
rect 2206 56006 2258 56058
rect 6950 56006 7002 56058
rect 7014 56006 7066 56058
rect 7078 56006 7130 56058
rect 7142 56006 7194 56058
rect 7206 56006 7258 56058
rect 11950 56006 12002 56058
rect 12014 56006 12066 56058
rect 12078 56006 12130 56058
rect 12142 56006 12194 56058
rect 12206 56006 12258 56058
rect 16950 56006 17002 56058
rect 17014 56006 17066 56058
rect 17078 56006 17130 56058
rect 17142 56006 17194 56058
rect 17206 56006 17258 56058
rect 21950 56006 22002 56058
rect 22014 56006 22066 56058
rect 22078 56006 22130 56058
rect 22142 56006 22194 56058
rect 22206 56006 22258 56058
rect 26950 56006 27002 56058
rect 27014 56006 27066 56058
rect 27078 56006 27130 56058
rect 27142 56006 27194 56058
rect 27206 56006 27258 56058
rect 31950 56006 32002 56058
rect 32014 56006 32066 56058
rect 32078 56006 32130 56058
rect 32142 56006 32194 56058
rect 32206 56006 32258 56058
rect 36950 56006 37002 56058
rect 37014 56006 37066 56058
rect 37078 56006 37130 56058
rect 37142 56006 37194 56058
rect 37206 56006 37258 56058
rect 10692 55904 10744 55956
rect 39304 55904 39356 55956
rect 3792 55836 3844 55888
rect 10968 55836 11020 55888
rect 15936 55879 15988 55888
rect 15936 55845 15945 55879
rect 15945 55845 15979 55879
rect 15979 55845 15988 55879
rect 15936 55836 15988 55845
rect 19432 55836 19484 55888
rect 34704 55836 34756 55888
rect 9404 55768 9456 55820
rect 22376 55768 22428 55820
rect 23204 55768 23256 55820
rect 9496 55743 9548 55752
rect 9496 55709 9505 55743
rect 9505 55709 9539 55743
rect 9539 55709 9548 55743
rect 9496 55700 9548 55709
rect 9956 55743 10008 55752
rect 9956 55709 9964 55743
rect 9964 55709 9998 55743
rect 9998 55709 10008 55743
rect 9956 55700 10008 55709
rect 11704 55700 11756 55752
rect 17960 55700 18012 55752
rect 19248 55700 19300 55752
rect 24124 55632 24176 55684
rect 16304 55607 16356 55616
rect 16304 55573 16313 55607
rect 16313 55573 16347 55607
rect 16347 55573 16356 55607
rect 16304 55564 16356 55573
rect 16488 55607 16540 55616
rect 16488 55573 16497 55607
rect 16497 55573 16531 55607
rect 16531 55573 16540 55607
rect 16488 55564 16540 55573
rect 2610 55462 2662 55514
rect 2674 55462 2726 55514
rect 2738 55462 2790 55514
rect 2802 55462 2854 55514
rect 2866 55462 2918 55514
rect 7610 55462 7662 55514
rect 7674 55462 7726 55514
rect 7738 55462 7790 55514
rect 7802 55462 7854 55514
rect 7866 55462 7918 55514
rect 12610 55462 12662 55514
rect 12674 55462 12726 55514
rect 12738 55462 12790 55514
rect 12802 55462 12854 55514
rect 12866 55462 12918 55514
rect 17610 55462 17662 55514
rect 17674 55462 17726 55514
rect 17738 55462 17790 55514
rect 17802 55462 17854 55514
rect 17866 55462 17918 55514
rect 22610 55462 22662 55514
rect 22674 55462 22726 55514
rect 22738 55462 22790 55514
rect 22802 55462 22854 55514
rect 22866 55462 22918 55514
rect 27610 55462 27662 55514
rect 27674 55462 27726 55514
rect 27738 55462 27790 55514
rect 27802 55462 27854 55514
rect 27866 55462 27918 55514
rect 32610 55462 32662 55514
rect 32674 55462 32726 55514
rect 32738 55462 32790 55514
rect 32802 55462 32854 55514
rect 32866 55462 32918 55514
rect 37610 55462 37662 55514
rect 37674 55462 37726 55514
rect 37738 55462 37790 55514
rect 37802 55462 37854 55514
rect 37866 55462 37918 55514
rect 13728 55292 13780 55344
rect 14464 55292 14516 55344
rect 6184 55224 6236 55276
rect 13452 55156 13504 55208
rect 14648 55156 14700 55208
rect 6276 55020 6328 55072
rect 1950 54918 2002 54970
rect 2014 54918 2066 54970
rect 2078 54918 2130 54970
rect 2142 54918 2194 54970
rect 2206 54918 2258 54970
rect 6950 54918 7002 54970
rect 7014 54918 7066 54970
rect 7078 54918 7130 54970
rect 7142 54918 7194 54970
rect 7206 54918 7258 54970
rect 11950 54918 12002 54970
rect 12014 54918 12066 54970
rect 12078 54918 12130 54970
rect 12142 54918 12194 54970
rect 12206 54918 12258 54970
rect 16950 54918 17002 54970
rect 17014 54918 17066 54970
rect 17078 54918 17130 54970
rect 17142 54918 17194 54970
rect 17206 54918 17258 54970
rect 21950 54918 22002 54970
rect 22014 54918 22066 54970
rect 22078 54918 22130 54970
rect 22142 54918 22194 54970
rect 22206 54918 22258 54970
rect 26950 54918 27002 54970
rect 27014 54918 27066 54970
rect 27078 54918 27130 54970
rect 27142 54918 27194 54970
rect 27206 54918 27258 54970
rect 31950 54918 32002 54970
rect 32014 54918 32066 54970
rect 32078 54918 32130 54970
rect 32142 54918 32194 54970
rect 32206 54918 32258 54970
rect 36950 54918 37002 54970
rect 37014 54918 37066 54970
rect 37078 54918 37130 54970
rect 37142 54918 37194 54970
rect 37206 54918 37258 54970
rect 6736 54680 6788 54732
rect 7472 54680 7524 54732
rect 15476 54723 15528 54732
rect 15476 54689 15485 54723
rect 15485 54689 15519 54723
rect 15519 54689 15528 54723
rect 15476 54680 15528 54689
rect 24860 54680 24912 54732
rect 35072 54748 35124 54800
rect 8208 54612 8260 54664
rect 34888 54680 34940 54732
rect 29920 54612 29972 54664
rect 5540 54587 5592 54596
rect 5540 54553 5549 54587
rect 5549 54553 5583 54587
rect 5583 54553 5592 54587
rect 5540 54544 5592 54553
rect 5908 54544 5960 54596
rect 6552 54587 6604 54596
rect 6552 54553 6561 54587
rect 6561 54553 6595 54587
rect 6595 54553 6604 54587
rect 6552 54544 6604 54553
rect 9312 54544 9364 54596
rect 14372 54544 14424 54596
rect 30288 54544 30340 54596
rect 4252 54519 4304 54528
rect 4252 54485 4261 54519
rect 4261 54485 4295 54519
rect 4295 54485 4304 54519
rect 4252 54476 4304 54485
rect 4712 54476 4764 54528
rect 6736 54519 6788 54528
rect 6736 54485 6745 54519
rect 6745 54485 6779 54519
rect 6779 54485 6788 54519
rect 6736 54476 6788 54485
rect 7104 54519 7156 54528
rect 7104 54485 7113 54519
rect 7113 54485 7147 54519
rect 7147 54485 7156 54519
rect 7104 54476 7156 54485
rect 33968 54519 34020 54528
rect 33968 54485 33977 54519
rect 33977 54485 34011 54519
rect 34011 54485 34020 54519
rect 33968 54476 34020 54485
rect 2610 54374 2662 54426
rect 2674 54374 2726 54426
rect 2738 54374 2790 54426
rect 2802 54374 2854 54426
rect 2866 54374 2918 54426
rect 7610 54374 7662 54426
rect 7674 54374 7726 54426
rect 7738 54374 7790 54426
rect 7802 54374 7854 54426
rect 7866 54374 7918 54426
rect 12610 54374 12662 54426
rect 12674 54374 12726 54426
rect 12738 54374 12790 54426
rect 12802 54374 12854 54426
rect 12866 54374 12918 54426
rect 17610 54374 17662 54426
rect 17674 54374 17726 54426
rect 17738 54374 17790 54426
rect 17802 54374 17854 54426
rect 17866 54374 17918 54426
rect 22610 54374 22662 54426
rect 22674 54374 22726 54426
rect 22738 54374 22790 54426
rect 22802 54374 22854 54426
rect 22866 54374 22918 54426
rect 27610 54374 27662 54426
rect 27674 54374 27726 54426
rect 27738 54374 27790 54426
rect 27802 54374 27854 54426
rect 27866 54374 27918 54426
rect 32610 54374 32662 54426
rect 32674 54374 32726 54426
rect 32738 54374 32790 54426
rect 32802 54374 32854 54426
rect 32866 54374 32918 54426
rect 37610 54374 37662 54426
rect 37674 54374 37726 54426
rect 37738 54374 37790 54426
rect 37802 54374 37854 54426
rect 37866 54374 37918 54426
rect 7104 54272 7156 54324
rect 29920 54272 29972 54324
rect 21548 54204 21600 54256
rect 15292 54136 15344 54188
rect 19156 54136 19208 54188
rect 20352 54136 20404 54188
rect 28080 54136 28132 54188
rect 28264 54179 28316 54188
rect 28264 54145 28273 54179
rect 28273 54145 28307 54179
rect 28307 54145 28316 54179
rect 28264 54136 28316 54145
rect 29000 54179 29052 54188
rect 29000 54145 29009 54179
rect 29009 54145 29043 54179
rect 29043 54145 29052 54179
rect 29000 54136 29052 54145
rect 13176 54000 13228 54052
rect 15936 54000 15988 54052
rect 6092 53932 6144 53984
rect 6552 53932 6604 53984
rect 28356 53975 28408 53984
rect 28356 53941 28365 53975
rect 28365 53941 28399 53975
rect 28399 53941 28408 53975
rect 28356 53932 28408 53941
rect 1950 53830 2002 53882
rect 2014 53830 2066 53882
rect 2078 53830 2130 53882
rect 2142 53830 2194 53882
rect 2206 53830 2258 53882
rect 6950 53830 7002 53882
rect 7014 53830 7066 53882
rect 7078 53830 7130 53882
rect 7142 53830 7194 53882
rect 7206 53830 7258 53882
rect 11950 53830 12002 53882
rect 12014 53830 12066 53882
rect 12078 53830 12130 53882
rect 12142 53830 12194 53882
rect 12206 53830 12258 53882
rect 16950 53830 17002 53882
rect 17014 53830 17066 53882
rect 17078 53830 17130 53882
rect 17142 53830 17194 53882
rect 17206 53830 17258 53882
rect 21950 53830 22002 53882
rect 22014 53830 22066 53882
rect 22078 53830 22130 53882
rect 22142 53830 22194 53882
rect 22206 53830 22258 53882
rect 26950 53830 27002 53882
rect 27014 53830 27066 53882
rect 27078 53830 27130 53882
rect 27142 53830 27194 53882
rect 27206 53830 27258 53882
rect 31950 53830 32002 53882
rect 32014 53830 32066 53882
rect 32078 53830 32130 53882
rect 32142 53830 32194 53882
rect 32206 53830 32258 53882
rect 36950 53830 37002 53882
rect 37014 53830 37066 53882
rect 37078 53830 37130 53882
rect 37142 53830 37194 53882
rect 37206 53830 37258 53882
rect 14924 53660 14976 53712
rect 15384 53660 15436 53712
rect 6000 53592 6052 53644
rect 9312 53592 9364 53644
rect 4436 53524 4488 53576
rect 8208 53456 8260 53508
rect 14924 53456 14976 53508
rect 15384 53567 15436 53576
rect 15384 53533 15393 53567
rect 15393 53533 15427 53567
rect 15427 53533 15436 53567
rect 15384 53524 15436 53533
rect 7288 53388 7340 53440
rect 15292 53431 15344 53440
rect 15292 53397 15301 53431
rect 15301 53397 15335 53431
rect 15335 53397 15344 53431
rect 15292 53388 15344 53397
rect 15476 53499 15528 53508
rect 15476 53465 15485 53499
rect 15485 53465 15519 53499
rect 15519 53465 15528 53499
rect 15476 53456 15528 53465
rect 15844 53499 15896 53508
rect 15844 53465 15853 53499
rect 15853 53465 15887 53499
rect 15887 53465 15896 53499
rect 15844 53456 15896 53465
rect 38292 53567 38344 53576
rect 38292 53533 38301 53567
rect 38301 53533 38335 53567
rect 38335 53533 38344 53567
rect 38292 53524 38344 53533
rect 26792 53456 26844 53508
rect 39212 53499 39264 53508
rect 39212 53465 39221 53499
rect 39221 53465 39255 53499
rect 39255 53465 39264 53499
rect 39212 53456 39264 53465
rect 23112 53388 23164 53440
rect 28448 53388 28500 53440
rect 2610 53286 2662 53338
rect 2674 53286 2726 53338
rect 2738 53286 2790 53338
rect 2802 53286 2854 53338
rect 2866 53286 2918 53338
rect 7610 53286 7662 53338
rect 7674 53286 7726 53338
rect 7738 53286 7790 53338
rect 7802 53286 7854 53338
rect 7866 53286 7918 53338
rect 12610 53286 12662 53338
rect 12674 53286 12726 53338
rect 12738 53286 12790 53338
rect 12802 53286 12854 53338
rect 12866 53286 12918 53338
rect 17610 53286 17662 53338
rect 17674 53286 17726 53338
rect 17738 53286 17790 53338
rect 17802 53286 17854 53338
rect 17866 53286 17918 53338
rect 22610 53286 22662 53338
rect 22674 53286 22726 53338
rect 22738 53286 22790 53338
rect 22802 53286 22854 53338
rect 22866 53286 22918 53338
rect 27610 53286 27662 53338
rect 27674 53286 27726 53338
rect 27738 53286 27790 53338
rect 27802 53286 27854 53338
rect 27866 53286 27918 53338
rect 32610 53286 32662 53338
rect 32674 53286 32726 53338
rect 32738 53286 32790 53338
rect 32802 53286 32854 53338
rect 32866 53286 32918 53338
rect 37610 53286 37662 53338
rect 37674 53286 37726 53338
rect 37738 53286 37790 53338
rect 37802 53286 37854 53338
rect 37866 53286 37918 53338
rect 2504 53116 2556 53168
rect 21732 53116 21784 53168
rect 36452 53116 36504 53168
rect 36728 53116 36780 53168
rect 15292 53091 15344 53100
rect 15292 53057 15301 53091
rect 15301 53057 15335 53091
rect 15335 53057 15344 53091
rect 15292 53048 15344 53057
rect 15568 53091 15620 53100
rect 15568 53057 15577 53091
rect 15577 53057 15611 53091
rect 15611 53057 15620 53091
rect 15568 53048 15620 53057
rect 16212 53048 16264 53100
rect 33692 53048 33744 53100
rect 34060 53048 34112 53100
rect 15936 53023 15988 53032
rect 15936 52989 15945 53023
rect 15945 52989 15979 53023
rect 15979 52989 15988 53023
rect 15936 52980 15988 52989
rect 15200 52912 15252 52964
rect 38752 52912 38804 52964
rect 36728 52887 36780 52896
rect 36728 52853 36737 52887
rect 36737 52853 36771 52887
rect 36771 52853 36780 52887
rect 36728 52844 36780 52853
rect 1950 52742 2002 52794
rect 2014 52742 2066 52794
rect 2078 52742 2130 52794
rect 2142 52742 2194 52794
rect 2206 52742 2258 52794
rect 6950 52742 7002 52794
rect 7014 52742 7066 52794
rect 7078 52742 7130 52794
rect 7142 52742 7194 52794
rect 7206 52742 7258 52794
rect 11950 52742 12002 52794
rect 12014 52742 12066 52794
rect 12078 52742 12130 52794
rect 12142 52742 12194 52794
rect 12206 52742 12258 52794
rect 16950 52742 17002 52794
rect 17014 52742 17066 52794
rect 17078 52742 17130 52794
rect 17142 52742 17194 52794
rect 17206 52742 17258 52794
rect 21950 52742 22002 52794
rect 22014 52742 22066 52794
rect 22078 52742 22130 52794
rect 22142 52742 22194 52794
rect 22206 52742 22258 52794
rect 26950 52742 27002 52794
rect 27014 52742 27066 52794
rect 27078 52742 27130 52794
rect 27142 52742 27194 52794
rect 27206 52742 27258 52794
rect 31950 52742 32002 52794
rect 32014 52742 32066 52794
rect 32078 52742 32130 52794
rect 32142 52742 32194 52794
rect 32206 52742 32258 52794
rect 36950 52742 37002 52794
rect 37014 52742 37066 52794
rect 37078 52742 37130 52794
rect 37142 52742 37194 52794
rect 37206 52742 37258 52794
rect 6000 52640 6052 52692
rect 6552 52640 6604 52692
rect 36820 52640 36872 52692
rect 8208 52572 8260 52624
rect 20996 52572 21048 52624
rect 23480 52572 23532 52624
rect 29460 52572 29512 52624
rect 20536 52504 20588 52556
rect 13912 52436 13964 52488
rect 21732 52436 21784 52488
rect 35808 52479 35860 52488
rect 35808 52445 35817 52479
rect 35817 52445 35851 52479
rect 35851 52445 35860 52479
rect 35808 52436 35860 52445
rect 36544 52479 36596 52488
rect 36544 52445 36553 52479
rect 36553 52445 36587 52479
rect 36587 52445 36596 52479
rect 36544 52436 36596 52445
rect 38200 52436 38252 52488
rect 34704 52411 34756 52420
rect 34704 52377 34713 52411
rect 34713 52377 34747 52411
rect 34747 52377 34756 52411
rect 34704 52368 34756 52377
rect 34888 52343 34940 52352
rect 34888 52309 34897 52343
rect 34897 52309 34931 52343
rect 34931 52309 34940 52343
rect 34888 52300 34940 52309
rect 34980 52343 35032 52352
rect 34980 52309 34989 52343
rect 34989 52309 35023 52343
rect 35023 52309 35032 52343
rect 34980 52300 35032 52309
rect 2610 52198 2662 52250
rect 2674 52198 2726 52250
rect 2738 52198 2790 52250
rect 2802 52198 2854 52250
rect 2866 52198 2918 52250
rect 7610 52198 7662 52250
rect 7674 52198 7726 52250
rect 7738 52198 7790 52250
rect 7802 52198 7854 52250
rect 7866 52198 7918 52250
rect 12610 52198 12662 52250
rect 12674 52198 12726 52250
rect 12738 52198 12790 52250
rect 12802 52198 12854 52250
rect 12866 52198 12918 52250
rect 17610 52198 17662 52250
rect 17674 52198 17726 52250
rect 17738 52198 17790 52250
rect 17802 52198 17854 52250
rect 17866 52198 17918 52250
rect 22610 52198 22662 52250
rect 22674 52198 22726 52250
rect 22738 52198 22790 52250
rect 22802 52198 22854 52250
rect 22866 52198 22918 52250
rect 27610 52198 27662 52250
rect 27674 52198 27726 52250
rect 27738 52198 27790 52250
rect 27802 52198 27854 52250
rect 27866 52198 27918 52250
rect 32610 52198 32662 52250
rect 32674 52198 32726 52250
rect 32738 52198 32790 52250
rect 32802 52198 32854 52250
rect 32866 52198 32918 52250
rect 37610 52198 37662 52250
rect 37674 52198 37726 52250
rect 37738 52198 37790 52250
rect 37802 52198 37854 52250
rect 37866 52198 37918 52250
rect 16856 52096 16908 52148
rect 21640 52096 21692 52148
rect 35808 52139 35860 52148
rect 35808 52105 35817 52139
rect 35817 52105 35851 52139
rect 35851 52105 35860 52139
rect 35808 52096 35860 52105
rect 10876 52028 10928 52080
rect 20536 52028 20588 52080
rect 4896 52003 4948 52012
rect 4896 51969 4905 52003
rect 4905 51969 4939 52003
rect 4939 51969 4948 52003
rect 4896 51960 4948 51969
rect 11244 51960 11296 52012
rect 15384 51960 15436 52012
rect 18144 51892 18196 51944
rect 20628 51935 20680 51944
rect 20628 51901 20637 51935
rect 20637 51901 20671 51935
rect 20671 51901 20680 51935
rect 20628 51892 20680 51901
rect 21456 52028 21508 52080
rect 25688 52028 25740 52080
rect 21548 52003 21600 52012
rect 21548 51969 21557 52003
rect 21557 51969 21591 52003
rect 21591 51969 21600 52003
rect 21548 51960 21600 51969
rect 10784 51824 10836 51876
rect 4988 51756 5040 51808
rect 21640 51892 21692 51944
rect 38292 51960 38344 52012
rect 36268 51935 36320 51944
rect 36268 51901 36277 51935
rect 36277 51901 36311 51935
rect 36311 51901 36320 51935
rect 36268 51892 36320 51901
rect 21732 51756 21784 51808
rect 1950 51654 2002 51706
rect 2014 51654 2066 51706
rect 2078 51654 2130 51706
rect 2142 51654 2194 51706
rect 2206 51654 2258 51706
rect 6950 51654 7002 51706
rect 7014 51654 7066 51706
rect 7078 51654 7130 51706
rect 7142 51654 7194 51706
rect 7206 51654 7258 51706
rect 11950 51654 12002 51706
rect 12014 51654 12066 51706
rect 12078 51654 12130 51706
rect 12142 51654 12194 51706
rect 12206 51654 12258 51706
rect 16950 51654 17002 51706
rect 17014 51654 17066 51706
rect 17078 51654 17130 51706
rect 17142 51654 17194 51706
rect 17206 51654 17258 51706
rect 21950 51654 22002 51706
rect 22014 51654 22066 51706
rect 22078 51654 22130 51706
rect 22142 51654 22194 51706
rect 22206 51654 22258 51706
rect 26950 51654 27002 51706
rect 27014 51654 27066 51706
rect 27078 51654 27130 51706
rect 27142 51654 27194 51706
rect 27206 51654 27258 51706
rect 31950 51654 32002 51706
rect 32014 51654 32066 51706
rect 32078 51654 32130 51706
rect 32142 51654 32194 51706
rect 32206 51654 32258 51706
rect 36950 51654 37002 51706
rect 37014 51654 37066 51706
rect 37078 51654 37130 51706
rect 37142 51654 37194 51706
rect 37206 51654 37258 51706
rect 31760 51391 31812 51400
rect 31760 51357 31769 51391
rect 31769 51357 31803 51391
rect 31803 51357 31812 51391
rect 31760 51348 31812 51357
rect 36820 51348 36872 51400
rect 6828 51280 6880 51332
rect 2610 51110 2662 51162
rect 2674 51110 2726 51162
rect 2738 51110 2790 51162
rect 2802 51110 2854 51162
rect 2866 51110 2918 51162
rect 7610 51110 7662 51162
rect 7674 51110 7726 51162
rect 7738 51110 7790 51162
rect 7802 51110 7854 51162
rect 7866 51110 7918 51162
rect 12610 51110 12662 51162
rect 12674 51110 12726 51162
rect 12738 51110 12790 51162
rect 12802 51110 12854 51162
rect 12866 51110 12918 51162
rect 17610 51110 17662 51162
rect 17674 51110 17726 51162
rect 17738 51110 17790 51162
rect 17802 51110 17854 51162
rect 17866 51110 17918 51162
rect 22610 51110 22662 51162
rect 22674 51110 22726 51162
rect 22738 51110 22790 51162
rect 22802 51110 22854 51162
rect 22866 51110 22918 51162
rect 27610 51110 27662 51162
rect 27674 51110 27726 51162
rect 27738 51110 27790 51162
rect 27802 51110 27854 51162
rect 27866 51110 27918 51162
rect 32610 51110 32662 51162
rect 32674 51110 32726 51162
rect 32738 51110 32790 51162
rect 32802 51110 32854 51162
rect 32866 51110 32918 51162
rect 37610 51110 37662 51162
rect 37674 51110 37726 51162
rect 37738 51110 37790 51162
rect 37802 51110 37854 51162
rect 37866 51110 37918 51162
rect 8208 51008 8260 51060
rect 13452 51008 13504 51060
rect 22284 51008 22336 51060
rect 23112 51008 23164 51060
rect 32404 51008 32456 51060
rect 37464 51008 37516 51060
rect 11612 50940 11664 50992
rect 22376 50940 22428 50992
rect 7932 50872 7984 50924
rect 8208 50872 8260 50924
rect 10692 50915 10744 50924
rect 10692 50881 10701 50915
rect 10701 50881 10735 50915
rect 10735 50881 10744 50915
rect 10692 50872 10744 50881
rect 10876 50915 10928 50924
rect 10876 50881 10885 50915
rect 10885 50881 10919 50915
rect 10919 50881 10928 50915
rect 10876 50872 10928 50881
rect 12992 50915 13044 50924
rect 12992 50881 13001 50915
rect 13001 50881 13044 50915
rect 12992 50872 13044 50881
rect 21824 50915 21876 50924
rect 21824 50881 21833 50915
rect 21833 50881 21867 50915
rect 21867 50881 21876 50915
rect 21824 50872 21876 50881
rect 11428 50804 11480 50856
rect 17500 50804 17552 50856
rect 21732 50804 21784 50856
rect 22284 50915 22336 50924
rect 22284 50881 22293 50915
rect 22293 50881 22327 50915
rect 22327 50881 22336 50915
rect 22284 50872 22336 50881
rect 26148 50804 26200 50856
rect 12440 50711 12492 50720
rect 12440 50677 12449 50711
rect 12449 50677 12483 50711
rect 12483 50677 12492 50711
rect 12440 50668 12492 50677
rect 12808 50711 12860 50720
rect 12808 50677 12817 50711
rect 12817 50677 12851 50711
rect 12851 50677 12860 50711
rect 12808 50668 12860 50677
rect 13268 50668 13320 50720
rect 23204 50668 23256 50720
rect 1950 50566 2002 50618
rect 2014 50566 2066 50618
rect 2078 50566 2130 50618
rect 2142 50566 2194 50618
rect 2206 50566 2258 50618
rect 6950 50566 7002 50618
rect 7014 50566 7066 50618
rect 7078 50566 7130 50618
rect 7142 50566 7194 50618
rect 7206 50566 7258 50618
rect 11950 50566 12002 50618
rect 12014 50566 12066 50618
rect 12078 50566 12130 50618
rect 12142 50566 12194 50618
rect 12206 50566 12258 50618
rect 16950 50566 17002 50618
rect 17014 50566 17066 50618
rect 17078 50566 17130 50618
rect 17142 50566 17194 50618
rect 17206 50566 17258 50618
rect 21950 50566 22002 50618
rect 22014 50566 22066 50618
rect 22078 50566 22130 50618
rect 22142 50566 22194 50618
rect 22206 50566 22258 50618
rect 26950 50566 27002 50618
rect 27014 50566 27066 50618
rect 27078 50566 27130 50618
rect 27142 50566 27194 50618
rect 27206 50566 27258 50618
rect 31950 50566 32002 50618
rect 32014 50566 32066 50618
rect 32078 50566 32130 50618
rect 32142 50566 32194 50618
rect 32206 50566 32258 50618
rect 36950 50566 37002 50618
rect 37014 50566 37066 50618
rect 37078 50566 37130 50618
rect 37142 50566 37194 50618
rect 37206 50566 37258 50618
rect 19892 50464 19944 50516
rect 29828 50464 29880 50516
rect 3056 50396 3108 50448
rect 9220 50396 9272 50448
rect 10600 50396 10652 50448
rect 14188 50396 14240 50448
rect 20628 50396 20680 50448
rect 23480 50396 23532 50448
rect 35256 50396 35308 50448
rect 8024 50328 8076 50380
rect 8208 50328 8260 50380
rect 8944 50260 8996 50312
rect 6736 50192 6788 50244
rect 12808 50260 12860 50312
rect 20536 50260 20588 50312
rect 39672 50328 39724 50380
rect 11612 50192 11664 50244
rect 25596 50124 25648 50176
rect 2610 50022 2662 50074
rect 2674 50022 2726 50074
rect 2738 50022 2790 50074
rect 2802 50022 2854 50074
rect 2866 50022 2918 50074
rect 7610 50022 7662 50074
rect 7674 50022 7726 50074
rect 7738 50022 7790 50074
rect 7802 50022 7854 50074
rect 7866 50022 7918 50074
rect 12610 50022 12662 50074
rect 12674 50022 12726 50074
rect 12738 50022 12790 50074
rect 12802 50022 12854 50074
rect 12866 50022 12918 50074
rect 17610 50022 17662 50074
rect 17674 50022 17726 50074
rect 17738 50022 17790 50074
rect 17802 50022 17854 50074
rect 17866 50022 17918 50074
rect 22610 50022 22662 50074
rect 22674 50022 22726 50074
rect 22738 50022 22790 50074
rect 22802 50022 22854 50074
rect 22866 50022 22918 50074
rect 27610 50022 27662 50074
rect 27674 50022 27726 50074
rect 27738 50022 27790 50074
rect 27802 50022 27854 50074
rect 27866 50022 27918 50074
rect 32610 50022 32662 50074
rect 32674 50022 32726 50074
rect 32738 50022 32790 50074
rect 32802 50022 32854 50074
rect 32866 50022 32918 50074
rect 37610 50022 37662 50074
rect 37674 50022 37726 50074
rect 37738 50022 37790 50074
rect 37802 50022 37854 50074
rect 37866 50022 37918 50074
rect 3884 49920 3936 49972
rect 7288 49852 7340 49904
rect 23112 49920 23164 49972
rect 1400 49827 1452 49836
rect 1400 49793 1409 49827
rect 1409 49793 1443 49827
rect 1443 49793 1452 49827
rect 1400 49784 1452 49793
rect 13912 49827 13964 49836
rect 13912 49793 13921 49827
rect 13921 49793 13955 49827
rect 13955 49793 13964 49827
rect 13912 49784 13964 49793
rect 14188 49827 14240 49836
rect 14188 49793 14197 49827
rect 14197 49793 14231 49827
rect 14231 49793 14240 49827
rect 14188 49784 14240 49793
rect 23664 49827 23716 49836
rect 23664 49793 23673 49827
rect 23673 49793 23707 49827
rect 23707 49793 23716 49827
rect 23664 49784 23716 49793
rect 23756 49784 23808 49836
rect 8944 49716 8996 49768
rect 11152 49716 11204 49768
rect 22376 49716 22428 49768
rect 23112 49716 23164 49768
rect 23572 49716 23624 49768
rect 24308 49827 24360 49836
rect 24308 49793 24317 49827
rect 24317 49793 24351 49827
rect 24351 49793 24360 49827
rect 24308 49784 24360 49793
rect 24676 49827 24728 49836
rect 24676 49793 24685 49827
rect 24685 49793 24719 49827
rect 24719 49793 24728 49827
rect 24676 49784 24728 49793
rect 33784 49784 33836 49836
rect 35808 49827 35860 49836
rect 35808 49793 35817 49827
rect 35817 49793 35851 49827
rect 35851 49793 35860 49827
rect 35808 49784 35860 49793
rect 25044 49759 25096 49768
rect 25044 49725 25053 49759
rect 25053 49725 25087 49759
rect 25087 49725 25096 49759
rect 25044 49716 25096 49725
rect 31576 49716 31628 49768
rect 36636 49827 36688 49836
rect 36636 49793 36645 49827
rect 36645 49793 36679 49827
rect 36679 49793 36688 49827
rect 36636 49784 36688 49793
rect 40500 49827 40552 49836
rect 40500 49793 40509 49827
rect 40509 49793 40543 49827
rect 40543 49793 40552 49827
rect 40500 49784 40552 49793
rect 13084 49648 13136 49700
rect 13360 49648 13412 49700
rect 29552 49648 29604 49700
rect 33784 49648 33836 49700
rect 34152 49648 34204 49700
rect 1950 49478 2002 49530
rect 2014 49478 2066 49530
rect 2078 49478 2130 49530
rect 2142 49478 2194 49530
rect 2206 49478 2258 49530
rect 6950 49478 7002 49530
rect 7014 49478 7066 49530
rect 7078 49478 7130 49530
rect 7142 49478 7194 49530
rect 7206 49478 7258 49530
rect 11950 49478 12002 49530
rect 12014 49478 12066 49530
rect 12078 49478 12130 49530
rect 12142 49478 12194 49530
rect 12206 49478 12258 49530
rect 16950 49478 17002 49530
rect 17014 49478 17066 49530
rect 17078 49478 17130 49530
rect 17142 49478 17194 49530
rect 17206 49478 17258 49530
rect 21950 49478 22002 49530
rect 22014 49478 22066 49530
rect 22078 49478 22130 49530
rect 22142 49478 22194 49530
rect 22206 49478 22258 49530
rect 26950 49478 27002 49530
rect 27014 49478 27066 49530
rect 27078 49478 27130 49530
rect 27142 49478 27194 49530
rect 27206 49478 27258 49530
rect 31950 49478 32002 49530
rect 32014 49478 32066 49530
rect 32078 49478 32130 49530
rect 32142 49478 32194 49530
rect 32206 49478 32258 49530
rect 36950 49478 37002 49530
rect 37014 49478 37066 49530
rect 37078 49478 37130 49530
rect 37142 49478 37194 49530
rect 37206 49478 37258 49530
rect 22284 49308 22336 49360
rect 23480 49308 23532 49360
rect 20168 49240 20220 49292
rect 24400 49215 24452 49224
rect 24400 49181 24409 49215
rect 24409 49181 24443 49215
rect 24443 49181 24452 49215
rect 24400 49172 24452 49181
rect 19248 49036 19300 49088
rect 37372 49104 37424 49156
rect 24860 49079 24912 49088
rect 24860 49045 24869 49079
rect 24869 49045 24903 49079
rect 24903 49045 24912 49079
rect 24860 49036 24912 49045
rect 2610 48934 2662 48986
rect 2674 48934 2726 48986
rect 2738 48934 2790 48986
rect 2802 48934 2854 48986
rect 2866 48934 2918 48986
rect 7610 48934 7662 48986
rect 7674 48934 7726 48986
rect 7738 48934 7790 48986
rect 7802 48934 7854 48986
rect 7866 48934 7918 48986
rect 12610 48934 12662 48986
rect 12674 48934 12726 48986
rect 12738 48934 12790 48986
rect 12802 48934 12854 48986
rect 12866 48934 12918 48986
rect 17610 48934 17662 48986
rect 17674 48934 17726 48986
rect 17738 48934 17790 48986
rect 17802 48934 17854 48986
rect 17866 48934 17918 48986
rect 22610 48934 22662 48986
rect 22674 48934 22726 48986
rect 22738 48934 22790 48986
rect 22802 48934 22854 48986
rect 22866 48934 22918 48986
rect 27610 48934 27662 48986
rect 27674 48934 27726 48986
rect 27738 48934 27790 48986
rect 27802 48934 27854 48986
rect 27866 48934 27918 48986
rect 32610 48934 32662 48986
rect 32674 48934 32726 48986
rect 32738 48934 32790 48986
rect 32802 48934 32854 48986
rect 32866 48934 32918 48986
rect 37610 48934 37662 48986
rect 37674 48934 37726 48986
rect 37738 48934 37790 48986
rect 37802 48934 37854 48986
rect 37866 48934 37918 48986
rect 16580 48832 16632 48884
rect 37372 48875 37424 48884
rect 37372 48841 37381 48875
rect 37381 48841 37415 48875
rect 37415 48841 37424 48875
rect 37372 48832 37424 48841
rect 13360 48764 13412 48816
rect 11428 48696 11480 48748
rect 19984 48764 20036 48816
rect 8944 48628 8996 48680
rect 11520 48628 11572 48680
rect 16948 48628 17000 48680
rect 17316 48696 17368 48748
rect 22376 48739 22428 48748
rect 22376 48705 22385 48739
rect 22385 48705 22419 48739
rect 22419 48705 22428 48739
rect 22376 48696 22428 48705
rect 24124 48696 24176 48748
rect 32956 48696 33008 48748
rect 38384 48696 38436 48748
rect 17408 48628 17460 48680
rect 37464 48628 37516 48680
rect 10692 48603 10744 48612
rect 10692 48569 10701 48603
rect 10701 48569 10735 48603
rect 10735 48569 10744 48603
rect 10692 48560 10744 48569
rect 13728 48560 13780 48612
rect 11428 48492 11480 48544
rect 16764 48492 16816 48544
rect 16948 48492 17000 48544
rect 22284 48492 22336 48544
rect 1950 48390 2002 48442
rect 2014 48390 2066 48442
rect 2078 48390 2130 48442
rect 2142 48390 2194 48442
rect 2206 48390 2258 48442
rect 6950 48390 7002 48442
rect 7014 48390 7066 48442
rect 7078 48390 7130 48442
rect 7142 48390 7194 48442
rect 7206 48390 7258 48442
rect 11950 48390 12002 48442
rect 12014 48390 12066 48442
rect 12078 48390 12130 48442
rect 12142 48390 12194 48442
rect 12206 48390 12258 48442
rect 16950 48390 17002 48442
rect 17014 48390 17066 48442
rect 17078 48390 17130 48442
rect 17142 48390 17194 48442
rect 17206 48390 17258 48442
rect 21950 48390 22002 48442
rect 22014 48390 22066 48442
rect 22078 48390 22130 48442
rect 22142 48390 22194 48442
rect 22206 48390 22258 48442
rect 26950 48390 27002 48442
rect 27014 48390 27066 48442
rect 27078 48390 27130 48442
rect 27142 48390 27194 48442
rect 27206 48390 27258 48442
rect 31950 48390 32002 48442
rect 32014 48390 32066 48442
rect 32078 48390 32130 48442
rect 32142 48390 32194 48442
rect 32206 48390 32258 48442
rect 36950 48390 37002 48442
rect 37014 48390 37066 48442
rect 37078 48390 37130 48442
rect 37142 48390 37194 48442
rect 37206 48390 37258 48442
rect 13544 48288 13596 48340
rect 24860 48288 24912 48340
rect 10508 48220 10560 48272
rect 11336 48220 11388 48272
rect 14096 48084 14148 48136
rect 19156 48084 19208 48136
rect 6460 47948 6512 48000
rect 14740 47948 14792 48000
rect 19156 47948 19208 48000
rect 38844 47948 38896 48000
rect 2610 47846 2662 47898
rect 2674 47846 2726 47898
rect 2738 47846 2790 47898
rect 2802 47846 2854 47898
rect 2866 47846 2918 47898
rect 7610 47846 7662 47898
rect 7674 47846 7726 47898
rect 7738 47846 7790 47898
rect 7802 47846 7854 47898
rect 7866 47846 7918 47898
rect 12610 47846 12662 47898
rect 12674 47846 12726 47898
rect 12738 47846 12790 47898
rect 12802 47846 12854 47898
rect 12866 47846 12918 47898
rect 17610 47846 17662 47898
rect 17674 47846 17726 47898
rect 17738 47846 17790 47898
rect 17802 47846 17854 47898
rect 17866 47846 17918 47898
rect 22610 47846 22662 47898
rect 22674 47846 22726 47898
rect 22738 47846 22790 47898
rect 22802 47846 22854 47898
rect 22866 47846 22918 47898
rect 27610 47846 27662 47898
rect 27674 47846 27726 47898
rect 27738 47846 27790 47898
rect 27802 47846 27854 47898
rect 27866 47846 27918 47898
rect 32610 47846 32662 47898
rect 32674 47846 32726 47898
rect 32738 47846 32790 47898
rect 32802 47846 32854 47898
rect 32866 47846 32918 47898
rect 37610 47846 37662 47898
rect 37674 47846 37726 47898
rect 37738 47846 37790 47898
rect 37802 47846 37854 47898
rect 37866 47846 37918 47898
rect 14464 47744 14516 47796
rect 38844 47744 38896 47796
rect 9680 47676 9732 47728
rect 35808 47676 35860 47728
rect 3976 47608 4028 47660
rect 21824 47608 21876 47660
rect 27988 47608 28040 47660
rect 2320 47540 2372 47592
rect 28172 47540 28224 47592
rect 29920 47540 29972 47592
rect 1950 47302 2002 47354
rect 2014 47302 2066 47354
rect 2078 47302 2130 47354
rect 2142 47302 2194 47354
rect 2206 47302 2258 47354
rect 6950 47302 7002 47354
rect 7014 47302 7066 47354
rect 7078 47302 7130 47354
rect 7142 47302 7194 47354
rect 7206 47302 7258 47354
rect 11950 47302 12002 47354
rect 12014 47302 12066 47354
rect 12078 47302 12130 47354
rect 12142 47302 12194 47354
rect 12206 47302 12258 47354
rect 16950 47302 17002 47354
rect 17014 47302 17066 47354
rect 17078 47302 17130 47354
rect 17142 47302 17194 47354
rect 17206 47302 17258 47354
rect 21950 47302 22002 47354
rect 22014 47302 22066 47354
rect 22078 47302 22130 47354
rect 22142 47302 22194 47354
rect 22206 47302 22258 47354
rect 26950 47302 27002 47354
rect 27014 47302 27066 47354
rect 27078 47302 27130 47354
rect 27142 47302 27194 47354
rect 27206 47302 27258 47354
rect 31950 47302 32002 47354
rect 32014 47302 32066 47354
rect 32078 47302 32130 47354
rect 32142 47302 32194 47354
rect 32206 47302 32258 47354
rect 36950 47302 37002 47354
rect 37014 47302 37066 47354
rect 37078 47302 37130 47354
rect 37142 47302 37194 47354
rect 37206 47302 37258 47354
rect 25872 46928 25924 46980
rect 31300 46928 31352 46980
rect 2610 46758 2662 46810
rect 2674 46758 2726 46810
rect 2738 46758 2790 46810
rect 2802 46758 2854 46810
rect 2866 46758 2918 46810
rect 7610 46758 7662 46810
rect 7674 46758 7726 46810
rect 7738 46758 7790 46810
rect 7802 46758 7854 46810
rect 7866 46758 7918 46810
rect 12610 46758 12662 46810
rect 12674 46758 12726 46810
rect 12738 46758 12790 46810
rect 12802 46758 12854 46810
rect 12866 46758 12918 46810
rect 17610 46758 17662 46810
rect 17674 46758 17726 46810
rect 17738 46758 17790 46810
rect 17802 46758 17854 46810
rect 17866 46758 17918 46810
rect 22610 46758 22662 46810
rect 22674 46758 22726 46810
rect 22738 46758 22790 46810
rect 22802 46758 22854 46810
rect 22866 46758 22918 46810
rect 27610 46758 27662 46810
rect 27674 46758 27726 46810
rect 27738 46758 27790 46810
rect 27802 46758 27854 46810
rect 27866 46758 27918 46810
rect 32610 46758 32662 46810
rect 32674 46758 32726 46810
rect 32738 46758 32790 46810
rect 32802 46758 32854 46810
rect 32866 46758 32918 46810
rect 37610 46758 37662 46810
rect 37674 46758 37726 46810
rect 37738 46758 37790 46810
rect 37802 46758 37854 46810
rect 37866 46758 37918 46810
rect 14464 46520 14516 46572
rect 22376 46520 22428 46572
rect 20628 46452 20680 46504
rect 30380 46452 30432 46504
rect 10324 46384 10376 46436
rect 20352 46384 20404 46436
rect 22376 46384 22428 46436
rect 23020 46384 23072 46436
rect 23204 46384 23256 46436
rect 39488 46384 39540 46436
rect 10784 46316 10836 46368
rect 36728 46316 36780 46368
rect 1950 46214 2002 46266
rect 2014 46214 2066 46266
rect 2078 46214 2130 46266
rect 2142 46214 2194 46266
rect 2206 46214 2258 46266
rect 6950 46214 7002 46266
rect 7014 46214 7066 46266
rect 7078 46214 7130 46266
rect 7142 46214 7194 46266
rect 7206 46214 7258 46266
rect 11950 46214 12002 46266
rect 12014 46214 12066 46266
rect 12078 46214 12130 46266
rect 12142 46214 12194 46266
rect 12206 46214 12258 46266
rect 16950 46214 17002 46266
rect 17014 46214 17066 46266
rect 17078 46214 17130 46266
rect 17142 46214 17194 46266
rect 17206 46214 17258 46266
rect 21950 46214 22002 46266
rect 22014 46214 22066 46266
rect 22078 46214 22130 46266
rect 22142 46214 22194 46266
rect 22206 46214 22258 46266
rect 26950 46214 27002 46266
rect 27014 46214 27066 46266
rect 27078 46214 27130 46266
rect 27142 46214 27194 46266
rect 27206 46214 27258 46266
rect 31950 46214 32002 46266
rect 32014 46214 32066 46266
rect 32078 46214 32130 46266
rect 32142 46214 32194 46266
rect 32206 46214 32258 46266
rect 36950 46214 37002 46266
rect 37014 46214 37066 46266
rect 37078 46214 37130 46266
rect 37142 46214 37194 46266
rect 37206 46214 37258 46266
rect 23020 46112 23072 46164
rect 23388 46112 23440 46164
rect 30380 45976 30432 46028
rect 31300 45976 31352 46028
rect 18144 45840 18196 45892
rect 31024 45840 31076 45892
rect 2610 45670 2662 45722
rect 2674 45670 2726 45722
rect 2738 45670 2790 45722
rect 2802 45670 2854 45722
rect 2866 45670 2918 45722
rect 7610 45670 7662 45722
rect 7674 45670 7726 45722
rect 7738 45670 7790 45722
rect 7802 45670 7854 45722
rect 7866 45670 7918 45722
rect 12610 45670 12662 45722
rect 12674 45670 12726 45722
rect 12738 45670 12790 45722
rect 12802 45670 12854 45722
rect 12866 45670 12918 45722
rect 17610 45670 17662 45722
rect 17674 45670 17726 45722
rect 17738 45670 17790 45722
rect 17802 45670 17854 45722
rect 17866 45670 17918 45722
rect 22610 45670 22662 45722
rect 22674 45670 22726 45722
rect 22738 45670 22790 45722
rect 22802 45670 22854 45722
rect 22866 45670 22918 45722
rect 27610 45670 27662 45722
rect 27674 45670 27726 45722
rect 27738 45670 27790 45722
rect 27802 45670 27854 45722
rect 27866 45670 27918 45722
rect 32610 45670 32662 45722
rect 32674 45670 32726 45722
rect 32738 45670 32790 45722
rect 32802 45670 32854 45722
rect 32866 45670 32918 45722
rect 37610 45670 37662 45722
rect 37674 45670 37726 45722
rect 37738 45670 37790 45722
rect 37802 45670 37854 45722
rect 37866 45670 37918 45722
rect 3424 45432 3476 45484
rect 20168 45500 20220 45552
rect 23204 45543 23256 45552
rect 23204 45509 23213 45543
rect 23213 45509 23247 45543
rect 23247 45509 23256 45543
rect 23204 45500 23256 45509
rect 23756 45500 23808 45552
rect 8944 45432 8996 45484
rect 9036 45364 9088 45416
rect 6460 45228 6512 45280
rect 20168 45228 20220 45280
rect 24492 45271 24544 45280
rect 24492 45237 24501 45271
rect 24501 45237 24535 45271
rect 24535 45237 24544 45271
rect 24492 45228 24544 45237
rect 1950 45126 2002 45178
rect 2014 45126 2066 45178
rect 2078 45126 2130 45178
rect 2142 45126 2194 45178
rect 2206 45126 2258 45178
rect 6950 45126 7002 45178
rect 7014 45126 7066 45178
rect 7078 45126 7130 45178
rect 7142 45126 7194 45178
rect 7206 45126 7258 45178
rect 11950 45126 12002 45178
rect 12014 45126 12066 45178
rect 12078 45126 12130 45178
rect 12142 45126 12194 45178
rect 12206 45126 12258 45178
rect 16950 45126 17002 45178
rect 17014 45126 17066 45178
rect 17078 45126 17130 45178
rect 17142 45126 17194 45178
rect 17206 45126 17258 45178
rect 21950 45126 22002 45178
rect 22014 45126 22066 45178
rect 22078 45126 22130 45178
rect 22142 45126 22194 45178
rect 22206 45126 22258 45178
rect 26950 45126 27002 45178
rect 27014 45126 27066 45178
rect 27078 45126 27130 45178
rect 27142 45126 27194 45178
rect 27206 45126 27258 45178
rect 31950 45126 32002 45178
rect 32014 45126 32066 45178
rect 32078 45126 32130 45178
rect 32142 45126 32194 45178
rect 32206 45126 32258 45178
rect 36950 45126 37002 45178
rect 37014 45126 37066 45178
rect 37078 45126 37130 45178
rect 37142 45126 37194 45178
rect 37206 45126 37258 45178
rect 10416 44956 10468 45008
rect 19524 44956 19576 45008
rect 12348 44888 12400 44940
rect 19800 44931 19852 44940
rect 19800 44897 19809 44931
rect 19809 44897 19843 44931
rect 19843 44897 19852 44931
rect 19800 44888 19852 44897
rect 21364 44956 21416 45008
rect 38752 44956 38804 45008
rect 26884 44888 26936 44940
rect 30104 44888 30156 44940
rect 32404 44931 32456 44940
rect 32404 44897 32413 44931
rect 32413 44897 32447 44931
rect 32447 44897 32456 44931
rect 32404 44888 32456 44897
rect 6460 44820 6512 44872
rect 6736 44863 6788 44872
rect 6736 44829 6745 44863
rect 6745 44829 6779 44863
rect 6779 44829 6788 44863
rect 6736 44820 6788 44829
rect 22376 44820 22428 44872
rect 31852 44752 31904 44804
rect 32588 44820 32640 44872
rect 19432 44727 19484 44736
rect 19432 44693 19441 44727
rect 19441 44693 19475 44727
rect 19475 44693 19484 44727
rect 19432 44684 19484 44693
rect 32312 44684 32364 44736
rect 2610 44582 2662 44634
rect 2674 44582 2726 44634
rect 2738 44582 2790 44634
rect 2802 44582 2854 44634
rect 2866 44582 2918 44634
rect 7610 44582 7662 44634
rect 7674 44582 7726 44634
rect 7738 44582 7790 44634
rect 7802 44582 7854 44634
rect 7866 44582 7918 44634
rect 12610 44582 12662 44634
rect 12674 44582 12726 44634
rect 12738 44582 12790 44634
rect 12802 44582 12854 44634
rect 12866 44582 12918 44634
rect 17610 44582 17662 44634
rect 17674 44582 17726 44634
rect 17738 44582 17790 44634
rect 17802 44582 17854 44634
rect 17866 44582 17918 44634
rect 22610 44582 22662 44634
rect 22674 44582 22726 44634
rect 22738 44582 22790 44634
rect 22802 44582 22854 44634
rect 22866 44582 22918 44634
rect 27610 44582 27662 44634
rect 27674 44582 27726 44634
rect 27738 44582 27790 44634
rect 27802 44582 27854 44634
rect 27866 44582 27918 44634
rect 32610 44582 32662 44634
rect 32674 44582 32726 44634
rect 32738 44582 32790 44634
rect 32802 44582 32854 44634
rect 32866 44582 32918 44634
rect 37610 44582 37662 44634
rect 37674 44582 37726 44634
rect 37738 44582 37790 44634
rect 37802 44582 37854 44634
rect 37866 44582 37918 44634
rect 18696 44480 18748 44532
rect 19064 44480 19116 44532
rect 12440 44412 12492 44464
rect 9220 44344 9272 44396
rect 19064 44344 19116 44396
rect 9956 44276 10008 44328
rect 19156 44276 19208 44328
rect 9496 44208 9548 44260
rect 10232 44251 10284 44260
rect 10232 44217 10241 44251
rect 10241 44217 10275 44251
rect 10275 44217 10284 44251
rect 10232 44208 10284 44217
rect 26884 44412 26936 44464
rect 33600 44412 33652 44464
rect 34980 44276 35032 44328
rect 35440 44276 35492 44328
rect 35900 44208 35952 44260
rect 36452 44208 36504 44260
rect 4896 44140 4948 44192
rect 5080 44183 5132 44192
rect 5080 44149 5089 44183
rect 5089 44149 5123 44183
rect 5123 44149 5132 44183
rect 5080 44140 5132 44149
rect 9036 44140 9088 44192
rect 9312 44140 9364 44192
rect 9956 44140 10008 44192
rect 14280 44140 14332 44192
rect 33692 44140 33744 44192
rect 1950 44038 2002 44090
rect 2014 44038 2066 44090
rect 2078 44038 2130 44090
rect 2142 44038 2194 44090
rect 2206 44038 2258 44090
rect 6950 44038 7002 44090
rect 7014 44038 7066 44090
rect 7078 44038 7130 44090
rect 7142 44038 7194 44090
rect 7206 44038 7258 44090
rect 11950 44038 12002 44090
rect 12014 44038 12066 44090
rect 12078 44038 12130 44090
rect 12142 44038 12194 44090
rect 12206 44038 12258 44090
rect 16950 44038 17002 44090
rect 17014 44038 17066 44090
rect 17078 44038 17130 44090
rect 17142 44038 17194 44090
rect 17206 44038 17258 44090
rect 21950 44038 22002 44090
rect 22014 44038 22066 44090
rect 22078 44038 22130 44090
rect 22142 44038 22194 44090
rect 22206 44038 22258 44090
rect 26950 44038 27002 44090
rect 27014 44038 27066 44090
rect 27078 44038 27130 44090
rect 27142 44038 27194 44090
rect 27206 44038 27258 44090
rect 31950 44038 32002 44090
rect 32014 44038 32066 44090
rect 32078 44038 32130 44090
rect 32142 44038 32194 44090
rect 32206 44038 32258 44090
rect 36950 44038 37002 44090
rect 37014 44038 37066 44090
rect 37078 44038 37130 44090
rect 37142 44038 37194 44090
rect 37206 44038 37258 44090
rect 19616 43936 19668 43988
rect 32496 43936 32548 43988
rect 25964 43596 26016 43648
rect 36636 43596 36688 43648
rect 2610 43494 2662 43546
rect 2674 43494 2726 43546
rect 2738 43494 2790 43546
rect 2802 43494 2854 43546
rect 2866 43494 2918 43546
rect 7610 43494 7662 43546
rect 7674 43494 7726 43546
rect 7738 43494 7790 43546
rect 7802 43494 7854 43546
rect 7866 43494 7918 43546
rect 12610 43494 12662 43546
rect 12674 43494 12726 43546
rect 12738 43494 12790 43546
rect 12802 43494 12854 43546
rect 12866 43494 12918 43546
rect 17610 43494 17662 43546
rect 17674 43494 17726 43546
rect 17738 43494 17790 43546
rect 17802 43494 17854 43546
rect 17866 43494 17918 43546
rect 22610 43494 22662 43546
rect 22674 43494 22726 43546
rect 22738 43494 22790 43546
rect 22802 43494 22854 43546
rect 22866 43494 22918 43546
rect 27610 43494 27662 43546
rect 27674 43494 27726 43546
rect 27738 43494 27790 43546
rect 27802 43494 27854 43546
rect 27866 43494 27918 43546
rect 32610 43494 32662 43546
rect 32674 43494 32726 43546
rect 32738 43494 32790 43546
rect 32802 43494 32854 43546
rect 32866 43494 32918 43546
rect 37610 43494 37662 43546
rect 37674 43494 37726 43546
rect 37738 43494 37790 43546
rect 37802 43494 37854 43546
rect 37866 43494 37918 43546
rect 10876 43392 10928 43444
rect 5080 43324 5132 43376
rect 14188 43392 14240 43444
rect 33048 43392 33100 43444
rect 9588 43299 9640 43308
rect 9588 43265 9597 43299
rect 9597 43265 9631 43299
rect 9631 43265 9640 43299
rect 9588 43256 9640 43265
rect 9680 43299 9732 43308
rect 9680 43265 9689 43299
rect 9689 43265 9723 43299
rect 9723 43265 9732 43299
rect 9680 43256 9732 43265
rect 10048 43256 10100 43308
rect 9404 43095 9456 43104
rect 9404 43061 9413 43095
rect 9413 43061 9447 43095
rect 9447 43061 9456 43095
rect 9404 43052 9456 43061
rect 10508 43188 10560 43240
rect 11244 43188 11296 43240
rect 11428 43188 11480 43240
rect 27988 43256 28040 43308
rect 16580 43188 16632 43240
rect 16764 43188 16816 43240
rect 12348 43120 12400 43172
rect 16764 43052 16816 43104
rect 19616 43052 19668 43104
rect 1950 42950 2002 43002
rect 2014 42950 2066 43002
rect 2078 42950 2130 43002
rect 2142 42950 2194 43002
rect 2206 42950 2258 43002
rect 6950 42950 7002 43002
rect 7014 42950 7066 43002
rect 7078 42950 7130 43002
rect 7142 42950 7194 43002
rect 7206 42950 7258 43002
rect 11950 42950 12002 43002
rect 12014 42950 12066 43002
rect 12078 42950 12130 43002
rect 12142 42950 12194 43002
rect 12206 42950 12258 43002
rect 16950 42950 17002 43002
rect 17014 42950 17066 43002
rect 17078 42950 17130 43002
rect 17142 42950 17194 43002
rect 17206 42950 17258 43002
rect 21950 42950 22002 43002
rect 22014 42950 22066 43002
rect 22078 42950 22130 43002
rect 22142 42950 22194 43002
rect 22206 42950 22258 43002
rect 26950 42950 27002 43002
rect 27014 42950 27066 43002
rect 27078 42950 27130 43002
rect 27142 42950 27194 43002
rect 27206 42950 27258 43002
rect 31950 42950 32002 43002
rect 32014 42950 32066 43002
rect 32078 42950 32130 43002
rect 32142 42950 32194 43002
rect 32206 42950 32258 43002
rect 36950 42950 37002 43002
rect 37014 42950 37066 43002
rect 37078 42950 37130 43002
rect 37142 42950 37194 43002
rect 37206 42950 37258 43002
rect 22192 42848 22244 42900
rect 23204 42848 23256 42900
rect 21548 42823 21600 42832
rect 21548 42789 21557 42823
rect 21557 42789 21591 42823
rect 21591 42789 21600 42823
rect 21548 42780 21600 42789
rect 3056 42712 3108 42764
rect 8392 42712 8444 42764
rect 19524 42712 19576 42764
rect 12992 42644 13044 42696
rect 22284 42712 22336 42764
rect 22744 42712 22796 42764
rect 23940 42712 23992 42764
rect 18604 42576 18656 42628
rect 19156 42576 19208 42628
rect 22100 42644 22152 42696
rect 21180 42576 21232 42628
rect 23388 42644 23440 42696
rect 5172 42508 5224 42560
rect 23204 42576 23256 42628
rect 22376 42508 22428 42560
rect 22744 42551 22796 42560
rect 22744 42517 22753 42551
rect 22753 42517 22787 42551
rect 22787 42517 22796 42551
rect 22744 42508 22796 42517
rect 23388 42508 23440 42560
rect 2610 42406 2662 42458
rect 2674 42406 2726 42458
rect 2738 42406 2790 42458
rect 2802 42406 2854 42458
rect 2866 42406 2918 42458
rect 7610 42406 7662 42458
rect 7674 42406 7726 42458
rect 7738 42406 7790 42458
rect 7802 42406 7854 42458
rect 7866 42406 7918 42458
rect 12610 42406 12662 42458
rect 12674 42406 12726 42458
rect 12738 42406 12790 42458
rect 12802 42406 12854 42458
rect 12866 42406 12918 42458
rect 17610 42406 17662 42458
rect 17674 42406 17726 42458
rect 17738 42406 17790 42458
rect 17802 42406 17854 42458
rect 17866 42406 17918 42458
rect 22610 42406 22662 42458
rect 22674 42406 22726 42458
rect 22738 42406 22790 42458
rect 22802 42406 22854 42458
rect 22866 42406 22918 42458
rect 27610 42406 27662 42458
rect 27674 42406 27726 42458
rect 27738 42406 27790 42458
rect 27802 42406 27854 42458
rect 27866 42406 27918 42458
rect 32610 42406 32662 42458
rect 32674 42406 32726 42458
rect 32738 42406 32790 42458
rect 32802 42406 32854 42458
rect 32866 42406 32918 42458
rect 37610 42406 37662 42458
rect 37674 42406 37726 42458
rect 37738 42406 37790 42458
rect 37802 42406 37854 42458
rect 37866 42406 37918 42458
rect 14004 42304 14056 42356
rect 25688 42304 25740 42356
rect 18512 42236 18564 42288
rect 19892 42168 19944 42220
rect 22376 42168 22428 42220
rect 5540 42032 5592 42084
rect 6092 42032 6144 42084
rect 18604 42032 18656 42084
rect 23572 42211 23624 42220
rect 23572 42177 23581 42211
rect 23581 42177 23615 42211
rect 23615 42177 23624 42211
rect 23572 42168 23624 42177
rect 23664 42211 23716 42220
rect 23664 42177 23673 42211
rect 23673 42177 23707 42211
rect 23707 42177 23716 42211
rect 23664 42168 23716 42177
rect 24676 42236 24728 42288
rect 27988 42236 28040 42288
rect 24032 42168 24084 42220
rect 24308 42168 24360 42220
rect 26332 42168 26384 42220
rect 26792 42168 26844 42220
rect 27344 42168 27396 42220
rect 26056 42100 26108 42152
rect 29552 42100 29604 42152
rect 32864 42143 32916 42152
rect 32864 42109 32873 42143
rect 32873 42109 32907 42143
rect 32907 42109 32916 42143
rect 32864 42100 32916 42109
rect 33232 42168 33284 42220
rect 36084 42100 36136 42152
rect 23940 42032 23992 42084
rect 35992 42032 36044 42084
rect 26424 41964 26476 42016
rect 1950 41862 2002 41914
rect 2014 41862 2066 41914
rect 2078 41862 2130 41914
rect 2142 41862 2194 41914
rect 2206 41862 2258 41914
rect 6950 41862 7002 41914
rect 7014 41862 7066 41914
rect 7078 41862 7130 41914
rect 7142 41862 7194 41914
rect 7206 41862 7258 41914
rect 11950 41862 12002 41914
rect 12014 41862 12066 41914
rect 12078 41862 12130 41914
rect 12142 41862 12194 41914
rect 12206 41862 12258 41914
rect 16950 41862 17002 41914
rect 17014 41862 17066 41914
rect 17078 41862 17130 41914
rect 17142 41862 17194 41914
rect 17206 41862 17258 41914
rect 21950 41862 22002 41914
rect 22014 41862 22066 41914
rect 22078 41862 22130 41914
rect 22142 41862 22194 41914
rect 22206 41862 22258 41914
rect 26950 41862 27002 41914
rect 27014 41862 27066 41914
rect 27078 41862 27130 41914
rect 27142 41862 27194 41914
rect 27206 41862 27258 41914
rect 31950 41862 32002 41914
rect 32014 41862 32066 41914
rect 32078 41862 32130 41914
rect 32142 41862 32194 41914
rect 32206 41862 32258 41914
rect 36950 41862 37002 41914
rect 37014 41862 37066 41914
rect 37078 41862 37130 41914
rect 37142 41862 37194 41914
rect 37206 41862 37258 41914
rect 9128 41760 9180 41812
rect 9496 41760 9548 41812
rect 8944 41692 8996 41744
rect 27344 41760 27396 41812
rect 29736 41624 29788 41676
rect 15568 41556 15620 41608
rect 16488 41556 16540 41608
rect 32772 41556 32824 41608
rect 33232 41667 33284 41676
rect 33232 41633 33241 41667
rect 33241 41633 33275 41667
rect 33275 41633 33284 41667
rect 33232 41624 33284 41633
rect 34980 41556 35032 41608
rect 8484 41488 8536 41540
rect 8944 41488 8996 41540
rect 28264 41488 28316 41540
rect 32312 41488 32364 41540
rect 8760 41420 8812 41472
rect 11796 41420 11848 41472
rect 23112 41420 23164 41472
rect 23756 41420 23808 41472
rect 28356 41420 28408 41472
rect 28816 41420 28868 41472
rect 31116 41420 31168 41472
rect 33324 41420 33376 41472
rect 36636 41420 36688 41472
rect 38660 41420 38712 41472
rect 2610 41318 2662 41370
rect 2674 41318 2726 41370
rect 2738 41318 2790 41370
rect 2802 41318 2854 41370
rect 2866 41318 2918 41370
rect 7610 41318 7662 41370
rect 7674 41318 7726 41370
rect 7738 41318 7790 41370
rect 7802 41318 7854 41370
rect 7866 41318 7918 41370
rect 12610 41318 12662 41370
rect 12674 41318 12726 41370
rect 12738 41318 12790 41370
rect 12802 41318 12854 41370
rect 12866 41318 12918 41370
rect 17610 41318 17662 41370
rect 17674 41318 17726 41370
rect 17738 41318 17790 41370
rect 17802 41318 17854 41370
rect 17866 41318 17918 41370
rect 22610 41318 22662 41370
rect 22674 41318 22726 41370
rect 22738 41318 22790 41370
rect 22802 41318 22854 41370
rect 22866 41318 22918 41370
rect 27610 41318 27662 41370
rect 27674 41318 27726 41370
rect 27738 41318 27790 41370
rect 27802 41318 27854 41370
rect 27866 41318 27918 41370
rect 32610 41318 32662 41370
rect 32674 41318 32726 41370
rect 32738 41318 32790 41370
rect 32802 41318 32854 41370
rect 32866 41318 32918 41370
rect 37610 41318 37662 41370
rect 37674 41318 37726 41370
rect 37738 41318 37790 41370
rect 37802 41318 37854 41370
rect 37866 41318 37918 41370
rect 16580 41216 16632 41268
rect 17316 41216 17368 41268
rect 19984 41216 20036 41268
rect 5540 41080 5592 41132
rect 21548 41148 21600 41200
rect 17316 41080 17368 41132
rect 3424 41055 3476 41064
rect 3424 41021 3433 41055
rect 3433 41021 3467 41055
rect 3467 41021 3476 41055
rect 3424 41012 3476 41021
rect 3884 41012 3936 41064
rect 10416 41012 10468 41064
rect 29184 41148 29236 41200
rect 22836 41080 22888 41132
rect 23388 41080 23440 41132
rect 25136 41080 25188 41132
rect 25872 41123 25924 41132
rect 25872 41089 25881 41123
rect 25881 41089 25915 41123
rect 25915 41089 25924 41123
rect 25872 41080 25924 41089
rect 27988 41080 28040 41132
rect 29276 41123 29328 41132
rect 29276 41089 29285 41123
rect 29285 41089 29319 41123
rect 29319 41089 29328 41123
rect 29276 41080 29328 41089
rect 29644 41216 29696 41268
rect 29920 41216 29972 41268
rect 29920 41123 29972 41132
rect 29920 41089 29929 41123
rect 29929 41089 29963 41123
rect 29963 41089 29972 41123
rect 29920 41080 29972 41089
rect 30564 41123 30616 41132
rect 30564 41089 30573 41123
rect 30573 41089 30607 41123
rect 30607 41089 30616 41123
rect 30564 41080 30616 41089
rect 30840 41080 30892 41132
rect 22744 40944 22796 40996
rect 10600 40876 10652 40928
rect 31024 41055 31076 41064
rect 31024 41021 31033 41055
rect 31033 41021 31067 41055
rect 31067 41021 31076 41055
rect 31024 41012 31076 41021
rect 23664 40944 23716 40996
rect 29276 40944 29328 40996
rect 34060 41148 34112 41200
rect 23112 40876 23164 40928
rect 29184 40876 29236 40928
rect 30104 40876 30156 40928
rect 1950 40774 2002 40826
rect 2014 40774 2066 40826
rect 2078 40774 2130 40826
rect 2142 40774 2194 40826
rect 2206 40774 2258 40826
rect 6950 40774 7002 40826
rect 7014 40774 7066 40826
rect 7078 40774 7130 40826
rect 7142 40774 7194 40826
rect 7206 40774 7258 40826
rect 11950 40774 12002 40826
rect 12014 40774 12066 40826
rect 12078 40774 12130 40826
rect 12142 40774 12194 40826
rect 12206 40774 12258 40826
rect 16950 40774 17002 40826
rect 17014 40774 17066 40826
rect 17078 40774 17130 40826
rect 17142 40774 17194 40826
rect 17206 40774 17258 40826
rect 21950 40774 22002 40826
rect 22014 40774 22066 40826
rect 22078 40774 22130 40826
rect 22142 40774 22194 40826
rect 22206 40774 22258 40826
rect 26950 40774 27002 40826
rect 27014 40774 27066 40826
rect 27078 40774 27130 40826
rect 27142 40774 27194 40826
rect 27206 40774 27258 40826
rect 31950 40774 32002 40826
rect 32014 40774 32066 40826
rect 32078 40774 32130 40826
rect 32142 40774 32194 40826
rect 32206 40774 32258 40826
rect 36950 40774 37002 40826
rect 37014 40774 37066 40826
rect 37078 40774 37130 40826
rect 37142 40774 37194 40826
rect 37206 40774 37258 40826
rect 13268 40672 13320 40724
rect 21364 40672 21416 40724
rect 23020 40672 23072 40724
rect 10968 40604 11020 40656
rect 29368 40536 29420 40588
rect 36268 40536 36320 40588
rect 39304 40536 39356 40588
rect 1768 40468 1820 40520
rect 2964 40468 3016 40520
rect 3516 40511 3568 40520
rect 3516 40477 3525 40511
rect 3525 40477 3559 40511
rect 3559 40477 3568 40511
rect 3516 40468 3568 40477
rect 16764 40468 16816 40520
rect 22468 40468 22520 40520
rect 23112 40511 23164 40520
rect 23112 40477 23121 40511
rect 23121 40477 23155 40511
rect 23155 40477 23164 40511
rect 23112 40468 23164 40477
rect 23572 40511 23624 40520
rect 23572 40477 23581 40511
rect 23581 40477 23615 40511
rect 23615 40477 23624 40511
rect 23572 40468 23624 40477
rect 24676 40468 24728 40520
rect 25136 40511 25188 40520
rect 25136 40477 25145 40511
rect 25145 40477 25179 40511
rect 25179 40477 25188 40511
rect 25136 40468 25188 40477
rect 31852 40468 31904 40520
rect 32404 40468 32456 40520
rect 3056 40443 3108 40452
rect 3056 40409 3065 40443
rect 3065 40409 3099 40443
rect 3099 40409 3108 40443
rect 3056 40400 3108 40409
rect 24400 40400 24452 40452
rect 13544 40332 13596 40384
rect 22744 40332 22796 40384
rect 29460 40332 29512 40384
rect 38660 40375 38712 40384
rect 38660 40341 38669 40375
rect 38669 40341 38703 40375
rect 38703 40341 38712 40375
rect 38660 40332 38712 40341
rect 2610 40230 2662 40282
rect 2674 40230 2726 40282
rect 2738 40230 2790 40282
rect 2802 40230 2854 40282
rect 2866 40230 2918 40282
rect 7610 40230 7662 40282
rect 7674 40230 7726 40282
rect 7738 40230 7790 40282
rect 7802 40230 7854 40282
rect 7866 40230 7918 40282
rect 12610 40230 12662 40282
rect 12674 40230 12726 40282
rect 12738 40230 12790 40282
rect 12802 40230 12854 40282
rect 12866 40230 12918 40282
rect 17610 40230 17662 40282
rect 17674 40230 17726 40282
rect 17738 40230 17790 40282
rect 17802 40230 17854 40282
rect 17866 40230 17918 40282
rect 22610 40230 22662 40282
rect 22674 40230 22726 40282
rect 22738 40230 22790 40282
rect 22802 40230 22854 40282
rect 22866 40230 22918 40282
rect 27610 40230 27662 40282
rect 27674 40230 27726 40282
rect 27738 40230 27790 40282
rect 27802 40230 27854 40282
rect 27866 40230 27918 40282
rect 32610 40230 32662 40282
rect 32674 40230 32726 40282
rect 32738 40230 32790 40282
rect 32802 40230 32854 40282
rect 32866 40230 32918 40282
rect 37610 40230 37662 40282
rect 37674 40230 37726 40282
rect 37738 40230 37790 40282
rect 37802 40230 37854 40282
rect 37866 40230 37918 40282
rect 16488 40128 16540 40180
rect 16764 40128 16816 40180
rect 848 40060 900 40112
rect 10600 40060 10652 40112
rect 10876 40060 10928 40112
rect 17316 40060 17368 40112
rect 24860 40060 24912 40112
rect 39304 40103 39356 40112
rect 39304 40069 39313 40103
rect 39313 40069 39347 40103
rect 39347 40069 39356 40103
rect 39304 40060 39356 40069
rect 32312 39992 32364 40044
rect 40868 40060 40920 40112
rect 8300 39924 8352 39976
rect 10416 39856 10468 39908
rect 30564 39856 30616 39908
rect 2504 39788 2556 39840
rect 13452 39788 13504 39840
rect 15016 39788 15068 39840
rect 23388 39788 23440 39840
rect 23664 39788 23716 39840
rect 36728 39788 36780 39840
rect 1950 39686 2002 39738
rect 2014 39686 2066 39738
rect 2078 39686 2130 39738
rect 2142 39686 2194 39738
rect 2206 39686 2258 39738
rect 6950 39686 7002 39738
rect 7014 39686 7066 39738
rect 7078 39686 7130 39738
rect 7142 39686 7194 39738
rect 7206 39686 7258 39738
rect 11950 39686 12002 39738
rect 12014 39686 12066 39738
rect 12078 39686 12130 39738
rect 12142 39686 12194 39738
rect 12206 39686 12258 39738
rect 16950 39686 17002 39738
rect 17014 39686 17066 39738
rect 17078 39686 17130 39738
rect 17142 39686 17194 39738
rect 17206 39686 17258 39738
rect 21950 39686 22002 39738
rect 22014 39686 22066 39738
rect 22078 39686 22130 39738
rect 22142 39686 22194 39738
rect 22206 39686 22258 39738
rect 26950 39686 27002 39738
rect 27014 39686 27066 39738
rect 27078 39686 27130 39738
rect 27142 39686 27194 39738
rect 27206 39686 27258 39738
rect 31950 39686 32002 39738
rect 32014 39686 32066 39738
rect 32078 39686 32130 39738
rect 32142 39686 32194 39738
rect 32206 39686 32258 39738
rect 36950 39686 37002 39738
rect 37014 39686 37066 39738
rect 37078 39686 37130 39738
rect 37142 39686 37194 39738
rect 37206 39686 37258 39738
rect 14556 39584 14608 39636
rect 4252 39516 4304 39568
rect 14924 39516 14976 39568
rect 16304 39448 16356 39500
rect 23572 39584 23624 39636
rect 30748 39584 30800 39636
rect 23388 39516 23440 39568
rect 26240 39516 26292 39568
rect 28724 39516 28776 39568
rect 29736 39516 29788 39568
rect 33140 39516 33192 39568
rect 13268 39423 13320 39432
rect 13268 39389 13277 39423
rect 13277 39389 13311 39423
rect 13311 39389 13320 39423
rect 13268 39380 13320 39389
rect 19432 39380 19484 39432
rect 19616 39380 19668 39432
rect 19800 39380 19852 39432
rect 21456 39312 21508 39364
rect 23204 39423 23256 39432
rect 23204 39389 23213 39423
rect 23213 39389 23247 39423
rect 23247 39389 23256 39423
rect 23204 39380 23256 39389
rect 23296 39423 23348 39432
rect 23296 39389 23305 39423
rect 23305 39389 23339 39423
rect 23339 39389 23348 39423
rect 23296 39380 23348 39389
rect 23572 39380 23624 39432
rect 23664 39423 23716 39432
rect 23664 39389 23673 39423
rect 23673 39389 23707 39423
rect 23707 39389 23716 39423
rect 23664 39380 23716 39389
rect 25872 39380 25924 39432
rect 26148 39423 26200 39432
rect 26148 39389 26157 39423
rect 26157 39389 26191 39423
rect 26191 39389 26200 39423
rect 26148 39380 26200 39389
rect 22192 39244 22244 39296
rect 23020 39287 23072 39296
rect 23020 39253 23029 39287
rect 23029 39253 23063 39287
rect 23063 39253 23072 39287
rect 23020 39244 23072 39253
rect 23756 39244 23808 39296
rect 28632 39312 28684 39364
rect 30196 39380 30248 39432
rect 30748 39423 30800 39432
rect 30748 39389 30757 39423
rect 30757 39389 30791 39423
rect 30791 39389 30800 39423
rect 30748 39380 30800 39389
rect 33140 39423 33192 39432
rect 33140 39389 33149 39423
rect 33149 39389 33183 39423
rect 33183 39389 33192 39423
rect 33140 39380 33192 39389
rect 38200 39380 38252 39432
rect 32956 39312 33008 39364
rect 29920 39244 29972 39296
rect 31852 39244 31904 39296
rect 2610 39142 2662 39194
rect 2674 39142 2726 39194
rect 2738 39142 2790 39194
rect 2802 39142 2854 39194
rect 2866 39142 2918 39194
rect 7610 39142 7662 39194
rect 7674 39142 7726 39194
rect 7738 39142 7790 39194
rect 7802 39142 7854 39194
rect 7866 39142 7918 39194
rect 12610 39142 12662 39194
rect 12674 39142 12726 39194
rect 12738 39142 12790 39194
rect 12802 39142 12854 39194
rect 12866 39142 12918 39194
rect 17610 39142 17662 39194
rect 17674 39142 17726 39194
rect 17738 39142 17790 39194
rect 17802 39142 17854 39194
rect 17866 39142 17918 39194
rect 22610 39142 22662 39194
rect 22674 39142 22726 39194
rect 22738 39142 22790 39194
rect 22802 39142 22854 39194
rect 22866 39142 22918 39194
rect 27610 39142 27662 39194
rect 27674 39142 27726 39194
rect 27738 39142 27790 39194
rect 27802 39142 27854 39194
rect 27866 39142 27918 39194
rect 32610 39142 32662 39194
rect 32674 39142 32726 39194
rect 32738 39142 32790 39194
rect 32802 39142 32854 39194
rect 32866 39142 32918 39194
rect 37610 39142 37662 39194
rect 37674 39142 37726 39194
rect 37738 39142 37790 39194
rect 37802 39142 37854 39194
rect 37866 39142 37918 39194
rect 9864 39040 9916 39092
rect 16304 39040 16356 39092
rect 20444 39040 20496 39092
rect 28724 39040 28776 39092
rect 30104 39040 30156 39092
rect 33140 39040 33192 39092
rect 20444 38947 20496 38956
rect 20444 38913 20453 38947
rect 20453 38913 20487 38947
rect 20487 38913 20496 38947
rect 20444 38904 20496 38913
rect 26240 38972 26292 39024
rect 28816 38972 28868 39024
rect 28954 38972 29006 39024
rect 30472 38972 30524 39024
rect 30564 38972 30616 39024
rect 28632 38904 28684 38956
rect 29092 38904 29144 38956
rect 29184 38947 29236 38956
rect 29184 38913 29193 38947
rect 29193 38913 29227 38947
rect 29227 38913 29236 38947
rect 29184 38904 29236 38913
rect 29736 38904 29788 38956
rect 30748 38947 30800 38956
rect 30748 38913 30757 38947
rect 30757 38913 30791 38947
rect 30791 38913 30800 38947
rect 30748 38904 30800 38913
rect 30932 38947 30984 38956
rect 30932 38913 30941 38947
rect 30941 38913 30975 38947
rect 30975 38913 30984 38947
rect 30932 38904 30984 38913
rect 20352 38836 20404 38888
rect 20168 38768 20220 38820
rect 5080 38700 5132 38752
rect 10232 38700 10284 38752
rect 23388 38743 23440 38752
rect 23388 38709 23397 38743
rect 23397 38709 23431 38743
rect 23431 38709 23440 38743
rect 23388 38700 23440 38709
rect 23848 38879 23900 38888
rect 23848 38845 23857 38879
rect 23857 38845 23891 38879
rect 23891 38845 23900 38879
rect 23848 38836 23900 38845
rect 24308 38836 24360 38888
rect 24584 38768 24636 38820
rect 29000 38768 29052 38820
rect 29368 38836 29420 38888
rect 29552 38879 29604 38888
rect 29552 38845 29561 38879
rect 29561 38845 29595 38879
rect 29595 38845 29604 38879
rect 29552 38836 29604 38845
rect 29184 38768 29236 38820
rect 28816 38700 28868 38752
rect 29092 38700 29144 38752
rect 30196 38743 30248 38752
rect 30196 38709 30205 38743
rect 30205 38709 30239 38743
rect 30239 38709 30248 38743
rect 30196 38700 30248 38709
rect 32312 38743 32364 38752
rect 32312 38709 32321 38743
rect 32321 38709 32355 38743
rect 32355 38709 32364 38743
rect 32312 38700 32364 38709
rect 1950 38598 2002 38650
rect 2014 38598 2066 38650
rect 2078 38598 2130 38650
rect 2142 38598 2194 38650
rect 2206 38598 2258 38650
rect 6950 38598 7002 38650
rect 7014 38598 7066 38650
rect 7078 38598 7130 38650
rect 7142 38598 7194 38650
rect 7206 38598 7258 38650
rect 11950 38598 12002 38650
rect 12014 38598 12066 38650
rect 12078 38598 12130 38650
rect 12142 38598 12194 38650
rect 12206 38598 12258 38650
rect 16950 38598 17002 38650
rect 17014 38598 17066 38650
rect 17078 38598 17130 38650
rect 17142 38598 17194 38650
rect 17206 38598 17258 38650
rect 21950 38598 22002 38650
rect 22014 38598 22066 38650
rect 22078 38598 22130 38650
rect 22142 38598 22194 38650
rect 22206 38598 22258 38650
rect 26950 38598 27002 38650
rect 27014 38598 27066 38650
rect 27078 38598 27130 38650
rect 27142 38598 27194 38650
rect 27206 38598 27258 38650
rect 31950 38598 32002 38650
rect 32014 38598 32066 38650
rect 32078 38598 32130 38650
rect 32142 38598 32194 38650
rect 32206 38598 32258 38650
rect 36950 38598 37002 38650
rect 37014 38598 37066 38650
rect 37078 38598 37130 38650
rect 37142 38598 37194 38650
rect 37206 38598 37258 38650
rect 19524 38539 19576 38548
rect 19524 38505 19533 38539
rect 19533 38505 19567 38539
rect 19567 38505 19576 38539
rect 19524 38496 19576 38505
rect 24124 38496 24176 38548
rect 32312 38496 32364 38548
rect 33048 38496 33100 38548
rect 6460 38428 6512 38480
rect 23848 38360 23900 38412
rect 24768 38403 24820 38412
rect 24768 38369 24777 38403
rect 24777 38369 24811 38403
rect 24811 38369 24820 38403
rect 24768 38360 24820 38369
rect 19800 38335 19852 38344
rect 19800 38301 19809 38335
rect 19809 38301 19843 38335
rect 19843 38301 19852 38335
rect 19800 38292 19852 38301
rect 14832 38224 14884 38276
rect 24584 38335 24636 38344
rect 24584 38301 24593 38335
rect 24593 38301 24627 38335
rect 24627 38301 24636 38335
rect 24584 38292 24636 38301
rect 33692 38292 33744 38344
rect 25872 38224 25924 38276
rect 10324 38156 10376 38208
rect 2610 38054 2662 38106
rect 2674 38054 2726 38106
rect 2738 38054 2790 38106
rect 2802 38054 2854 38106
rect 2866 38054 2918 38106
rect 7610 38054 7662 38106
rect 7674 38054 7726 38106
rect 7738 38054 7790 38106
rect 7802 38054 7854 38106
rect 7866 38054 7918 38106
rect 12610 38054 12662 38106
rect 12674 38054 12726 38106
rect 12738 38054 12790 38106
rect 12802 38054 12854 38106
rect 12866 38054 12918 38106
rect 17610 38054 17662 38106
rect 17674 38054 17726 38106
rect 17738 38054 17790 38106
rect 17802 38054 17854 38106
rect 17866 38054 17918 38106
rect 22610 38054 22662 38106
rect 22674 38054 22726 38106
rect 22738 38054 22790 38106
rect 22802 38054 22854 38106
rect 22866 38054 22918 38106
rect 27610 38054 27662 38106
rect 27674 38054 27726 38106
rect 27738 38054 27790 38106
rect 27802 38054 27854 38106
rect 27866 38054 27918 38106
rect 32610 38054 32662 38106
rect 32674 38054 32726 38106
rect 32738 38054 32790 38106
rect 32802 38054 32854 38106
rect 32866 38054 32918 38106
rect 37610 38054 37662 38106
rect 37674 38054 37726 38106
rect 37738 38054 37790 38106
rect 37802 38054 37854 38106
rect 37866 38054 37918 38106
rect 32404 37952 32456 38004
rect 38384 37952 38436 38004
rect 11060 37884 11112 37936
rect 15292 37884 15344 37936
rect 25228 37927 25280 37936
rect 25228 37893 25237 37927
rect 25237 37893 25271 37927
rect 25271 37893 25280 37927
rect 25228 37884 25280 37893
rect 25504 37884 25556 37936
rect 35532 37884 35584 37936
rect 8300 37816 8352 37868
rect 16856 37816 16908 37868
rect 25688 37859 25740 37868
rect 25688 37825 25697 37859
rect 25697 37825 25731 37859
rect 25731 37825 25740 37859
rect 25688 37816 25740 37825
rect 25504 37748 25556 37800
rect 26792 37816 26844 37868
rect 27436 37816 27488 37868
rect 32588 37748 32640 37800
rect 18052 37680 18104 37732
rect 30472 37680 30524 37732
rect 29552 37612 29604 37664
rect 1950 37510 2002 37562
rect 2014 37510 2066 37562
rect 2078 37510 2130 37562
rect 2142 37510 2194 37562
rect 2206 37510 2258 37562
rect 6950 37510 7002 37562
rect 7014 37510 7066 37562
rect 7078 37510 7130 37562
rect 7142 37510 7194 37562
rect 7206 37510 7258 37562
rect 11950 37510 12002 37562
rect 12014 37510 12066 37562
rect 12078 37510 12130 37562
rect 12142 37510 12194 37562
rect 12206 37510 12258 37562
rect 16950 37510 17002 37562
rect 17014 37510 17066 37562
rect 17078 37510 17130 37562
rect 17142 37510 17194 37562
rect 17206 37510 17258 37562
rect 21950 37510 22002 37562
rect 22014 37510 22066 37562
rect 22078 37510 22130 37562
rect 22142 37510 22194 37562
rect 22206 37510 22258 37562
rect 26950 37510 27002 37562
rect 27014 37510 27066 37562
rect 27078 37510 27130 37562
rect 27142 37510 27194 37562
rect 27206 37510 27258 37562
rect 31950 37510 32002 37562
rect 32014 37510 32066 37562
rect 32078 37510 32130 37562
rect 32142 37510 32194 37562
rect 32206 37510 32258 37562
rect 36950 37510 37002 37562
rect 37014 37510 37066 37562
rect 37078 37510 37130 37562
rect 37142 37510 37194 37562
rect 37206 37510 37258 37562
rect 18604 37408 18656 37460
rect 28080 37408 28132 37460
rect 8392 37340 8444 37392
rect 25504 37340 25556 37392
rect 26608 37340 26660 37392
rect 28540 37340 28592 37392
rect 17408 37272 17460 37324
rect 18972 37272 19024 37324
rect 32496 37340 32548 37392
rect 16764 37068 16816 37120
rect 34704 37204 34756 37256
rect 34888 37204 34940 37256
rect 38844 37247 38896 37256
rect 38844 37213 38853 37247
rect 38853 37213 38887 37247
rect 38887 37213 38896 37247
rect 38844 37204 38896 37213
rect 39028 37247 39080 37256
rect 39028 37213 39037 37247
rect 39037 37213 39071 37247
rect 39071 37213 39080 37247
rect 39028 37204 39080 37213
rect 31208 37136 31260 37188
rect 17960 37068 18012 37120
rect 38016 37068 38068 37120
rect 2610 36966 2662 37018
rect 2674 36966 2726 37018
rect 2738 36966 2790 37018
rect 2802 36966 2854 37018
rect 2866 36966 2918 37018
rect 7610 36966 7662 37018
rect 7674 36966 7726 37018
rect 7738 36966 7790 37018
rect 7802 36966 7854 37018
rect 7866 36966 7918 37018
rect 12610 36966 12662 37018
rect 12674 36966 12726 37018
rect 12738 36966 12790 37018
rect 12802 36966 12854 37018
rect 12866 36966 12918 37018
rect 17610 36966 17662 37018
rect 17674 36966 17726 37018
rect 17738 36966 17790 37018
rect 17802 36966 17854 37018
rect 17866 36966 17918 37018
rect 22610 36966 22662 37018
rect 22674 36966 22726 37018
rect 22738 36966 22790 37018
rect 22802 36966 22854 37018
rect 22866 36966 22918 37018
rect 27610 36966 27662 37018
rect 27674 36966 27726 37018
rect 27738 36966 27790 37018
rect 27802 36966 27854 37018
rect 27866 36966 27918 37018
rect 32610 36966 32662 37018
rect 32674 36966 32726 37018
rect 32738 36966 32790 37018
rect 32802 36966 32854 37018
rect 32866 36966 32918 37018
rect 37610 36966 37662 37018
rect 37674 36966 37726 37018
rect 37738 36966 37790 37018
rect 37802 36966 37854 37018
rect 37866 36966 37918 37018
rect 26608 36796 26660 36848
rect 38108 36796 38160 36848
rect 23480 36728 23532 36780
rect 23940 36771 23992 36780
rect 23940 36737 23949 36771
rect 23949 36737 23983 36771
rect 23983 36737 23992 36771
rect 23940 36728 23992 36737
rect 30380 36728 30432 36780
rect 38016 36771 38068 36780
rect 38016 36737 38025 36771
rect 38025 36737 38059 36771
rect 38059 36737 38068 36771
rect 38016 36728 38068 36737
rect 38568 36660 38620 36712
rect 15292 36524 15344 36576
rect 18696 36524 18748 36576
rect 1950 36422 2002 36474
rect 2014 36422 2066 36474
rect 2078 36422 2130 36474
rect 2142 36422 2194 36474
rect 2206 36422 2258 36474
rect 6950 36422 7002 36474
rect 7014 36422 7066 36474
rect 7078 36422 7130 36474
rect 7142 36422 7194 36474
rect 7206 36422 7258 36474
rect 11950 36422 12002 36474
rect 12014 36422 12066 36474
rect 12078 36422 12130 36474
rect 12142 36422 12194 36474
rect 12206 36422 12258 36474
rect 16950 36422 17002 36474
rect 17014 36422 17066 36474
rect 17078 36422 17130 36474
rect 17142 36422 17194 36474
rect 17206 36422 17258 36474
rect 21950 36422 22002 36474
rect 22014 36422 22066 36474
rect 22078 36422 22130 36474
rect 22142 36422 22194 36474
rect 22206 36422 22258 36474
rect 26950 36422 27002 36474
rect 27014 36422 27066 36474
rect 27078 36422 27130 36474
rect 27142 36422 27194 36474
rect 27206 36422 27258 36474
rect 31950 36422 32002 36474
rect 32014 36422 32066 36474
rect 32078 36422 32130 36474
rect 32142 36422 32194 36474
rect 32206 36422 32258 36474
rect 36950 36422 37002 36474
rect 37014 36422 37066 36474
rect 37078 36422 37130 36474
rect 37142 36422 37194 36474
rect 37206 36422 37258 36474
rect 11704 36320 11756 36372
rect 30288 36252 30340 36304
rect 30748 36252 30800 36304
rect 9588 36116 9640 36168
rect 10968 36184 11020 36236
rect 20076 36184 20128 36236
rect 28264 36116 28316 36168
rect 35072 36159 35124 36168
rect 35072 36125 35081 36159
rect 35081 36125 35115 36159
rect 35115 36125 35124 36159
rect 35072 36116 35124 36125
rect 35256 36159 35308 36168
rect 35256 36125 35265 36159
rect 35265 36125 35299 36159
rect 35299 36125 35308 36159
rect 35256 36116 35308 36125
rect 2610 35878 2662 35930
rect 2674 35878 2726 35930
rect 2738 35878 2790 35930
rect 2802 35878 2854 35930
rect 2866 35878 2918 35930
rect 7610 35878 7662 35930
rect 7674 35878 7726 35930
rect 7738 35878 7790 35930
rect 7802 35878 7854 35930
rect 7866 35878 7918 35930
rect 12610 35878 12662 35930
rect 12674 35878 12726 35930
rect 12738 35878 12790 35930
rect 12802 35878 12854 35930
rect 12866 35878 12918 35930
rect 17610 35878 17662 35930
rect 17674 35878 17726 35930
rect 17738 35878 17790 35930
rect 17802 35878 17854 35930
rect 17866 35878 17918 35930
rect 22610 35878 22662 35930
rect 22674 35878 22726 35930
rect 22738 35878 22790 35930
rect 22802 35878 22854 35930
rect 22866 35878 22918 35930
rect 27610 35878 27662 35930
rect 27674 35878 27726 35930
rect 27738 35878 27790 35930
rect 27802 35878 27854 35930
rect 27866 35878 27918 35930
rect 32610 35878 32662 35930
rect 32674 35878 32726 35930
rect 32738 35878 32790 35930
rect 32802 35878 32854 35930
rect 32866 35878 32918 35930
rect 37610 35878 37662 35930
rect 37674 35878 37726 35930
rect 37738 35878 37790 35930
rect 37802 35878 37854 35930
rect 37866 35878 37918 35930
rect 3976 35776 4028 35828
rect 7472 35776 7524 35828
rect 7656 35776 7708 35828
rect 10232 35776 10284 35828
rect 23204 35776 23256 35828
rect 23388 35776 23440 35828
rect 9772 35708 9824 35760
rect 4160 35683 4212 35692
rect 4160 35649 4169 35683
rect 4169 35649 4203 35683
rect 4203 35649 4212 35683
rect 4160 35640 4212 35649
rect 14188 35640 14240 35692
rect 15016 35640 15068 35692
rect 16672 35708 16724 35760
rect 31760 35776 31812 35828
rect 31852 35708 31904 35760
rect 6092 35572 6144 35624
rect 16488 35572 16540 35624
rect 16856 35572 16908 35624
rect 17224 35640 17276 35692
rect 17592 35640 17644 35692
rect 24952 35640 25004 35692
rect 26148 35640 26200 35692
rect 26608 35640 26660 35692
rect 3976 35504 4028 35556
rect 16396 35504 16448 35556
rect 17684 35572 17736 35624
rect 19248 35504 19300 35556
rect 24952 35436 25004 35488
rect 29460 35572 29512 35624
rect 25136 35504 25188 35556
rect 30472 35640 30524 35692
rect 36544 35572 36596 35624
rect 30472 35436 30524 35488
rect 1950 35334 2002 35386
rect 2014 35334 2066 35386
rect 2078 35334 2130 35386
rect 2142 35334 2194 35386
rect 2206 35334 2258 35386
rect 6950 35334 7002 35386
rect 7014 35334 7066 35386
rect 7078 35334 7130 35386
rect 7142 35334 7194 35386
rect 7206 35334 7258 35386
rect 11950 35334 12002 35386
rect 12014 35334 12066 35386
rect 12078 35334 12130 35386
rect 12142 35334 12194 35386
rect 12206 35334 12258 35386
rect 16950 35334 17002 35386
rect 17014 35334 17066 35386
rect 17078 35334 17130 35386
rect 17142 35334 17194 35386
rect 17206 35334 17258 35386
rect 21950 35334 22002 35386
rect 22014 35334 22066 35386
rect 22078 35334 22130 35386
rect 22142 35334 22194 35386
rect 22206 35334 22258 35386
rect 26950 35334 27002 35386
rect 27014 35334 27066 35386
rect 27078 35334 27130 35386
rect 27142 35334 27194 35386
rect 27206 35334 27258 35386
rect 31950 35334 32002 35386
rect 32014 35334 32066 35386
rect 32078 35334 32130 35386
rect 32142 35334 32194 35386
rect 32206 35334 32258 35386
rect 36950 35334 37002 35386
rect 37014 35334 37066 35386
rect 37078 35334 37130 35386
rect 37142 35334 37194 35386
rect 37206 35334 37258 35386
rect 3792 35232 3844 35284
rect 6736 35232 6788 35284
rect 7196 35232 7248 35284
rect 9772 35232 9824 35284
rect 10508 35232 10560 35284
rect 6644 35164 6696 35216
rect 19892 35164 19944 35216
rect 6000 35096 6052 35148
rect 6460 35028 6512 35080
rect 7472 35028 7524 35080
rect 7656 35028 7708 35080
rect 9772 35071 9824 35080
rect 9772 35037 9781 35071
rect 9781 35037 9815 35071
rect 9815 35037 9824 35071
rect 9772 35028 9824 35037
rect 9864 35071 9916 35080
rect 9864 35037 9873 35071
rect 9873 35037 9907 35071
rect 9907 35037 9916 35071
rect 9864 35028 9916 35037
rect 11060 35096 11112 35148
rect 12440 35139 12492 35148
rect 12440 35105 12449 35139
rect 12449 35105 12483 35139
rect 12483 35105 12492 35139
rect 12440 35096 12492 35105
rect 10232 35071 10284 35080
rect 10232 35037 10241 35071
rect 10241 35037 10275 35071
rect 10275 35037 10284 35071
rect 10232 35028 10284 35037
rect 13084 35028 13136 35080
rect 14004 35096 14056 35148
rect 14832 35096 14884 35148
rect 16396 35096 16448 35148
rect 13544 35071 13596 35080
rect 13544 35037 13553 35071
rect 13553 35037 13587 35071
rect 13587 35037 13596 35071
rect 13544 35028 13596 35037
rect 13728 35071 13780 35080
rect 13728 35037 13737 35071
rect 13737 35037 13771 35071
rect 13771 35037 13780 35071
rect 13728 35028 13780 35037
rect 13820 35071 13872 35080
rect 13820 35037 13829 35071
rect 13829 35037 13863 35071
rect 13863 35037 13872 35071
rect 13820 35028 13872 35037
rect 16672 35139 16724 35148
rect 16672 35105 16681 35139
rect 16681 35105 16715 35139
rect 16715 35105 16724 35139
rect 16672 35096 16724 35105
rect 23112 35164 23164 35216
rect 33140 35164 33192 35216
rect 34152 35164 34204 35216
rect 38936 35164 38988 35216
rect 4068 34935 4120 34944
rect 4068 34901 4077 34935
rect 4077 34901 4111 34935
rect 4111 34901 4120 34935
rect 4068 34892 4120 34901
rect 8116 34960 8168 35012
rect 6460 34892 6512 34944
rect 17684 35028 17736 35080
rect 25872 35028 25924 35080
rect 17592 34960 17644 35012
rect 26608 34892 26660 34944
rect 35440 34960 35492 35012
rect 29644 34892 29696 34944
rect 38384 34892 38436 34944
rect 2610 34790 2662 34842
rect 2674 34790 2726 34842
rect 2738 34790 2790 34842
rect 2802 34790 2854 34842
rect 2866 34790 2918 34842
rect 7610 34790 7662 34842
rect 7674 34790 7726 34842
rect 7738 34790 7790 34842
rect 7802 34790 7854 34842
rect 7866 34790 7918 34842
rect 12610 34790 12662 34842
rect 12674 34790 12726 34842
rect 12738 34790 12790 34842
rect 12802 34790 12854 34842
rect 12866 34790 12918 34842
rect 17610 34790 17662 34842
rect 17674 34790 17726 34842
rect 17738 34790 17790 34842
rect 17802 34790 17854 34842
rect 17866 34790 17918 34842
rect 22610 34790 22662 34842
rect 22674 34790 22726 34842
rect 22738 34790 22790 34842
rect 22802 34790 22854 34842
rect 22866 34790 22918 34842
rect 27610 34790 27662 34842
rect 27674 34790 27726 34842
rect 27738 34790 27790 34842
rect 27802 34790 27854 34842
rect 27866 34790 27918 34842
rect 32610 34790 32662 34842
rect 32674 34790 32726 34842
rect 32738 34790 32790 34842
rect 32802 34790 32854 34842
rect 32866 34790 32918 34842
rect 37610 34790 37662 34842
rect 37674 34790 37726 34842
rect 37738 34790 37790 34842
rect 37802 34790 37854 34842
rect 37866 34790 37918 34842
rect 7196 34663 7248 34672
rect 7196 34629 7205 34663
rect 7205 34629 7239 34663
rect 7239 34629 7248 34663
rect 7196 34620 7248 34629
rect 7472 34620 7524 34672
rect 8116 34620 8168 34672
rect 7380 34595 7432 34604
rect 7380 34561 7389 34595
rect 7389 34561 7423 34595
rect 7423 34561 7432 34595
rect 7380 34552 7432 34561
rect 18696 34688 18748 34740
rect 23112 34688 23164 34740
rect 36728 34688 36780 34740
rect 16856 34620 16908 34672
rect 12992 34552 13044 34604
rect 13544 34552 13596 34604
rect 15568 34595 15620 34604
rect 15568 34561 15577 34595
rect 15577 34561 15611 34595
rect 15611 34561 15620 34595
rect 15568 34552 15620 34561
rect 15752 34595 15804 34604
rect 15752 34561 15761 34595
rect 15761 34561 15795 34595
rect 15795 34561 15804 34595
rect 15752 34552 15804 34561
rect 21640 34552 21692 34604
rect 21732 34552 21784 34604
rect 29920 34620 29972 34672
rect 34244 34620 34296 34672
rect 16672 34484 16724 34536
rect 33140 34484 33192 34536
rect 36176 34484 36228 34536
rect 38568 34527 38620 34536
rect 38568 34493 38577 34527
rect 38577 34493 38611 34527
rect 38611 34493 38620 34527
rect 38568 34484 38620 34493
rect 13728 34416 13780 34468
rect 19616 34416 19668 34468
rect 1950 34246 2002 34298
rect 2014 34246 2066 34298
rect 2078 34246 2130 34298
rect 2142 34246 2194 34298
rect 2206 34246 2258 34298
rect 6950 34246 7002 34298
rect 7014 34246 7066 34298
rect 7078 34246 7130 34298
rect 7142 34246 7194 34298
rect 7206 34246 7258 34298
rect 11950 34246 12002 34298
rect 12014 34246 12066 34298
rect 12078 34246 12130 34298
rect 12142 34246 12194 34298
rect 12206 34246 12258 34298
rect 16950 34246 17002 34298
rect 17014 34246 17066 34298
rect 17078 34246 17130 34298
rect 17142 34246 17194 34298
rect 17206 34246 17258 34298
rect 21950 34246 22002 34298
rect 22014 34246 22066 34298
rect 22078 34246 22130 34298
rect 22142 34246 22194 34298
rect 22206 34246 22258 34298
rect 26950 34246 27002 34298
rect 27014 34246 27066 34298
rect 27078 34246 27130 34298
rect 27142 34246 27194 34298
rect 27206 34246 27258 34298
rect 31950 34246 32002 34298
rect 32014 34246 32066 34298
rect 32078 34246 32130 34298
rect 32142 34246 32194 34298
rect 32206 34246 32258 34298
rect 36950 34246 37002 34298
rect 37014 34246 37066 34298
rect 37078 34246 37130 34298
rect 37142 34246 37194 34298
rect 37206 34246 37258 34298
rect 14740 34144 14792 34196
rect 25412 34144 25464 34196
rect 2964 34076 3016 34128
rect 5540 34076 5592 34128
rect 21824 34076 21876 34128
rect 7472 34008 7524 34060
rect 24860 34008 24912 34060
rect 1768 33940 1820 33992
rect 14924 33940 14976 33992
rect 15660 33940 15712 33992
rect 3516 33872 3568 33924
rect 11704 33872 11756 33924
rect 13268 33872 13320 33924
rect 17316 33872 17368 33924
rect 23572 33872 23624 33924
rect 24124 33872 24176 33924
rect 36452 33872 36504 33924
rect 16120 33804 16172 33856
rect 27988 33804 28040 33856
rect 2610 33702 2662 33754
rect 2674 33702 2726 33754
rect 2738 33702 2790 33754
rect 2802 33702 2854 33754
rect 2866 33702 2918 33754
rect 7610 33702 7662 33754
rect 7674 33702 7726 33754
rect 7738 33702 7790 33754
rect 7802 33702 7854 33754
rect 7866 33702 7918 33754
rect 12610 33702 12662 33754
rect 12674 33702 12726 33754
rect 12738 33702 12790 33754
rect 12802 33702 12854 33754
rect 12866 33702 12918 33754
rect 17610 33702 17662 33754
rect 17674 33702 17726 33754
rect 17738 33702 17790 33754
rect 17802 33702 17854 33754
rect 17866 33702 17918 33754
rect 22610 33702 22662 33754
rect 22674 33702 22726 33754
rect 22738 33702 22790 33754
rect 22802 33702 22854 33754
rect 22866 33702 22918 33754
rect 27610 33702 27662 33754
rect 27674 33702 27726 33754
rect 27738 33702 27790 33754
rect 27802 33702 27854 33754
rect 27866 33702 27918 33754
rect 32610 33702 32662 33754
rect 32674 33702 32726 33754
rect 32738 33702 32790 33754
rect 32802 33702 32854 33754
rect 32866 33702 32918 33754
rect 37610 33702 37662 33754
rect 37674 33702 37726 33754
rect 37738 33702 37790 33754
rect 37802 33702 37854 33754
rect 37866 33702 37918 33754
rect 7380 33600 7432 33652
rect 14832 33600 14884 33652
rect 14924 33600 14976 33652
rect 6368 33575 6420 33584
rect 6368 33541 6377 33575
rect 6377 33541 6411 33575
rect 6411 33541 6420 33575
rect 6368 33532 6420 33541
rect 13544 33464 13596 33516
rect 13728 33507 13780 33516
rect 13728 33473 13737 33507
rect 13737 33473 13771 33507
rect 13771 33473 13780 33507
rect 13728 33464 13780 33473
rect 14188 33507 14240 33516
rect 14188 33473 14197 33507
rect 14197 33473 14231 33507
rect 14231 33473 14240 33507
rect 14188 33464 14240 33473
rect 14832 33464 14884 33516
rect 17500 33600 17552 33652
rect 17316 33532 17368 33584
rect 18236 33532 18288 33584
rect 19248 33600 19300 33652
rect 19340 33532 19392 33584
rect 19892 33532 19944 33584
rect 22376 33532 22428 33584
rect 7380 33396 7432 33448
rect 8392 33396 8444 33448
rect 14280 33439 14332 33448
rect 14280 33405 14289 33439
rect 14289 33405 14323 33439
rect 14323 33405 14332 33439
rect 14280 33396 14332 33405
rect 15016 33396 15068 33448
rect 17868 33507 17920 33516
rect 17868 33473 17877 33507
rect 17877 33473 17911 33507
rect 17911 33473 17920 33507
rect 17868 33464 17920 33473
rect 24216 33532 24268 33584
rect 24860 33575 24912 33584
rect 24860 33541 24869 33575
rect 24869 33541 24903 33575
rect 24903 33541 24912 33575
rect 24860 33532 24912 33541
rect 23296 33464 23348 33516
rect 25412 33507 25464 33516
rect 25412 33473 25421 33507
rect 25421 33473 25455 33507
rect 25455 33473 25464 33507
rect 25412 33464 25464 33473
rect 25872 33464 25924 33516
rect 26148 33507 26200 33516
rect 26148 33473 26157 33507
rect 26157 33473 26191 33507
rect 26191 33473 26200 33507
rect 26148 33464 26200 33473
rect 18880 33396 18932 33448
rect 6368 33328 6420 33380
rect 12992 33328 13044 33380
rect 15752 33328 15804 33380
rect 14004 33260 14056 33312
rect 14648 33260 14700 33312
rect 14832 33260 14884 33312
rect 19984 33328 20036 33380
rect 18420 33260 18472 33312
rect 18696 33260 18748 33312
rect 1950 33158 2002 33210
rect 2014 33158 2066 33210
rect 2078 33158 2130 33210
rect 2142 33158 2194 33210
rect 2206 33158 2258 33210
rect 6950 33158 7002 33210
rect 7014 33158 7066 33210
rect 7078 33158 7130 33210
rect 7142 33158 7194 33210
rect 7206 33158 7258 33210
rect 11950 33158 12002 33210
rect 12014 33158 12066 33210
rect 12078 33158 12130 33210
rect 12142 33158 12194 33210
rect 12206 33158 12258 33210
rect 16950 33158 17002 33210
rect 17014 33158 17066 33210
rect 17078 33158 17130 33210
rect 17142 33158 17194 33210
rect 17206 33158 17258 33210
rect 21950 33158 22002 33210
rect 22014 33158 22066 33210
rect 22078 33158 22130 33210
rect 22142 33158 22194 33210
rect 22206 33158 22258 33210
rect 26950 33158 27002 33210
rect 27014 33158 27066 33210
rect 27078 33158 27130 33210
rect 27142 33158 27194 33210
rect 27206 33158 27258 33210
rect 31950 33158 32002 33210
rect 32014 33158 32066 33210
rect 32078 33158 32130 33210
rect 32142 33158 32194 33210
rect 32206 33158 32258 33210
rect 36950 33158 37002 33210
rect 37014 33158 37066 33210
rect 37078 33158 37130 33210
rect 37142 33158 37194 33210
rect 37206 33158 37258 33210
rect 4896 33056 4948 33108
rect 10232 33056 10284 33108
rect 13084 33056 13136 33108
rect 14188 33056 14240 33108
rect 24492 33056 24544 33108
rect 35992 33056 36044 33108
rect 3148 32988 3200 33040
rect 11520 32988 11572 33040
rect 13544 32988 13596 33040
rect 13728 32988 13780 33040
rect 15936 32988 15988 33040
rect 30380 32988 30432 33040
rect 31484 32988 31536 33040
rect 5724 32920 5776 32972
rect 11612 32920 11664 32972
rect 13820 32920 13872 32972
rect 18052 32920 18104 32972
rect 17408 32852 17460 32904
rect 33232 32895 33284 32904
rect 33232 32861 33241 32895
rect 33241 32861 33275 32895
rect 33275 32861 33284 32895
rect 33232 32852 33284 32861
rect 16856 32784 16908 32836
rect 36544 32852 36596 32904
rect 35992 32784 36044 32836
rect 38200 32852 38252 32904
rect 38200 32716 38252 32768
rect 2610 32614 2662 32666
rect 2674 32614 2726 32666
rect 2738 32614 2790 32666
rect 2802 32614 2854 32666
rect 2866 32614 2918 32666
rect 7610 32614 7662 32666
rect 7674 32614 7726 32666
rect 7738 32614 7790 32666
rect 7802 32614 7854 32666
rect 7866 32614 7918 32666
rect 12610 32614 12662 32666
rect 12674 32614 12726 32666
rect 12738 32614 12790 32666
rect 12802 32614 12854 32666
rect 12866 32614 12918 32666
rect 17610 32614 17662 32666
rect 17674 32614 17726 32666
rect 17738 32614 17790 32666
rect 17802 32614 17854 32666
rect 17866 32614 17918 32666
rect 22610 32614 22662 32666
rect 22674 32614 22726 32666
rect 22738 32614 22790 32666
rect 22802 32614 22854 32666
rect 22866 32614 22918 32666
rect 27610 32614 27662 32666
rect 27674 32614 27726 32666
rect 27738 32614 27790 32666
rect 27802 32614 27854 32666
rect 27866 32614 27918 32666
rect 32610 32614 32662 32666
rect 32674 32614 32726 32666
rect 32738 32614 32790 32666
rect 32802 32614 32854 32666
rect 32866 32614 32918 32666
rect 37610 32614 37662 32666
rect 37674 32614 37726 32666
rect 37738 32614 37790 32666
rect 37802 32614 37854 32666
rect 37866 32614 37918 32666
rect 9772 32512 9824 32564
rect 16028 32512 16080 32564
rect 6092 32444 6144 32496
rect 11428 32444 11480 32496
rect 16948 32444 17000 32496
rect 19064 32512 19116 32564
rect 17132 32444 17184 32496
rect 6000 32376 6052 32428
rect 6368 32419 6420 32428
rect 6368 32385 6377 32419
rect 6377 32385 6411 32419
rect 6411 32385 6420 32419
rect 6368 32376 6420 32385
rect 6644 32419 6696 32428
rect 6644 32385 6653 32419
rect 6653 32385 6687 32419
rect 6687 32385 6696 32419
rect 6644 32376 6696 32385
rect 6736 32419 6788 32428
rect 6736 32385 6745 32419
rect 6745 32385 6779 32419
rect 6779 32385 6788 32419
rect 6736 32376 6788 32385
rect 6460 32351 6512 32360
rect 6460 32317 6469 32351
rect 6469 32317 6503 32351
rect 6503 32317 6512 32351
rect 6460 32308 6512 32317
rect 19248 32308 19300 32360
rect 18972 32240 19024 32292
rect 19064 32240 19116 32292
rect 28632 32419 28684 32428
rect 28632 32385 28641 32419
rect 28641 32385 28675 32419
rect 28675 32385 28684 32419
rect 28632 32376 28684 32385
rect 28816 32419 28868 32428
rect 28816 32385 28825 32419
rect 28825 32385 28859 32419
rect 28859 32385 28868 32419
rect 28816 32376 28868 32385
rect 24308 32308 24360 32360
rect 28724 32308 28776 32360
rect 29000 32419 29052 32428
rect 29000 32385 29010 32419
rect 29010 32385 29044 32419
rect 29044 32385 29052 32419
rect 30932 32444 30984 32496
rect 29000 32376 29052 32385
rect 30472 32376 30524 32428
rect 18052 32172 18104 32224
rect 18328 32172 18380 32224
rect 1950 32070 2002 32122
rect 2014 32070 2066 32122
rect 2078 32070 2130 32122
rect 2142 32070 2194 32122
rect 2206 32070 2258 32122
rect 6950 32070 7002 32122
rect 7014 32070 7066 32122
rect 7078 32070 7130 32122
rect 7142 32070 7194 32122
rect 7206 32070 7258 32122
rect 11950 32070 12002 32122
rect 12014 32070 12066 32122
rect 12078 32070 12130 32122
rect 12142 32070 12194 32122
rect 12206 32070 12258 32122
rect 16950 32070 17002 32122
rect 17014 32070 17066 32122
rect 17078 32070 17130 32122
rect 17142 32070 17194 32122
rect 17206 32070 17258 32122
rect 21950 32070 22002 32122
rect 22014 32070 22066 32122
rect 22078 32070 22130 32122
rect 22142 32070 22194 32122
rect 22206 32070 22258 32122
rect 26950 32070 27002 32122
rect 27014 32070 27066 32122
rect 27078 32070 27130 32122
rect 27142 32070 27194 32122
rect 27206 32070 27258 32122
rect 31950 32070 32002 32122
rect 32014 32070 32066 32122
rect 32078 32070 32130 32122
rect 32142 32070 32194 32122
rect 32206 32070 32258 32122
rect 36950 32070 37002 32122
rect 37014 32070 37066 32122
rect 37078 32070 37130 32122
rect 37142 32070 37194 32122
rect 37206 32070 37258 32122
rect 18328 31968 18380 32020
rect 16396 31900 16448 31952
rect 16764 31900 16816 31952
rect 17316 31900 17368 31952
rect 7380 31832 7432 31884
rect 9312 31832 9364 31884
rect 10232 31832 10284 31884
rect 18696 31900 18748 31952
rect 19340 31900 19392 31952
rect 18880 31832 18932 31884
rect 1400 31807 1452 31816
rect 1400 31773 1409 31807
rect 1409 31773 1443 31807
rect 1443 31773 1452 31807
rect 1400 31764 1452 31773
rect 1676 31807 1728 31816
rect 1676 31773 1685 31807
rect 1685 31773 1719 31807
rect 1719 31773 1728 31807
rect 1676 31764 1728 31773
rect 9036 31807 9088 31816
rect 9036 31773 9045 31807
rect 9045 31773 9079 31807
rect 9079 31773 9088 31807
rect 9036 31764 9088 31773
rect 17408 31807 17460 31816
rect 17408 31773 17417 31807
rect 17417 31773 17451 31807
rect 17451 31773 17460 31807
rect 17408 31764 17460 31773
rect 24584 31832 24636 31884
rect 30564 31832 30616 31884
rect 27344 31764 27396 31816
rect 31116 31807 31168 31816
rect 31116 31773 31125 31807
rect 31125 31773 31159 31807
rect 31159 31773 31168 31807
rect 31116 31764 31168 31773
rect 32496 31764 32548 31816
rect 34060 31764 34112 31816
rect 7472 31628 7524 31680
rect 16856 31628 16908 31680
rect 2610 31526 2662 31578
rect 2674 31526 2726 31578
rect 2738 31526 2790 31578
rect 2802 31526 2854 31578
rect 2866 31526 2918 31578
rect 7610 31526 7662 31578
rect 7674 31526 7726 31578
rect 7738 31526 7790 31578
rect 7802 31526 7854 31578
rect 7866 31526 7918 31578
rect 12610 31526 12662 31578
rect 12674 31526 12726 31578
rect 12738 31526 12790 31578
rect 12802 31526 12854 31578
rect 12866 31526 12918 31578
rect 17610 31526 17662 31578
rect 17674 31526 17726 31578
rect 17738 31526 17790 31578
rect 17802 31526 17854 31578
rect 17866 31526 17918 31578
rect 22610 31526 22662 31578
rect 22674 31526 22726 31578
rect 22738 31526 22790 31578
rect 22802 31526 22854 31578
rect 22866 31526 22918 31578
rect 27610 31526 27662 31578
rect 27674 31526 27726 31578
rect 27738 31526 27790 31578
rect 27802 31526 27854 31578
rect 27866 31526 27918 31578
rect 32610 31526 32662 31578
rect 32674 31526 32726 31578
rect 32738 31526 32790 31578
rect 32802 31526 32854 31578
rect 32866 31526 32918 31578
rect 37610 31526 37662 31578
rect 37674 31526 37726 31578
rect 37738 31526 37790 31578
rect 37802 31526 37854 31578
rect 37866 31526 37918 31578
rect 16672 31424 16724 31476
rect 17408 31288 17460 31340
rect 18328 31288 18380 31340
rect 31576 31288 31628 31340
rect 40500 31331 40552 31340
rect 40500 31297 40509 31331
rect 40509 31297 40543 31331
rect 40543 31297 40552 31331
rect 40500 31288 40552 31297
rect 10232 31220 10284 31272
rect 24584 31220 24636 31272
rect 24768 31220 24820 31272
rect 33784 31220 33836 31272
rect 38292 31220 38344 31272
rect 8300 31152 8352 31204
rect 24952 31152 25004 31204
rect 15936 31084 15988 31136
rect 18512 31084 18564 31136
rect 31208 31084 31260 31136
rect 31392 31084 31444 31136
rect 1950 30982 2002 31034
rect 2014 30982 2066 31034
rect 2078 30982 2130 31034
rect 2142 30982 2194 31034
rect 2206 30982 2258 31034
rect 6950 30982 7002 31034
rect 7014 30982 7066 31034
rect 7078 30982 7130 31034
rect 7142 30982 7194 31034
rect 7206 30982 7258 31034
rect 11950 30982 12002 31034
rect 12014 30982 12066 31034
rect 12078 30982 12130 31034
rect 12142 30982 12194 31034
rect 12206 30982 12258 31034
rect 16950 30982 17002 31034
rect 17014 30982 17066 31034
rect 17078 30982 17130 31034
rect 17142 30982 17194 31034
rect 17206 30982 17258 31034
rect 21950 30982 22002 31034
rect 22014 30982 22066 31034
rect 22078 30982 22130 31034
rect 22142 30982 22194 31034
rect 22206 30982 22258 31034
rect 26950 30982 27002 31034
rect 27014 30982 27066 31034
rect 27078 30982 27130 31034
rect 27142 30982 27194 31034
rect 27206 30982 27258 31034
rect 31950 30982 32002 31034
rect 32014 30982 32066 31034
rect 32078 30982 32130 31034
rect 32142 30982 32194 31034
rect 32206 30982 32258 31034
rect 36950 30982 37002 31034
rect 37014 30982 37066 31034
rect 37078 30982 37130 31034
rect 37142 30982 37194 31034
rect 37206 30982 37258 31034
rect 16120 30880 16172 30932
rect 16488 30880 16540 30932
rect 17868 30880 17920 30932
rect 24768 30880 24820 30932
rect 35992 30880 36044 30932
rect 36360 30880 36412 30932
rect 36728 30812 36780 30864
rect 1860 30676 1912 30728
rect 2504 30744 2556 30796
rect 17960 30744 18012 30796
rect 18236 30744 18288 30796
rect 1492 30608 1544 30660
rect 3516 30676 3568 30728
rect 9864 30676 9916 30728
rect 27436 30676 27488 30728
rect 36820 30676 36872 30728
rect 13176 30540 13228 30592
rect 36268 30583 36320 30592
rect 36268 30549 36277 30583
rect 36277 30549 36311 30583
rect 36311 30549 36320 30583
rect 36268 30540 36320 30549
rect 36452 30583 36504 30592
rect 36452 30549 36461 30583
rect 36461 30549 36495 30583
rect 36495 30549 36504 30583
rect 36452 30540 36504 30549
rect 2610 30438 2662 30490
rect 2674 30438 2726 30490
rect 2738 30438 2790 30490
rect 2802 30438 2854 30490
rect 2866 30438 2918 30490
rect 7610 30438 7662 30490
rect 7674 30438 7726 30490
rect 7738 30438 7790 30490
rect 7802 30438 7854 30490
rect 7866 30438 7918 30490
rect 12610 30438 12662 30490
rect 12674 30438 12726 30490
rect 12738 30438 12790 30490
rect 12802 30438 12854 30490
rect 12866 30438 12918 30490
rect 17610 30438 17662 30490
rect 17674 30438 17726 30490
rect 17738 30438 17790 30490
rect 17802 30438 17854 30490
rect 17866 30438 17918 30490
rect 22610 30438 22662 30490
rect 22674 30438 22726 30490
rect 22738 30438 22790 30490
rect 22802 30438 22854 30490
rect 22866 30438 22918 30490
rect 27610 30438 27662 30490
rect 27674 30438 27726 30490
rect 27738 30438 27790 30490
rect 27802 30438 27854 30490
rect 27866 30438 27918 30490
rect 32610 30438 32662 30490
rect 32674 30438 32726 30490
rect 32738 30438 32790 30490
rect 32802 30438 32854 30490
rect 32866 30438 32918 30490
rect 37610 30438 37662 30490
rect 37674 30438 37726 30490
rect 37738 30438 37790 30490
rect 37802 30438 37854 30490
rect 37866 30438 37918 30490
rect 9128 30268 9180 30320
rect 35440 30268 35492 30320
rect 16672 30200 16724 30252
rect 33416 30200 33468 30252
rect 8852 30132 8904 30184
rect 11336 30064 11388 30116
rect 30104 30064 30156 30116
rect 30380 30175 30432 30184
rect 30380 30141 30389 30175
rect 30389 30141 30423 30175
rect 30423 30141 30432 30175
rect 30380 30132 30432 30141
rect 30472 30175 30524 30184
rect 30472 30141 30481 30175
rect 30481 30141 30515 30175
rect 30515 30141 30524 30175
rect 30472 30132 30524 30141
rect 31208 30064 31260 30116
rect 15016 29996 15068 30048
rect 36084 29996 36136 30048
rect 1950 29894 2002 29946
rect 2014 29894 2066 29946
rect 2078 29894 2130 29946
rect 2142 29894 2194 29946
rect 2206 29894 2258 29946
rect 6950 29894 7002 29946
rect 7014 29894 7066 29946
rect 7078 29894 7130 29946
rect 7142 29894 7194 29946
rect 7206 29894 7258 29946
rect 11950 29894 12002 29946
rect 12014 29894 12066 29946
rect 12078 29894 12130 29946
rect 12142 29894 12194 29946
rect 12206 29894 12258 29946
rect 16950 29894 17002 29946
rect 17014 29894 17066 29946
rect 17078 29894 17130 29946
rect 17142 29894 17194 29946
rect 17206 29894 17258 29946
rect 21950 29894 22002 29946
rect 22014 29894 22066 29946
rect 22078 29894 22130 29946
rect 22142 29894 22194 29946
rect 22206 29894 22258 29946
rect 26950 29894 27002 29946
rect 27014 29894 27066 29946
rect 27078 29894 27130 29946
rect 27142 29894 27194 29946
rect 27206 29894 27258 29946
rect 31950 29894 32002 29946
rect 32014 29894 32066 29946
rect 32078 29894 32130 29946
rect 32142 29894 32194 29946
rect 32206 29894 32258 29946
rect 36950 29894 37002 29946
rect 37014 29894 37066 29946
rect 37078 29894 37130 29946
rect 37142 29894 37194 29946
rect 37206 29894 37258 29946
rect 9220 29792 9272 29844
rect 23572 29792 23624 29844
rect 35440 29792 35492 29844
rect 36176 29792 36228 29844
rect 30932 29724 30984 29776
rect 17408 29656 17460 29708
rect 18328 29656 18380 29708
rect 20904 29699 20956 29708
rect 20904 29665 20913 29699
rect 20913 29665 20947 29699
rect 20947 29665 20956 29699
rect 20904 29656 20956 29665
rect 21640 29631 21692 29640
rect 21640 29597 21649 29631
rect 21649 29597 21683 29631
rect 21683 29597 21692 29631
rect 21640 29588 21692 29597
rect 21824 29588 21876 29640
rect 22468 29656 22520 29708
rect 26056 29656 26108 29708
rect 28632 29656 28684 29708
rect 38936 29656 38988 29708
rect 23204 29588 23256 29640
rect 31208 29588 31260 29640
rect 35440 29588 35492 29640
rect 36084 29631 36136 29640
rect 36084 29597 36093 29631
rect 36093 29597 36127 29631
rect 36127 29597 36136 29631
rect 36084 29588 36136 29597
rect 36176 29588 36228 29640
rect 16948 29520 17000 29572
rect 17868 29520 17920 29572
rect 8668 29452 8720 29504
rect 8944 29452 8996 29504
rect 15844 29452 15896 29504
rect 25596 29520 25648 29572
rect 27436 29520 27488 29572
rect 32496 29520 32548 29572
rect 23296 29452 23348 29504
rect 31944 29452 31996 29504
rect 2610 29350 2662 29402
rect 2674 29350 2726 29402
rect 2738 29350 2790 29402
rect 2802 29350 2854 29402
rect 2866 29350 2918 29402
rect 7610 29350 7662 29402
rect 7674 29350 7726 29402
rect 7738 29350 7790 29402
rect 7802 29350 7854 29402
rect 7866 29350 7918 29402
rect 12610 29350 12662 29402
rect 12674 29350 12726 29402
rect 12738 29350 12790 29402
rect 12802 29350 12854 29402
rect 12866 29350 12918 29402
rect 17610 29350 17662 29402
rect 17674 29350 17726 29402
rect 17738 29350 17790 29402
rect 17802 29350 17854 29402
rect 17866 29350 17918 29402
rect 22610 29350 22662 29402
rect 22674 29350 22726 29402
rect 22738 29350 22790 29402
rect 22802 29350 22854 29402
rect 22866 29350 22918 29402
rect 27610 29350 27662 29402
rect 27674 29350 27726 29402
rect 27738 29350 27790 29402
rect 27802 29350 27854 29402
rect 27866 29350 27918 29402
rect 32610 29350 32662 29402
rect 32674 29350 32726 29402
rect 32738 29350 32790 29402
rect 32802 29350 32854 29402
rect 32866 29350 32918 29402
rect 37610 29350 37662 29402
rect 37674 29350 37726 29402
rect 37738 29350 37790 29402
rect 37802 29350 37854 29402
rect 37866 29350 37918 29402
rect 8852 29112 8904 29164
rect 12256 29248 12308 29300
rect 23572 29248 23624 29300
rect 24492 29248 24544 29300
rect 36176 29248 36228 29300
rect 38936 29291 38988 29300
rect 38936 29257 38945 29291
rect 38945 29257 38979 29291
rect 38979 29257 38988 29291
rect 38936 29248 38988 29257
rect 12532 29180 12584 29232
rect 31668 29180 31720 29232
rect 11980 29155 12032 29164
rect 4712 29044 4764 29096
rect 6828 29044 6880 29096
rect 11980 29121 11989 29155
rect 11989 29121 12023 29155
rect 12023 29121 12032 29155
rect 11980 29112 12032 29121
rect 12256 29112 12308 29164
rect 17408 29112 17460 29164
rect 30932 29112 30984 29164
rect 10600 29044 10652 29096
rect 11336 29087 11388 29096
rect 11336 29053 11345 29087
rect 11345 29053 11379 29087
rect 11379 29053 11388 29087
rect 11336 29044 11388 29053
rect 16304 29044 16356 29096
rect 16948 29044 17000 29096
rect 30104 29044 30156 29096
rect 11520 28976 11572 29028
rect 11796 29019 11848 29028
rect 11796 28985 11805 29019
rect 11805 28985 11839 29019
rect 11839 28985 11848 29019
rect 11796 28976 11848 28985
rect 11980 28976 12032 29028
rect 12532 28976 12584 29028
rect 16672 28976 16724 29028
rect 17868 28976 17920 29028
rect 33232 28976 33284 29028
rect 33968 28976 34020 29028
rect 9128 28951 9180 28960
rect 9128 28917 9137 28951
rect 9137 28917 9171 28951
rect 9171 28917 9180 28951
rect 9128 28908 9180 28917
rect 9680 28908 9732 28960
rect 10048 28908 10100 28960
rect 17776 28908 17828 28960
rect 25320 28908 25372 28960
rect 25964 28908 26016 28960
rect 1950 28806 2002 28858
rect 2014 28806 2066 28858
rect 2078 28806 2130 28858
rect 2142 28806 2194 28858
rect 2206 28806 2258 28858
rect 6950 28806 7002 28858
rect 7014 28806 7066 28858
rect 7078 28806 7130 28858
rect 7142 28806 7194 28858
rect 7206 28806 7258 28858
rect 11950 28806 12002 28858
rect 12014 28806 12066 28858
rect 12078 28806 12130 28858
rect 12142 28806 12194 28858
rect 12206 28806 12258 28858
rect 16950 28806 17002 28858
rect 17014 28806 17066 28858
rect 17078 28806 17130 28858
rect 17142 28806 17194 28858
rect 17206 28806 17258 28858
rect 21950 28806 22002 28858
rect 22014 28806 22066 28858
rect 22078 28806 22130 28858
rect 22142 28806 22194 28858
rect 22206 28806 22258 28858
rect 26950 28806 27002 28858
rect 27014 28806 27066 28858
rect 27078 28806 27130 28858
rect 27142 28806 27194 28858
rect 27206 28806 27258 28858
rect 31950 28806 32002 28858
rect 32014 28806 32066 28858
rect 32078 28806 32130 28858
rect 32142 28806 32194 28858
rect 32206 28806 32258 28858
rect 36950 28806 37002 28858
rect 37014 28806 37066 28858
rect 37078 28806 37130 28858
rect 37142 28806 37194 28858
rect 37206 28806 37258 28858
rect 16856 28704 16908 28756
rect 16948 28704 17000 28756
rect 18696 28704 18748 28756
rect 23940 28704 23992 28756
rect 10784 28543 10836 28552
rect 10784 28509 10793 28543
rect 10793 28509 10827 28543
rect 10827 28509 10836 28543
rect 10784 28500 10836 28509
rect 17408 28611 17460 28620
rect 17408 28577 17417 28611
rect 17417 28577 17451 28611
rect 17451 28577 17460 28611
rect 17408 28568 17460 28577
rect 17776 28611 17828 28620
rect 17776 28577 17785 28611
rect 17785 28577 17819 28611
rect 17819 28577 17828 28611
rect 17776 28568 17828 28577
rect 24400 28568 24452 28620
rect 15936 28500 15988 28552
rect 10692 28432 10744 28484
rect 16948 28500 17000 28552
rect 16672 28432 16724 28484
rect 20720 28500 20772 28552
rect 25320 28432 25372 28484
rect 19800 28364 19852 28416
rect 2610 28262 2662 28314
rect 2674 28262 2726 28314
rect 2738 28262 2790 28314
rect 2802 28262 2854 28314
rect 2866 28262 2918 28314
rect 7610 28262 7662 28314
rect 7674 28262 7726 28314
rect 7738 28262 7790 28314
rect 7802 28262 7854 28314
rect 7866 28262 7918 28314
rect 12610 28262 12662 28314
rect 12674 28262 12726 28314
rect 12738 28262 12790 28314
rect 12802 28262 12854 28314
rect 12866 28262 12918 28314
rect 17610 28262 17662 28314
rect 17674 28262 17726 28314
rect 17738 28262 17790 28314
rect 17802 28262 17854 28314
rect 17866 28262 17918 28314
rect 22610 28262 22662 28314
rect 22674 28262 22726 28314
rect 22738 28262 22790 28314
rect 22802 28262 22854 28314
rect 22866 28262 22918 28314
rect 27610 28262 27662 28314
rect 27674 28262 27726 28314
rect 27738 28262 27790 28314
rect 27802 28262 27854 28314
rect 27866 28262 27918 28314
rect 32610 28262 32662 28314
rect 32674 28262 32726 28314
rect 32738 28262 32790 28314
rect 32802 28262 32854 28314
rect 32866 28262 32918 28314
rect 37610 28262 37662 28314
rect 37674 28262 37726 28314
rect 37738 28262 37790 28314
rect 37802 28262 37854 28314
rect 37866 28262 37918 28314
rect 16948 28160 17000 28212
rect 17408 28160 17460 28212
rect 24860 28203 24912 28212
rect 24860 28169 24869 28203
rect 24869 28169 24903 28203
rect 24903 28169 24912 28203
rect 24860 28160 24912 28169
rect 5540 28092 5592 28144
rect 24400 28067 24452 28076
rect 24400 28033 24409 28067
rect 24409 28033 24443 28067
rect 24443 28033 24452 28067
rect 24400 28024 24452 28033
rect 24676 28067 24728 28076
rect 24676 28033 24685 28067
rect 24685 28033 24719 28067
rect 24719 28033 24728 28067
rect 24676 28024 24728 28033
rect 30932 28024 30984 28076
rect 11704 27956 11756 28008
rect 22376 27888 22428 27940
rect 20812 27820 20864 27872
rect 21548 27820 21600 27872
rect 32956 27820 33008 27872
rect 35992 27820 36044 27872
rect 1950 27718 2002 27770
rect 2014 27718 2066 27770
rect 2078 27718 2130 27770
rect 2142 27718 2194 27770
rect 2206 27718 2258 27770
rect 6950 27718 7002 27770
rect 7014 27718 7066 27770
rect 7078 27718 7130 27770
rect 7142 27718 7194 27770
rect 7206 27718 7258 27770
rect 11950 27718 12002 27770
rect 12014 27718 12066 27770
rect 12078 27718 12130 27770
rect 12142 27718 12194 27770
rect 12206 27718 12258 27770
rect 16950 27718 17002 27770
rect 17014 27718 17066 27770
rect 17078 27718 17130 27770
rect 17142 27718 17194 27770
rect 17206 27718 17258 27770
rect 21950 27718 22002 27770
rect 22014 27718 22066 27770
rect 22078 27718 22130 27770
rect 22142 27718 22194 27770
rect 22206 27718 22258 27770
rect 26950 27718 27002 27770
rect 27014 27718 27066 27770
rect 27078 27718 27130 27770
rect 27142 27718 27194 27770
rect 27206 27718 27258 27770
rect 31950 27718 32002 27770
rect 32014 27718 32066 27770
rect 32078 27718 32130 27770
rect 32142 27718 32194 27770
rect 32206 27718 32258 27770
rect 36950 27718 37002 27770
rect 37014 27718 37066 27770
rect 37078 27718 37130 27770
rect 37142 27718 37194 27770
rect 37206 27718 37258 27770
rect 17224 27616 17276 27668
rect 17408 27616 17460 27668
rect 19800 27616 19852 27668
rect 20628 27616 20680 27668
rect 34520 27616 34572 27668
rect 23296 27548 23348 27600
rect 24216 27548 24268 27600
rect 33416 27480 33468 27532
rect 32496 27412 32548 27464
rect 30380 27344 30432 27396
rect 2610 27174 2662 27226
rect 2674 27174 2726 27226
rect 2738 27174 2790 27226
rect 2802 27174 2854 27226
rect 2866 27174 2918 27226
rect 7610 27174 7662 27226
rect 7674 27174 7726 27226
rect 7738 27174 7790 27226
rect 7802 27174 7854 27226
rect 7866 27174 7918 27226
rect 12610 27174 12662 27226
rect 12674 27174 12726 27226
rect 12738 27174 12790 27226
rect 12802 27174 12854 27226
rect 12866 27174 12918 27226
rect 17610 27174 17662 27226
rect 17674 27174 17726 27226
rect 17738 27174 17790 27226
rect 17802 27174 17854 27226
rect 17866 27174 17918 27226
rect 22610 27174 22662 27226
rect 22674 27174 22726 27226
rect 22738 27174 22790 27226
rect 22802 27174 22854 27226
rect 22866 27174 22918 27226
rect 27610 27174 27662 27226
rect 27674 27174 27726 27226
rect 27738 27174 27790 27226
rect 27802 27174 27854 27226
rect 27866 27174 27918 27226
rect 32610 27174 32662 27226
rect 32674 27174 32726 27226
rect 32738 27174 32790 27226
rect 32802 27174 32854 27226
rect 32866 27174 32918 27226
rect 37610 27174 37662 27226
rect 37674 27174 37726 27226
rect 37738 27174 37790 27226
rect 37802 27174 37854 27226
rect 37866 27174 37918 27226
rect 16580 27004 16632 27056
rect 17408 27004 17460 27056
rect 13912 26936 13964 26988
rect 4068 26800 4120 26852
rect 17592 26800 17644 26852
rect 18604 26868 18656 26920
rect 19156 26868 19208 26920
rect 23112 26868 23164 26920
rect 33416 26868 33468 26920
rect 38568 26868 38620 26920
rect 26516 26800 26568 26852
rect 1950 26630 2002 26682
rect 2014 26630 2066 26682
rect 2078 26630 2130 26682
rect 2142 26630 2194 26682
rect 2206 26630 2258 26682
rect 6950 26630 7002 26682
rect 7014 26630 7066 26682
rect 7078 26630 7130 26682
rect 7142 26630 7194 26682
rect 7206 26630 7258 26682
rect 11950 26630 12002 26682
rect 12014 26630 12066 26682
rect 12078 26630 12130 26682
rect 12142 26630 12194 26682
rect 12206 26630 12258 26682
rect 16950 26630 17002 26682
rect 17014 26630 17066 26682
rect 17078 26630 17130 26682
rect 17142 26630 17194 26682
rect 17206 26630 17258 26682
rect 21950 26630 22002 26682
rect 22014 26630 22066 26682
rect 22078 26630 22130 26682
rect 22142 26630 22194 26682
rect 22206 26630 22258 26682
rect 26950 26630 27002 26682
rect 27014 26630 27066 26682
rect 27078 26630 27130 26682
rect 27142 26630 27194 26682
rect 27206 26630 27258 26682
rect 31950 26630 32002 26682
rect 32014 26630 32066 26682
rect 32078 26630 32130 26682
rect 32142 26630 32194 26682
rect 32206 26630 32258 26682
rect 36950 26630 37002 26682
rect 37014 26630 37066 26682
rect 37078 26630 37130 26682
rect 37142 26630 37194 26682
rect 37206 26630 37258 26682
rect 24952 26460 25004 26512
rect 9588 26392 9640 26444
rect 16396 26392 16448 26444
rect 19248 26392 19300 26444
rect 4712 26324 4764 26376
rect 17224 26324 17276 26376
rect 17592 26324 17644 26376
rect 36636 26528 36688 26580
rect 9680 26256 9732 26308
rect 15200 26256 15252 26308
rect 31760 26367 31812 26376
rect 31760 26333 31770 26367
rect 31770 26333 31804 26367
rect 31804 26333 31812 26367
rect 31760 26324 31812 26333
rect 6276 26188 6328 26240
rect 6460 26188 6512 26240
rect 31760 26188 31812 26240
rect 37372 26188 37424 26240
rect 37556 26188 37608 26240
rect 2610 26086 2662 26138
rect 2674 26086 2726 26138
rect 2738 26086 2790 26138
rect 2802 26086 2854 26138
rect 2866 26086 2918 26138
rect 7610 26086 7662 26138
rect 7674 26086 7726 26138
rect 7738 26086 7790 26138
rect 7802 26086 7854 26138
rect 7866 26086 7918 26138
rect 12610 26086 12662 26138
rect 12674 26086 12726 26138
rect 12738 26086 12790 26138
rect 12802 26086 12854 26138
rect 12866 26086 12918 26138
rect 17610 26086 17662 26138
rect 17674 26086 17726 26138
rect 17738 26086 17790 26138
rect 17802 26086 17854 26138
rect 17866 26086 17918 26138
rect 22610 26086 22662 26138
rect 22674 26086 22726 26138
rect 22738 26086 22790 26138
rect 22802 26086 22854 26138
rect 22866 26086 22918 26138
rect 27610 26086 27662 26138
rect 27674 26086 27726 26138
rect 27738 26086 27790 26138
rect 27802 26086 27854 26138
rect 27866 26086 27918 26138
rect 32610 26086 32662 26138
rect 32674 26086 32726 26138
rect 32738 26086 32790 26138
rect 32802 26086 32854 26138
rect 32866 26086 32918 26138
rect 37610 26086 37662 26138
rect 37674 26086 37726 26138
rect 37738 26086 37790 26138
rect 37802 26086 37854 26138
rect 37866 26086 37918 26138
rect 6460 25984 6512 26036
rect 1676 25916 1728 25968
rect 2412 25916 2464 25968
rect 5908 25848 5960 25900
rect 6644 25891 6696 25900
rect 6644 25857 6653 25891
rect 6653 25857 6687 25891
rect 6687 25857 6696 25891
rect 6644 25848 6696 25857
rect 7472 25916 7524 25968
rect 8392 25916 8444 25968
rect 5540 25780 5592 25832
rect 9036 25848 9088 25900
rect 17500 25984 17552 26036
rect 18052 25959 18104 25968
rect 18052 25925 18061 25959
rect 18061 25925 18095 25959
rect 18095 25925 18104 25959
rect 18052 25916 18104 25925
rect 25320 25916 25372 25968
rect 25136 25848 25188 25900
rect 11060 25780 11112 25832
rect 17224 25780 17276 25832
rect 17408 25780 17460 25832
rect 18972 25780 19024 25832
rect 31024 25780 31076 25832
rect 16856 25712 16908 25764
rect 24308 25712 24360 25764
rect 38936 25712 38988 25764
rect 15660 25644 15712 25696
rect 26056 25644 26108 25696
rect 1950 25542 2002 25594
rect 2014 25542 2066 25594
rect 2078 25542 2130 25594
rect 2142 25542 2194 25594
rect 2206 25542 2258 25594
rect 6950 25542 7002 25594
rect 7014 25542 7066 25594
rect 7078 25542 7130 25594
rect 7142 25542 7194 25594
rect 7206 25542 7258 25594
rect 11950 25542 12002 25594
rect 12014 25542 12066 25594
rect 12078 25542 12130 25594
rect 12142 25542 12194 25594
rect 12206 25542 12258 25594
rect 16950 25542 17002 25594
rect 17014 25542 17066 25594
rect 17078 25542 17130 25594
rect 17142 25542 17194 25594
rect 17206 25542 17258 25594
rect 21950 25542 22002 25594
rect 22014 25542 22066 25594
rect 22078 25542 22130 25594
rect 22142 25542 22194 25594
rect 22206 25542 22258 25594
rect 26950 25542 27002 25594
rect 27014 25542 27066 25594
rect 27078 25542 27130 25594
rect 27142 25542 27194 25594
rect 27206 25542 27258 25594
rect 31950 25542 32002 25594
rect 32014 25542 32066 25594
rect 32078 25542 32130 25594
rect 32142 25542 32194 25594
rect 32206 25542 32258 25594
rect 36950 25542 37002 25594
rect 37014 25542 37066 25594
rect 37078 25542 37130 25594
rect 37142 25542 37194 25594
rect 37206 25542 37258 25594
rect 16304 25440 16356 25492
rect 16856 25440 16908 25492
rect 15936 25372 15988 25424
rect 34060 25372 34112 25424
rect 17316 25304 17368 25356
rect 38200 25304 38252 25356
rect 10692 25236 10744 25288
rect 38384 25279 38436 25288
rect 38384 25245 38393 25279
rect 38393 25245 38427 25279
rect 38427 25245 38436 25279
rect 38384 25236 38436 25245
rect 17316 25168 17368 25220
rect 17868 25168 17920 25220
rect 31484 25168 31536 25220
rect 19524 25100 19576 25152
rect 2610 24998 2662 25050
rect 2674 24998 2726 25050
rect 2738 24998 2790 25050
rect 2802 24998 2854 25050
rect 2866 24998 2918 25050
rect 7610 24998 7662 25050
rect 7674 24998 7726 25050
rect 7738 24998 7790 25050
rect 7802 24998 7854 25050
rect 7866 24998 7918 25050
rect 12610 24998 12662 25050
rect 12674 24998 12726 25050
rect 12738 24998 12790 25050
rect 12802 24998 12854 25050
rect 12866 24998 12918 25050
rect 17610 24998 17662 25050
rect 17674 24998 17726 25050
rect 17738 24998 17790 25050
rect 17802 24998 17854 25050
rect 17866 24998 17918 25050
rect 22610 24998 22662 25050
rect 22674 24998 22726 25050
rect 22738 24998 22790 25050
rect 22802 24998 22854 25050
rect 22866 24998 22918 25050
rect 27610 24998 27662 25050
rect 27674 24998 27726 25050
rect 27738 24998 27790 25050
rect 27802 24998 27854 25050
rect 27866 24998 27918 25050
rect 32610 24998 32662 25050
rect 32674 24998 32726 25050
rect 32738 24998 32790 25050
rect 32802 24998 32854 25050
rect 32866 24998 32918 25050
rect 37610 24998 37662 25050
rect 37674 24998 37726 25050
rect 37738 24998 37790 25050
rect 37802 24998 37854 25050
rect 37866 24998 37918 25050
rect 27528 24896 27580 24948
rect 3424 24760 3476 24812
rect 5172 24760 5224 24812
rect 8024 24760 8076 24812
rect 10508 24803 10560 24812
rect 10508 24769 10517 24803
rect 10517 24769 10551 24803
rect 10551 24769 10560 24803
rect 10508 24760 10560 24769
rect 7288 24692 7340 24744
rect 7472 24692 7524 24744
rect 10416 24667 10468 24676
rect 10416 24633 10425 24667
rect 10425 24633 10459 24667
rect 10459 24633 10468 24667
rect 10416 24624 10468 24633
rect 18604 24760 18656 24812
rect 19984 24803 20036 24812
rect 19984 24769 19993 24803
rect 19993 24769 20027 24803
rect 20027 24769 20036 24803
rect 19984 24760 20036 24769
rect 20536 24760 20588 24812
rect 26332 24760 26384 24812
rect 27436 24760 27488 24812
rect 20720 24692 20772 24744
rect 22376 24624 22428 24676
rect 7288 24556 7340 24608
rect 19984 24556 20036 24608
rect 27344 24556 27396 24608
rect 38568 24760 38620 24812
rect 39212 24760 39264 24812
rect 27620 24692 27672 24744
rect 38292 24692 38344 24744
rect 1950 24454 2002 24506
rect 2014 24454 2066 24506
rect 2078 24454 2130 24506
rect 2142 24454 2194 24506
rect 2206 24454 2258 24506
rect 6950 24454 7002 24506
rect 7014 24454 7066 24506
rect 7078 24454 7130 24506
rect 7142 24454 7194 24506
rect 7206 24454 7258 24506
rect 11950 24454 12002 24506
rect 12014 24454 12066 24506
rect 12078 24454 12130 24506
rect 12142 24454 12194 24506
rect 12206 24454 12258 24506
rect 16950 24454 17002 24506
rect 17014 24454 17066 24506
rect 17078 24454 17130 24506
rect 17142 24454 17194 24506
rect 17206 24454 17258 24506
rect 21950 24454 22002 24506
rect 22014 24454 22066 24506
rect 22078 24454 22130 24506
rect 22142 24454 22194 24506
rect 22206 24454 22258 24506
rect 26950 24454 27002 24506
rect 27014 24454 27066 24506
rect 27078 24454 27130 24506
rect 27142 24454 27194 24506
rect 27206 24454 27258 24506
rect 31950 24454 32002 24506
rect 32014 24454 32066 24506
rect 32078 24454 32130 24506
rect 32142 24454 32194 24506
rect 32206 24454 32258 24506
rect 36950 24454 37002 24506
rect 37014 24454 37066 24506
rect 37078 24454 37130 24506
rect 37142 24454 37194 24506
rect 37206 24454 37258 24506
rect 8116 24352 8168 24404
rect 8300 24352 8352 24404
rect 10508 24352 10560 24404
rect 24676 24352 24728 24404
rect 36360 24352 36412 24404
rect 1676 24284 1728 24336
rect 4988 24284 5040 24336
rect 1768 24216 1820 24268
rect 10968 24216 11020 24268
rect 18972 24259 19024 24268
rect 18972 24225 18981 24259
rect 18981 24225 19015 24259
rect 19015 24225 19024 24259
rect 18972 24216 19024 24225
rect 7472 24148 7524 24200
rect 12348 24148 12400 24200
rect 18144 24191 18196 24200
rect 18144 24157 18153 24191
rect 18153 24157 18187 24191
rect 18187 24157 18196 24191
rect 18144 24148 18196 24157
rect 18696 24191 18748 24200
rect 18696 24157 18705 24191
rect 18705 24157 18739 24191
rect 18739 24157 18748 24191
rect 18696 24148 18748 24157
rect 23296 24148 23348 24200
rect 33048 24148 33100 24200
rect 33416 24191 33468 24200
rect 33416 24157 33425 24191
rect 33425 24157 33459 24191
rect 33459 24157 33468 24191
rect 33416 24148 33468 24157
rect 34244 24148 34296 24200
rect 8024 24123 8076 24132
rect 8024 24089 8033 24123
rect 8033 24089 8067 24123
rect 8067 24089 8076 24123
rect 8024 24080 8076 24089
rect 26056 24123 26108 24132
rect 26056 24089 26065 24123
rect 26065 24089 26099 24123
rect 26099 24089 26108 24123
rect 26056 24080 26108 24089
rect 26148 24080 26200 24132
rect 29644 24080 29696 24132
rect 36544 24080 36596 24132
rect 19156 24012 19208 24064
rect 26332 24055 26384 24064
rect 26332 24021 26341 24055
rect 26341 24021 26375 24055
rect 26375 24021 26384 24055
rect 26332 24012 26384 24021
rect 26516 24055 26568 24064
rect 26516 24021 26525 24055
rect 26525 24021 26559 24055
rect 26559 24021 26568 24055
rect 26516 24012 26568 24021
rect 2610 23910 2662 23962
rect 2674 23910 2726 23962
rect 2738 23910 2790 23962
rect 2802 23910 2854 23962
rect 2866 23910 2918 23962
rect 7610 23910 7662 23962
rect 7674 23910 7726 23962
rect 7738 23910 7790 23962
rect 7802 23910 7854 23962
rect 7866 23910 7918 23962
rect 12610 23910 12662 23962
rect 12674 23910 12726 23962
rect 12738 23910 12790 23962
rect 12802 23910 12854 23962
rect 12866 23910 12918 23962
rect 17610 23910 17662 23962
rect 17674 23910 17726 23962
rect 17738 23910 17790 23962
rect 17802 23910 17854 23962
rect 17866 23910 17918 23962
rect 22610 23910 22662 23962
rect 22674 23910 22726 23962
rect 22738 23910 22790 23962
rect 22802 23910 22854 23962
rect 22866 23910 22918 23962
rect 27610 23910 27662 23962
rect 27674 23910 27726 23962
rect 27738 23910 27790 23962
rect 27802 23910 27854 23962
rect 27866 23910 27918 23962
rect 32610 23910 32662 23962
rect 32674 23910 32726 23962
rect 32738 23910 32790 23962
rect 32802 23910 32854 23962
rect 32866 23910 32918 23962
rect 37610 23910 37662 23962
rect 37674 23910 37726 23962
rect 37738 23910 37790 23962
rect 37802 23910 37854 23962
rect 37866 23910 37918 23962
rect 8300 23808 8352 23860
rect 25872 23808 25924 23860
rect 26148 23808 26200 23860
rect 26332 23808 26384 23860
rect 7472 23740 7524 23792
rect 8116 23740 8168 23792
rect 35440 23740 35492 23792
rect 8300 23604 8352 23656
rect 24584 23672 24636 23724
rect 34244 23715 34296 23724
rect 34244 23681 34253 23715
rect 34253 23681 34287 23715
rect 34287 23681 34296 23715
rect 34244 23672 34296 23681
rect 27528 23604 27580 23656
rect 33048 23604 33100 23656
rect 34152 23647 34204 23656
rect 34152 23613 34161 23647
rect 34161 23613 34195 23647
rect 34195 23613 34204 23647
rect 34152 23604 34204 23613
rect 26332 23536 26384 23588
rect 33784 23536 33836 23588
rect 8484 23468 8536 23520
rect 1950 23366 2002 23418
rect 2014 23366 2066 23418
rect 2078 23366 2130 23418
rect 2142 23366 2194 23418
rect 2206 23366 2258 23418
rect 6950 23366 7002 23418
rect 7014 23366 7066 23418
rect 7078 23366 7130 23418
rect 7142 23366 7194 23418
rect 7206 23366 7258 23418
rect 11950 23366 12002 23418
rect 12014 23366 12066 23418
rect 12078 23366 12130 23418
rect 12142 23366 12194 23418
rect 12206 23366 12258 23418
rect 16950 23366 17002 23418
rect 17014 23366 17066 23418
rect 17078 23366 17130 23418
rect 17142 23366 17194 23418
rect 17206 23366 17258 23418
rect 21950 23366 22002 23418
rect 22014 23366 22066 23418
rect 22078 23366 22130 23418
rect 22142 23366 22194 23418
rect 22206 23366 22258 23418
rect 26950 23366 27002 23418
rect 27014 23366 27066 23418
rect 27078 23366 27130 23418
rect 27142 23366 27194 23418
rect 27206 23366 27258 23418
rect 31950 23366 32002 23418
rect 32014 23366 32066 23418
rect 32078 23366 32130 23418
rect 32142 23366 32194 23418
rect 32206 23366 32258 23418
rect 36950 23366 37002 23418
rect 37014 23366 37066 23418
rect 37078 23366 37130 23418
rect 37142 23366 37194 23418
rect 37206 23366 37258 23418
rect 3608 23264 3660 23316
rect 3976 23264 4028 23316
rect 6828 23196 6880 23248
rect 17316 23264 17368 23316
rect 18328 23264 18380 23316
rect 21732 23264 21784 23316
rect 8944 23196 8996 23248
rect 11704 23196 11756 23248
rect 12256 23196 12308 23248
rect 10324 23128 10376 23180
rect 15016 23128 15068 23180
rect 27436 23128 27488 23180
rect 17960 23060 18012 23112
rect 18236 23060 18288 23112
rect 19892 22992 19944 23044
rect 30380 22992 30432 23044
rect 4988 22924 5040 22976
rect 8668 22924 8720 22976
rect 8944 22924 8996 22976
rect 18236 22924 18288 22976
rect 37372 22924 37424 22976
rect 2610 22822 2662 22874
rect 2674 22822 2726 22874
rect 2738 22822 2790 22874
rect 2802 22822 2854 22874
rect 2866 22822 2918 22874
rect 7610 22822 7662 22874
rect 7674 22822 7726 22874
rect 7738 22822 7790 22874
rect 7802 22822 7854 22874
rect 7866 22822 7918 22874
rect 12610 22822 12662 22874
rect 12674 22822 12726 22874
rect 12738 22822 12790 22874
rect 12802 22822 12854 22874
rect 12866 22822 12918 22874
rect 17610 22822 17662 22874
rect 17674 22822 17726 22874
rect 17738 22822 17790 22874
rect 17802 22822 17854 22874
rect 17866 22822 17918 22874
rect 22610 22822 22662 22874
rect 22674 22822 22726 22874
rect 22738 22822 22790 22874
rect 22802 22822 22854 22874
rect 22866 22822 22918 22874
rect 27610 22822 27662 22874
rect 27674 22822 27726 22874
rect 27738 22822 27790 22874
rect 27802 22822 27854 22874
rect 27866 22822 27918 22874
rect 32610 22822 32662 22874
rect 32674 22822 32726 22874
rect 32738 22822 32790 22874
rect 32802 22822 32854 22874
rect 32866 22822 32918 22874
rect 37610 22822 37662 22874
rect 37674 22822 37726 22874
rect 37738 22822 37790 22874
rect 37802 22822 37854 22874
rect 37866 22822 37918 22874
rect 11612 22720 11664 22772
rect 11980 22720 12032 22772
rect 8668 22652 8720 22704
rect 11060 22652 11112 22704
rect 12256 22695 12308 22704
rect 12256 22661 12265 22695
rect 12265 22661 12299 22695
rect 12299 22661 12308 22695
rect 12256 22652 12308 22661
rect 848 22584 900 22636
rect 14924 22695 14976 22704
rect 14924 22661 14933 22695
rect 14933 22661 14967 22695
rect 14967 22661 14976 22695
rect 14924 22652 14976 22661
rect 15016 22695 15068 22704
rect 15016 22661 15025 22695
rect 15025 22661 15059 22695
rect 15059 22661 15068 22695
rect 15016 22652 15068 22661
rect 17408 22720 17460 22772
rect 17868 22720 17920 22772
rect 17960 22720 18012 22772
rect 37372 22720 37424 22772
rect 18328 22652 18380 22704
rect 6644 22516 6696 22568
rect 14648 22627 14700 22636
rect 14648 22593 14657 22627
rect 14657 22593 14691 22627
rect 14691 22593 14700 22627
rect 14648 22584 14700 22593
rect 17316 22627 17368 22636
rect 17316 22593 17325 22627
rect 17325 22593 17359 22627
rect 17359 22593 17368 22627
rect 17316 22584 17368 22593
rect 17592 22627 17644 22636
rect 17592 22593 17601 22627
rect 17601 22593 17635 22627
rect 17635 22593 17644 22627
rect 17592 22584 17644 22593
rect 7472 22448 7524 22500
rect 8392 22448 8444 22500
rect 11980 22448 12032 22500
rect 3608 22380 3660 22432
rect 14280 22448 14332 22500
rect 40500 22627 40552 22636
rect 40500 22593 40509 22627
rect 40509 22593 40543 22627
rect 40543 22593 40552 22627
rect 40500 22584 40552 22593
rect 32956 22516 33008 22568
rect 38844 22516 38896 22568
rect 14372 22423 14424 22432
rect 14372 22389 14381 22423
rect 14381 22389 14415 22423
rect 14415 22389 14424 22423
rect 14372 22380 14424 22389
rect 1950 22278 2002 22330
rect 2014 22278 2066 22330
rect 2078 22278 2130 22330
rect 2142 22278 2194 22330
rect 2206 22278 2258 22330
rect 6950 22278 7002 22330
rect 7014 22278 7066 22330
rect 7078 22278 7130 22330
rect 7142 22278 7194 22330
rect 7206 22278 7258 22330
rect 11950 22278 12002 22330
rect 12014 22278 12066 22330
rect 12078 22278 12130 22330
rect 12142 22278 12194 22330
rect 12206 22278 12258 22330
rect 16950 22278 17002 22330
rect 17014 22278 17066 22330
rect 17078 22278 17130 22330
rect 17142 22278 17194 22330
rect 17206 22278 17258 22330
rect 21950 22278 22002 22330
rect 22014 22278 22066 22330
rect 22078 22278 22130 22330
rect 22142 22278 22194 22330
rect 22206 22278 22258 22330
rect 26950 22278 27002 22330
rect 27014 22278 27066 22330
rect 27078 22278 27130 22330
rect 27142 22278 27194 22330
rect 27206 22278 27258 22330
rect 31950 22278 32002 22330
rect 32014 22278 32066 22330
rect 32078 22278 32130 22330
rect 32142 22278 32194 22330
rect 32206 22278 32258 22330
rect 36950 22278 37002 22330
rect 37014 22278 37066 22330
rect 37078 22278 37130 22330
rect 37142 22278 37194 22330
rect 37206 22278 37258 22330
rect 17316 22176 17368 22228
rect 17592 22176 17644 22228
rect 9036 22108 9088 22160
rect 11612 22108 11664 22160
rect 18604 22108 18656 22160
rect 15292 22083 15344 22092
rect 15292 22049 15301 22083
rect 15301 22049 15335 22083
rect 15335 22049 15344 22083
rect 15292 22040 15344 22049
rect 17224 22040 17276 22092
rect 17408 22040 17460 22092
rect 25044 22040 25096 22092
rect 26240 22040 26292 22092
rect 14832 22015 14884 22024
rect 14832 21981 14841 22015
rect 14841 21981 14875 22015
rect 14875 21981 14884 22015
rect 14832 21972 14884 21981
rect 26148 21972 26200 22024
rect 38844 22040 38896 22092
rect 17500 21836 17552 21888
rect 17868 21836 17920 21888
rect 2610 21734 2662 21786
rect 2674 21734 2726 21786
rect 2738 21734 2790 21786
rect 2802 21734 2854 21786
rect 2866 21734 2918 21786
rect 7610 21734 7662 21786
rect 7674 21734 7726 21786
rect 7738 21734 7790 21786
rect 7802 21734 7854 21786
rect 7866 21734 7918 21786
rect 12610 21734 12662 21786
rect 12674 21734 12726 21786
rect 12738 21734 12790 21786
rect 12802 21734 12854 21786
rect 12866 21734 12918 21786
rect 17610 21734 17662 21786
rect 17674 21734 17726 21786
rect 17738 21734 17790 21786
rect 17802 21734 17854 21786
rect 17866 21734 17918 21786
rect 22610 21734 22662 21786
rect 22674 21734 22726 21786
rect 22738 21734 22790 21786
rect 22802 21734 22854 21786
rect 22866 21734 22918 21786
rect 27610 21734 27662 21786
rect 27674 21734 27726 21786
rect 27738 21734 27790 21786
rect 27802 21734 27854 21786
rect 27866 21734 27918 21786
rect 32610 21734 32662 21786
rect 32674 21734 32726 21786
rect 32738 21734 32790 21786
rect 32802 21734 32854 21786
rect 32866 21734 32918 21786
rect 37610 21734 37662 21786
rect 37674 21734 37726 21786
rect 37738 21734 37790 21786
rect 37802 21734 37854 21786
rect 37866 21734 37918 21786
rect 31760 21428 31812 21480
rect 39028 21428 39080 21480
rect 11704 21360 11756 21412
rect 12440 21360 12492 21412
rect 17224 21360 17276 21412
rect 38476 21360 38528 21412
rect 7840 21292 7892 21344
rect 33232 21292 33284 21344
rect 1950 21190 2002 21242
rect 2014 21190 2066 21242
rect 2078 21190 2130 21242
rect 2142 21190 2194 21242
rect 2206 21190 2258 21242
rect 6950 21190 7002 21242
rect 7014 21190 7066 21242
rect 7078 21190 7130 21242
rect 7142 21190 7194 21242
rect 7206 21190 7258 21242
rect 11950 21190 12002 21242
rect 12014 21190 12066 21242
rect 12078 21190 12130 21242
rect 12142 21190 12194 21242
rect 12206 21190 12258 21242
rect 16950 21190 17002 21242
rect 17014 21190 17066 21242
rect 17078 21190 17130 21242
rect 17142 21190 17194 21242
rect 17206 21190 17258 21242
rect 21950 21190 22002 21242
rect 22014 21190 22066 21242
rect 22078 21190 22130 21242
rect 22142 21190 22194 21242
rect 22206 21190 22258 21242
rect 26950 21190 27002 21242
rect 27014 21190 27066 21242
rect 27078 21190 27130 21242
rect 27142 21190 27194 21242
rect 27206 21190 27258 21242
rect 31950 21190 32002 21242
rect 32014 21190 32066 21242
rect 32078 21190 32130 21242
rect 32142 21190 32194 21242
rect 32206 21190 32258 21242
rect 36950 21190 37002 21242
rect 37014 21190 37066 21242
rect 37078 21190 37130 21242
rect 37142 21190 37194 21242
rect 37206 21190 37258 21242
rect 12992 21088 13044 21140
rect 15936 21020 15988 21072
rect 3424 20927 3476 20936
rect 3424 20893 3433 20927
rect 3433 20893 3467 20927
rect 3467 20893 3476 20927
rect 3424 20884 3476 20893
rect 3516 20927 3568 20936
rect 3516 20893 3525 20927
rect 3525 20893 3559 20927
rect 3559 20893 3568 20927
rect 3516 20884 3568 20893
rect 10600 20952 10652 21004
rect 7840 20927 7892 20936
rect 7840 20893 7849 20927
rect 7849 20893 7883 20927
rect 7883 20893 7892 20927
rect 7840 20884 7892 20893
rect 4988 20816 5040 20868
rect 9312 20816 9364 20868
rect 22468 21020 22520 21072
rect 22284 20995 22336 21004
rect 22284 20961 22293 20995
rect 22293 20961 22327 20995
rect 22327 20961 22336 20995
rect 22284 20952 22336 20961
rect 24032 20952 24084 21004
rect 21824 20884 21876 20936
rect 22376 20927 22428 20936
rect 22376 20893 22385 20927
rect 22385 20893 22419 20927
rect 22419 20893 22428 20927
rect 22376 20884 22428 20893
rect 27344 20816 27396 20868
rect 4804 20748 4856 20800
rect 2610 20646 2662 20698
rect 2674 20646 2726 20698
rect 2738 20646 2790 20698
rect 2802 20646 2854 20698
rect 2866 20646 2918 20698
rect 7610 20646 7662 20698
rect 7674 20646 7726 20698
rect 7738 20646 7790 20698
rect 7802 20646 7854 20698
rect 7866 20646 7918 20698
rect 12610 20646 12662 20698
rect 12674 20646 12726 20698
rect 12738 20646 12790 20698
rect 12802 20646 12854 20698
rect 12866 20646 12918 20698
rect 17610 20646 17662 20698
rect 17674 20646 17726 20698
rect 17738 20646 17790 20698
rect 17802 20646 17854 20698
rect 17866 20646 17918 20698
rect 22610 20646 22662 20698
rect 22674 20646 22726 20698
rect 22738 20646 22790 20698
rect 22802 20646 22854 20698
rect 22866 20646 22918 20698
rect 27610 20646 27662 20698
rect 27674 20646 27726 20698
rect 27738 20646 27790 20698
rect 27802 20646 27854 20698
rect 27866 20646 27918 20698
rect 32610 20646 32662 20698
rect 32674 20646 32726 20698
rect 32738 20646 32790 20698
rect 32802 20646 32854 20698
rect 32866 20646 32918 20698
rect 37610 20646 37662 20698
rect 37674 20646 37726 20698
rect 37738 20646 37790 20698
rect 37802 20646 37854 20698
rect 37866 20646 37918 20698
rect 1676 20587 1728 20596
rect 1676 20553 1685 20587
rect 1685 20553 1719 20587
rect 1719 20553 1728 20587
rect 1676 20544 1728 20553
rect 20628 20544 20680 20596
rect 1584 20476 1636 20528
rect 23020 20476 23072 20528
rect 24952 20544 25004 20596
rect 37464 20544 37516 20596
rect 5080 20408 5132 20460
rect 24124 20451 24176 20460
rect 24124 20417 24133 20451
rect 24133 20417 24167 20451
rect 24167 20417 24176 20451
rect 24124 20408 24176 20417
rect 35716 20476 35768 20528
rect 22376 20340 22428 20392
rect 23296 20340 23348 20392
rect 24676 20383 24728 20392
rect 24676 20349 24685 20383
rect 24685 20349 24719 20383
rect 24719 20349 24728 20383
rect 24676 20340 24728 20349
rect 24584 20315 24636 20324
rect 24584 20281 24593 20315
rect 24593 20281 24627 20315
rect 24627 20281 24636 20315
rect 24584 20272 24636 20281
rect 23296 20204 23348 20256
rect 27344 20408 27396 20460
rect 34980 20408 35032 20460
rect 33140 20247 33192 20256
rect 33140 20213 33149 20247
rect 33149 20213 33183 20247
rect 33183 20213 33192 20247
rect 33140 20204 33192 20213
rect 35072 20340 35124 20392
rect 35164 20204 35216 20256
rect 1950 20102 2002 20154
rect 2014 20102 2066 20154
rect 2078 20102 2130 20154
rect 2142 20102 2194 20154
rect 2206 20102 2258 20154
rect 6950 20102 7002 20154
rect 7014 20102 7066 20154
rect 7078 20102 7130 20154
rect 7142 20102 7194 20154
rect 7206 20102 7258 20154
rect 11950 20102 12002 20154
rect 12014 20102 12066 20154
rect 12078 20102 12130 20154
rect 12142 20102 12194 20154
rect 12206 20102 12258 20154
rect 16950 20102 17002 20154
rect 17014 20102 17066 20154
rect 17078 20102 17130 20154
rect 17142 20102 17194 20154
rect 17206 20102 17258 20154
rect 21950 20102 22002 20154
rect 22014 20102 22066 20154
rect 22078 20102 22130 20154
rect 22142 20102 22194 20154
rect 22206 20102 22258 20154
rect 26950 20102 27002 20154
rect 27014 20102 27066 20154
rect 27078 20102 27130 20154
rect 27142 20102 27194 20154
rect 27206 20102 27258 20154
rect 31950 20102 32002 20154
rect 32014 20102 32066 20154
rect 32078 20102 32130 20154
rect 32142 20102 32194 20154
rect 32206 20102 32258 20154
rect 36950 20102 37002 20154
rect 37014 20102 37066 20154
rect 37078 20102 37130 20154
rect 37142 20102 37194 20154
rect 37206 20102 37258 20154
rect 18420 20000 18472 20052
rect 27344 20000 27396 20052
rect 33232 20000 33284 20052
rect 33508 20000 33560 20052
rect 4620 19932 4672 19984
rect 19524 19932 19576 19984
rect 4344 19839 4396 19848
rect 4344 19805 4353 19839
rect 4353 19805 4387 19839
rect 4387 19805 4396 19839
rect 4344 19796 4396 19805
rect 8024 19864 8076 19916
rect 13176 19864 13228 19916
rect 18236 19864 18288 19916
rect 37464 19907 37516 19916
rect 37464 19873 37473 19907
rect 37473 19873 37507 19907
rect 37507 19873 37516 19907
rect 37464 19864 37516 19873
rect 15752 19839 15804 19848
rect 15752 19805 15761 19839
rect 15761 19805 15795 19839
rect 15795 19805 15804 19839
rect 15752 19796 15804 19805
rect 33232 19839 33284 19848
rect 33232 19805 33241 19839
rect 33241 19805 33275 19839
rect 33275 19805 33284 19839
rect 33232 19796 33284 19805
rect 33324 19796 33376 19848
rect 37372 19796 37424 19848
rect 38016 19932 38068 19984
rect 17408 19728 17460 19780
rect 18512 19728 18564 19780
rect 18696 19728 18748 19780
rect 6276 19660 6328 19712
rect 7196 19660 7248 19712
rect 8116 19660 8168 19712
rect 30840 19660 30892 19712
rect 33232 19660 33284 19712
rect 33784 19660 33836 19712
rect 2610 19558 2662 19610
rect 2674 19558 2726 19610
rect 2738 19558 2790 19610
rect 2802 19558 2854 19610
rect 2866 19558 2918 19610
rect 7610 19558 7662 19610
rect 7674 19558 7726 19610
rect 7738 19558 7790 19610
rect 7802 19558 7854 19610
rect 7866 19558 7918 19610
rect 12610 19558 12662 19610
rect 12674 19558 12726 19610
rect 12738 19558 12790 19610
rect 12802 19558 12854 19610
rect 12866 19558 12918 19610
rect 17610 19558 17662 19610
rect 17674 19558 17726 19610
rect 17738 19558 17790 19610
rect 17802 19558 17854 19610
rect 17866 19558 17918 19610
rect 22610 19558 22662 19610
rect 22674 19558 22726 19610
rect 22738 19558 22790 19610
rect 22802 19558 22854 19610
rect 22866 19558 22918 19610
rect 27610 19558 27662 19610
rect 27674 19558 27726 19610
rect 27738 19558 27790 19610
rect 27802 19558 27854 19610
rect 27866 19558 27918 19610
rect 32610 19558 32662 19610
rect 32674 19558 32726 19610
rect 32738 19558 32790 19610
rect 32802 19558 32854 19610
rect 32866 19558 32918 19610
rect 37610 19558 37662 19610
rect 37674 19558 37726 19610
rect 37738 19558 37790 19610
rect 37802 19558 37854 19610
rect 37866 19558 37918 19610
rect 18972 19456 19024 19508
rect 24676 19456 24728 19508
rect 33140 19456 33192 19508
rect 7196 19320 7248 19372
rect 8024 19388 8076 19440
rect 9496 19320 9548 19372
rect 18420 19388 18472 19440
rect 18696 19320 18748 19372
rect 8024 19252 8076 19304
rect 8208 19252 8260 19304
rect 17868 19116 17920 19168
rect 22284 19116 22336 19168
rect 1950 19014 2002 19066
rect 2014 19014 2066 19066
rect 2078 19014 2130 19066
rect 2142 19014 2194 19066
rect 2206 19014 2258 19066
rect 6950 19014 7002 19066
rect 7014 19014 7066 19066
rect 7078 19014 7130 19066
rect 7142 19014 7194 19066
rect 7206 19014 7258 19066
rect 11950 19014 12002 19066
rect 12014 19014 12066 19066
rect 12078 19014 12130 19066
rect 12142 19014 12194 19066
rect 12206 19014 12258 19066
rect 16950 19014 17002 19066
rect 17014 19014 17066 19066
rect 17078 19014 17130 19066
rect 17142 19014 17194 19066
rect 17206 19014 17258 19066
rect 21950 19014 22002 19066
rect 22014 19014 22066 19066
rect 22078 19014 22130 19066
rect 22142 19014 22194 19066
rect 22206 19014 22258 19066
rect 26950 19014 27002 19066
rect 27014 19014 27066 19066
rect 27078 19014 27130 19066
rect 27142 19014 27194 19066
rect 27206 19014 27258 19066
rect 31950 19014 32002 19066
rect 32014 19014 32066 19066
rect 32078 19014 32130 19066
rect 32142 19014 32194 19066
rect 32206 19014 32258 19066
rect 36950 19014 37002 19066
rect 37014 19014 37066 19066
rect 37078 19014 37130 19066
rect 37142 19014 37194 19066
rect 37206 19014 37258 19066
rect 10968 18776 11020 18828
rect 25596 18844 25648 18896
rect 21088 18776 21140 18828
rect 17868 18751 17920 18760
rect 17868 18717 17877 18751
rect 17877 18717 17911 18751
rect 17911 18717 17920 18751
rect 17868 18708 17920 18717
rect 18420 18708 18472 18760
rect 18604 18708 18656 18760
rect 18696 18751 18748 18760
rect 18696 18717 18705 18751
rect 18705 18717 18739 18751
rect 18739 18717 18748 18751
rect 18696 18708 18748 18717
rect 26240 18751 26292 18760
rect 26240 18717 26249 18751
rect 26249 18717 26283 18751
rect 26283 18717 26292 18751
rect 26240 18708 26292 18717
rect 26424 18751 26476 18760
rect 26424 18717 26433 18751
rect 26433 18717 26467 18751
rect 26467 18717 26476 18751
rect 26424 18708 26476 18717
rect 26608 18708 26660 18760
rect 30932 18640 30984 18692
rect 19524 18572 19576 18624
rect 2610 18470 2662 18522
rect 2674 18470 2726 18522
rect 2738 18470 2790 18522
rect 2802 18470 2854 18522
rect 2866 18470 2918 18522
rect 7610 18470 7662 18522
rect 7674 18470 7726 18522
rect 7738 18470 7790 18522
rect 7802 18470 7854 18522
rect 7866 18470 7918 18522
rect 12610 18470 12662 18522
rect 12674 18470 12726 18522
rect 12738 18470 12790 18522
rect 12802 18470 12854 18522
rect 12866 18470 12918 18522
rect 17610 18470 17662 18522
rect 17674 18470 17726 18522
rect 17738 18470 17790 18522
rect 17802 18470 17854 18522
rect 17866 18470 17918 18522
rect 22610 18470 22662 18522
rect 22674 18470 22726 18522
rect 22738 18470 22790 18522
rect 22802 18470 22854 18522
rect 22866 18470 22918 18522
rect 27610 18470 27662 18522
rect 27674 18470 27726 18522
rect 27738 18470 27790 18522
rect 27802 18470 27854 18522
rect 27866 18470 27918 18522
rect 32610 18470 32662 18522
rect 32674 18470 32726 18522
rect 32738 18470 32790 18522
rect 32802 18470 32854 18522
rect 32866 18470 32918 18522
rect 37610 18470 37662 18522
rect 37674 18470 37726 18522
rect 37738 18470 37790 18522
rect 37802 18470 37854 18522
rect 37866 18470 37918 18522
rect 7472 18368 7524 18420
rect 8116 18368 8168 18420
rect 29644 18368 29696 18420
rect 35624 18368 35676 18420
rect 25412 18232 25464 18284
rect 29552 18232 29604 18284
rect 30104 18232 30156 18284
rect 25688 18164 25740 18216
rect 33876 18028 33928 18080
rect 37372 18028 37424 18080
rect 1950 17926 2002 17978
rect 2014 17926 2066 17978
rect 2078 17926 2130 17978
rect 2142 17926 2194 17978
rect 2206 17926 2258 17978
rect 6950 17926 7002 17978
rect 7014 17926 7066 17978
rect 7078 17926 7130 17978
rect 7142 17926 7194 17978
rect 7206 17926 7258 17978
rect 11950 17926 12002 17978
rect 12014 17926 12066 17978
rect 12078 17926 12130 17978
rect 12142 17926 12194 17978
rect 12206 17926 12258 17978
rect 16950 17926 17002 17978
rect 17014 17926 17066 17978
rect 17078 17926 17130 17978
rect 17142 17926 17194 17978
rect 17206 17926 17258 17978
rect 21950 17926 22002 17978
rect 22014 17926 22066 17978
rect 22078 17926 22130 17978
rect 22142 17926 22194 17978
rect 22206 17926 22258 17978
rect 26950 17926 27002 17978
rect 27014 17926 27066 17978
rect 27078 17926 27130 17978
rect 27142 17926 27194 17978
rect 27206 17926 27258 17978
rect 31950 17926 32002 17978
rect 32014 17926 32066 17978
rect 32078 17926 32130 17978
rect 32142 17926 32194 17978
rect 32206 17926 32258 17978
rect 36950 17926 37002 17978
rect 37014 17926 37066 17978
rect 37078 17926 37130 17978
rect 37142 17926 37194 17978
rect 37206 17926 37258 17978
rect 34336 17824 34388 17876
rect 35348 17824 35400 17876
rect 36728 17824 36780 17876
rect 24216 17688 24268 17740
rect 18880 17620 18932 17672
rect 38936 17663 38988 17672
rect 38936 17629 38945 17663
rect 38945 17629 38979 17663
rect 38979 17629 38988 17663
rect 38936 17620 38988 17629
rect 35072 17552 35124 17604
rect 4528 17484 4580 17536
rect 14556 17484 14608 17536
rect 2610 17382 2662 17434
rect 2674 17382 2726 17434
rect 2738 17382 2790 17434
rect 2802 17382 2854 17434
rect 2866 17382 2918 17434
rect 7610 17382 7662 17434
rect 7674 17382 7726 17434
rect 7738 17382 7790 17434
rect 7802 17382 7854 17434
rect 7866 17382 7918 17434
rect 12610 17382 12662 17434
rect 12674 17382 12726 17434
rect 12738 17382 12790 17434
rect 12802 17382 12854 17434
rect 12866 17382 12918 17434
rect 17610 17382 17662 17434
rect 17674 17382 17726 17434
rect 17738 17382 17790 17434
rect 17802 17382 17854 17434
rect 17866 17382 17918 17434
rect 22610 17382 22662 17434
rect 22674 17382 22726 17434
rect 22738 17382 22790 17434
rect 22802 17382 22854 17434
rect 22866 17382 22918 17434
rect 27610 17382 27662 17434
rect 27674 17382 27726 17434
rect 27738 17382 27790 17434
rect 27802 17382 27854 17434
rect 27866 17382 27918 17434
rect 32610 17382 32662 17434
rect 32674 17382 32726 17434
rect 32738 17382 32790 17434
rect 32802 17382 32854 17434
rect 32866 17382 32918 17434
rect 37610 17382 37662 17434
rect 37674 17382 37726 17434
rect 37738 17382 37790 17434
rect 37802 17382 37854 17434
rect 37866 17382 37918 17434
rect 3056 17280 3108 17332
rect 18144 17280 18196 17332
rect 7472 17212 7524 17264
rect 30012 17212 30064 17264
rect 1950 16838 2002 16890
rect 2014 16838 2066 16890
rect 2078 16838 2130 16890
rect 2142 16838 2194 16890
rect 2206 16838 2258 16890
rect 6950 16838 7002 16890
rect 7014 16838 7066 16890
rect 7078 16838 7130 16890
rect 7142 16838 7194 16890
rect 7206 16838 7258 16890
rect 11950 16838 12002 16890
rect 12014 16838 12066 16890
rect 12078 16838 12130 16890
rect 12142 16838 12194 16890
rect 12206 16838 12258 16890
rect 16950 16838 17002 16890
rect 17014 16838 17066 16890
rect 17078 16838 17130 16890
rect 17142 16838 17194 16890
rect 17206 16838 17258 16890
rect 21950 16838 22002 16890
rect 22014 16838 22066 16890
rect 22078 16838 22130 16890
rect 22142 16838 22194 16890
rect 22206 16838 22258 16890
rect 26950 16838 27002 16890
rect 27014 16838 27066 16890
rect 27078 16838 27130 16890
rect 27142 16838 27194 16890
rect 27206 16838 27258 16890
rect 31950 16838 32002 16890
rect 32014 16838 32066 16890
rect 32078 16838 32130 16890
rect 32142 16838 32194 16890
rect 32206 16838 32258 16890
rect 36950 16838 37002 16890
rect 37014 16838 37066 16890
rect 37078 16838 37130 16890
rect 37142 16838 37194 16890
rect 37206 16838 37258 16890
rect 22284 16736 22336 16788
rect 6552 16643 6604 16652
rect 6552 16609 6561 16643
rect 6561 16609 6595 16643
rect 6595 16609 6604 16643
rect 6552 16600 6604 16609
rect 22376 16668 22428 16720
rect 24492 16643 24544 16652
rect 24492 16609 24501 16643
rect 24501 16609 24535 16643
rect 24535 16609 24544 16643
rect 24492 16600 24544 16609
rect 34612 16600 34664 16652
rect 7380 16532 7432 16584
rect 24952 16575 25004 16584
rect 24952 16541 24961 16575
rect 24961 16541 24995 16575
rect 24995 16541 25004 16575
rect 24952 16532 25004 16541
rect 25596 16532 25648 16584
rect 28448 16464 28500 16516
rect 35256 16464 35308 16516
rect 2610 16294 2662 16346
rect 2674 16294 2726 16346
rect 2738 16294 2790 16346
rect 2802 16294 2854 16346
rect 2866 16294 2918 16346
rect 7610 16294 7662 16346
rect 7674 16294 7726 16346
rect 7738 16294 7790 16346
rect 7802 16294 7854 16346
rect 7866 16294 7918 16346
rect 12610 16294 12662 16346
rect 12674 16294 12726 16346
rect 12738 16294 12790 16346
rect 12802 16294 12854 16346
rect 12866 16294 12918 16346
rect 17610 16294 17662 16346
rect 17674 16294 17726 16346
rect 17738 16294 17790 16346
rect 17802 16294 17854 16346
rect 17866 16294 17918 16346
rect 22610 16294 22662 16346
rect 22674 16294 22726 16346
rect 22738 16294 22790 16346
rect 22802 16294 22854 16346
rect 22866 16294 22918 16346
rect 27610 16294 27662 16346
rect 27674 16294 27726 16346
rect 27738 16294 27790 16346
rect 27802 16294 27854 16346
rect 27866 16294 27918 16346
rect 32610 16294 32662 16346
rect 32674 16294 32726 16346
rect 32738 16294 32790 16346
rect 32802 16294 32854 16346
rect 32866 16294 32918 16346
rect 37610 16294 37662 16346
rect 37674 16294 37726 16346
rect 37738 16294 37790 16346
rect 37802 16294 37854 16346
rect 37866 16294 37918 16346
rect 3516 16192 3568 16244
rect 2320 16056 2372 16108
rect 6368 16056 6420 16108
rect 9220 16056 9272 16108
rect 9404 15988 9456 16040
rect 24860 15988 24912 16040
rect 6184 15920 6236 15972
rect 31024 15920 31076 15972
rect 2320 15852 2372 15904
rect 11796 15852 11848 15904
rect 39304 15852 39356 15904
rect 1950 15750 2002 15802
rect 2014 15750 2066 15802
rect 2078 15750 2130 15802
rect 2142 15750 2194 15802
rect 2206 15750 2258 15802
rect 6950 15750 7002 15802
rect 7014 15750 7066 15802
rect 7078 15750 7130 15802
rect 7142 15750 7194 15802
rect 7206 15750 7258 15802
rect 11950 15750 12002 15802
rect 12014 15750 12066 15802
rect 12078 15750 12130 15802
rect 12142 15750 12194 15802
rect 12206 15750 12258 15802
rect 16950 15750 17002 15802
rect 17014 15750 17066 15802
rect 17078 15750 17130 15802
rect 17142 15750 17194 15802
rect 17206 15750 17258 15802
rect 21950 15750 22002 15802
rect 22014 15750 22066 15802
rect 22078 15750 22130 15802
rect 22142 15750 22194 15802
rect 22206 15750 22258 15802
rect 26950 15750 27002 15802
rect 27014 15750 27066 15802
rect 27078 15750 27130 15802
rect 27142 15750 27194 15802
rect 27206 15750 27258 15802
rect 31950 15750 32002 15802
rect 32014 15750 32066 15802
rect 32078 15750 32130 15802
rect 32142 15750 32194 15802
rect 32206 15750 32258 15802
rect 36950 15750 37002 15802
rect 37014 15750 37066 15802
rect 37078 15750 37130 15802
rect 37142 15750 37194 15802
rect 37206 15750 37258 15802
rect 12992 15691 13044 15700
rect 12992 15657 13001 15691
rect 13001 15657 13035 15691
rect 13035 15657 13044 15691
rect 12992 15648 13044 15657
rect 13452 15691 13504 15700
rect 13452 15657 13461 15691
rect 13461 15657 13495 15691
rect 13495 15657 13504 15691
rect 13452 15648 13504 15657
rect 13176 15487 13228 15496
rect 13176 15453 13185 15487
rect 13185 15453 13219 15487
rect 13219 15453 13228 15487
rect 13176 15444 13228 15453
rect 34704 15487 34756 15496
rect 34704 15453 34713 15487
rect 34713 15453 34747 15487
rect 34747 15453 34756 15487
rect 34704 15444 34756 15453
rect 38200 15444 38252 15496
rect 38568 15444 38620 15496
rect 13084 15376 13136 15428
rect 13268 15419 13320 15428
rect 13268 15385 13277 15419
rect 13277 15385 13311 15419
rect 13311 15385 13320 15419
rect 13268 15376 13320 15385
rect 35532 15419 35584 15428
rect 35532 15385 35541 15419
rect 35541 15385 35575 15419
rect 35575 15385 35584 15419
rect 35532 15376 35584 15385
rect 38384 15308 38436 15360
rect 38568 15308 38620 15360
rect 2610 15206 2662 15258
rect 2674 15206 2726 15258
rect 2738 15206 2790 15258
rect 2802 15206 2854 15258
rect 2866 15206 2918 15258
rect 7610 15206 7662 15258
rect 7674 15206 7726 15258
rect 7738 15206 7790 15258
rect 7802 15206 7854 15258
rect 7866 15206 7918 15258
rect 12610 15206 12662 15258
rect 12674 15206 12726 15258
rect 12738 15206 12790 15258
rect 12802 15206 12854 15258
rect 12866 15206 12918 15258
rect 17610 15206 17662 15258
rect 17674 15206 17726 15258
rect 17738 15206 17790 15258
rect 17802 15206 17854 15258
rect 17866 15206 17918 15258
rect 22610 15206 22662 15258
rect 22674 15206 22726 15258
rect 22738 15206 22790 15258
rect 22802 15206 22854 15258
rect 22866 15206 22918 15258
rect 27610 15206 27662 15258
rect 27674 15206 27726 15258
rect 27738 15206 27790 15258
rect 27802 15206 27854 15258
rect 27866 15206 27918 15258
rect 32610 15206 32662 15258
rect 32674 15206 32726 15258
rect 32738 15206 32790 15258
rect 32802 15206 32854 15258
rect 32866 15206 32918 15258
rect 37610 15206 37662 15258
rect 37674 15206 37726 15258
rect 37738 15206 37790 15258
rect 37802 15206 37854 15258
rect 37866 15206 37918 15258
rect 14556 15079 14608 15088
rect 14556 15045 14565 15079
rect 14565 15045 14599 15079
rect 14599 15045 14608 15079
rect 14556 15036 14608 15045
rect 17224 15104 17276 15156
rect 18420 15104 18472 15156
rect 20076 15104 20128 15156
rect 21824 15104 21876 15156
rect 16580 15036 16632 15088
rect 23572 14968 23624 15020
rect 17224 14900 17276 14952
rect 31024 15079 31076 15088
rect 31024 15045 31033 15079
rect 31033 15045 31067 15079
rect 31067 15045 31076 15079
rect 31024 15036 31076 15045
rect 31208 15036 31260 15088
rect 31392 15011 31444 15020
rect 31392 14977 31401 15011
rect 31401 14977 31435 15011
rect 31435 14977 31444 15011
rect 31392 14968 31444 14977
rect 33692 15011 33744 15020
rect 33692 14977 33701 15011
rect 33701 14977 33735 15011
rect 33735 14977 33744 15011
rect 33692 14968 33744 14977
rect 34244 15011 34296 15020
rect 34244 14977 34253 15011
rect 34253 14977 34287 15011
rect 34287 14977 34296 15011
rect 34244 14968 34296 14977
rect 37372 15036 37424 15088
rect 38660 15036 38712 15088
rect 31484 14832 31536 14884
rect 26608 14764 26660 14816
rect 34336 14943 34388 14952
rect 34336 14909 34345 14943
rect 34345 14909 34379 14943
rect 34379 14909 34388 14943
rect 34336 14900 34388 14909
rect 31760 14875 31812 14884
rect 31760 14841 31769 14875
rect 31769 14841 31803 14875
rect 31803 14841 31812 14875
rect 31760 14832 31812 14841
rect 35348 15011 35400 15020
rect 35348 14977 35357 15011
rect 35357 14977 35391 15011
rect 35391 14977 35400 15011
rect 35348 14968 35400 14977
rect 38292 15011 38344 15020
rect 38292 14977 38301 15011
rect 38301 14977 38335 15011
rect 38335 14977 38344 15011
rect 38292 14968 38344 14977
rect 34980 14943 35032 14952
rect 34980 14909 34989 14943
rect 34989 14909 35023 14943
rect 35023 14909 35032 14943
rect 34980 14900 35032 14909
rect 35256 14943 35308 14952
rect 35256 14909 35265 14943
rect 35265 14909 35299 14943
rect 35299 14909 35308 14943
rect 35256 14900 35308 14909
rect 39028 14832 39080 14884
rect 38200 14764 38252 14816
rect 1950 14662 2002 14714
rect 2014 14662 2066 14714
rect 2078 14662 2130 14714
rect 2142 14662 2194 14714
rect 2206 14662 2258 14714
rect 6950 14662 7002 14714
rect 7014 14662 7066 14714
rect 7078 14662 7130 14714
rect 7142 14662 7194 14714
rect 7206 14662 7258 14714
rect 11950 14662 12002 14714
rect 12014 14662 12066 14714
rect 12078 14662 12130 14714
rect 12142 14662 12194 14714
rect 12206 14662 12258 14714
rect 16950 14662 17002 14714
rect 17014 14662 17066 14714
rect 17078 14662 17130 14714
rect 17142 14662 17194 14714
rect 17206 14662 17258 14714
rect 21950 14662 22002 14714
rect 22014 14662 22066 14714
rect 22078 14662 22130 14714
rect 22142 14662 22194 14714
rect 22206 14662 22258 14714
rect 26950 14662 27002 14714
rect 27014 14662 27066 14714
rect 27078 14662 27130 14714
rect 27142 14662 27194 14714
rect 27206 14662 27258 14714
rect 31950 14662 32002 14714
rect 32014 14662 32066 14714
rect 32078 14662 32130 14714
rect 32142 14662 32194 14714
rect 32206 14662 32258 14714
rect 36950 14662 37002 14714
rect 37014 14662 37066 14714
rect 37078 14662 37130 14714
rect 37142 14662 37194 14714
rect 37206 14662 37258 14714
rect 9128 14560 9180 14612
rect 23480 14492 23532 14544
rect 29092 14492 29144 14544
rect 30104 14492 30156 14544
rect 32312 14492 32364 14544
rect 26516 14424 26568 14476
rect 30748 14356 30800 14408
rect 31300 14399 31352 14408
rect 31300 14365 31309 14399
rect 31309 14365 31343 14399
rect 31343 14365 31352 14399
rect 31300 14356 31352 14365
rect 32404 14424 32456 14476
rect 29828 14288 29880 14340
rect 31208 14288 31260 14340
rect 33416 14356 33468 14408
rect 39304 14399 39356 14408
rect 39304 14365 39313 14399
rect 39313 14365 39347 14399
rect 39347 14365 39356 14399
rect 39304 14356 39356 14365
rect 39488 14467 39540 14476
rect 39488 14433 39497 14467
rect 39497 14433 39531 14467
rect 39531 14433 39540 14467
rect 39488 14424 39540 14433
rect 35716 14220 35768 14272
rect 2610 14118 2662 14170
rect 2674 14118 2726 14170
rect 2738 14118 2790 14170
rect 2802 14118 2854 14170
rect 2866 14118 2918 14170
rect 7610 14118 7662 14170
rect 7674 14118 7726 14170
rect 7738 14118 7790 14170
rect 7802 14118 7854 14170
rect 7866 14118 7918 14170
rect 12610 14118 12662 14170
rect 12674 14118 12726 14170
rect 12738 14118 12790 14170
rect 12802 14118 12854 14170
rect 12866 14118 12918 14170
rect 17610 14118 17662 14170
rect 17674 14118 17726 14170
rect 17738 14118 17790 14170
rect 17802 14118 17854 14170
rect 17866 14118 17918 14170
rect 22610 14118 22662 14170
rect 22674 14118 22726 14170
rect 22738 14118 22790 14170
rect 22802 14118 22854 14170
rect 22866 14118 22918 14170
rect 27610 14118 27662 14170
rect 27674 14118 27726 14170
rect 27738 14118 27790 14170
rect 27802 14118 27854 14170
rect 27866 14118 27918 14170
rect 32610 14118 32662 14170
rect 32674 14118 32726 14170
rect 32738 14118 32790 14170
rect 32802 14118 32854 14170
rect 32866 14118 32918 14170
rect 37610 14118 37662 14170
rect 37674 14118 37726 14170
rect 37738 14118 37790 14170
rect 37802 14118 37854 14170
rect 37866 14118 37918 14170
rect 38752 14016 38804 14068
rect 1400 13923 1452 13932
rect 1400 13889 1409 13923
rect 1409 13889 1443 13923
rect 1443 13889 1452 13923
rect 1400 13880 1452 13889
rect 19156 13880 19208 13932
rect 38384 13923 38436 13932
rect 38384 13889 38393 13923
rect 38393 13889 38427 13923
rect 38427 13889 38436 13923
rect 38384 13880 38436 13889
rect 38844 13880 38896 13932
rect 39948 13880 40000 13932
rect 13544 13812 13596 13864
rect 33416 13812 33468 13864
rect 1950 13574 2002 13626
rect 2014 13574 2066 13626
rect 2078 13574 2130 13626
rect 2142 13574 2194 13626
rect 2206 13574 2258 13626
rect 6950 13574 7002 13626
rect 7014 13574 7066 13626
rect 7078 13574 7130 13626
rect 7142 13574 7194 13626
rect 7206 13574 7258 13626
rect 11950 13574 12002 13626
rect 12014 13574 12066 13626
rect 12078 13574 12130 13626
rect 12142 13574 12194 13626
rect 12206 13574 12258 13626
rect 16950 13574 17002 13626
rect 17014 13574 17066 13626
rect 17078 13574 17130 13626
rect 17142 13574 17194 13626
rect 17206 13574 17258 13626
rect 21950 13574 22002 13626
rect 22014 13574 22066 13626
rect 22078 13574 22130 13626
rect 22142 13574 22194 13626
rect 22206 13574 22258 13626
rect 26950 13574 27002 13626
rect 27014 13574 27066 13626
rect 27078 13574 27130 13626
rect 27142 13574 27194 13626
rect 27206 13574 27258 13626
rect 31950 13574 32002 13626
rect 32014 13574 32066 13626
rect 32078 13574 32130 13626
rect 32142 13574 32194 13626
rect 32206 13574 32258 13626
rect 36950 13574 37002 13626
rect 37014 13574 37066 13626
rect 37078 13574 37130 13626
rect 37142 13574 37194 13626
rect 37206 13574 37258 13626
rect 38752 13472 38804 13524
rect 34244 13336 34296 13388
rect 39028 13311 39080 13320
rect 39028 13277 39037 13311
rect 39037 13277 39071 13311
rect 39071 13277 39080 13311
rect 39028 13268 39080 13277
rect 35532 13200 35584 13252
rect 7380 13132 7432 13184
rect 21640 13132 21692 13184
rect 38568 13132 38620 13184
rect 2610 13030 2662 13082
rect 2674 13030 2726 13082
rect 2738 13030 2790 13082
rect 2802 13030 2854 13082
rect 2866 13030 2918 13082
rect 7610 13030 7662 13082
rect 7674 13030 7726 13082
rect 7738 13030 7790 13082
rect 7802 13030 7854 13082
rect 7866 13030 7918 13082
rect 12610 13030 12662 13082
rect 12674 13030 12726 13082
rect 12738 13030 12790 13082
rect 12802 13030 12854 13082
rect 12866 13030 12918 13082
rect 17610 13030 17662 13082
rect 17674 13030 17726 13082
rect 17738 13030 17790 13082
rect 17802 13030 17854 13082
rect 17866 13030 17918 13082
rect 22610 13030 22662 13082
rect 22674 13030 22726 13082
rect 22738 13030 22790 13082
rect 22802 13030 22854 13082
rect 22866 13030 22918 13082
rect 27610 13030 27662 13082
rect 27674 13030 27726 13082
rect 27738 13030 27790 13082
rect 27802 13030 27854 13082
rect 27866 13030 27918 13082
rect 32610 13030 32662 13082
rect 32674 13030 32726 13082
rect 32738 13030 32790 13082
rect 32802 13030 32854 13082
rect 32866 13030 32918 13082
rect 37610 13030 37662 13082
rect 37674 13030 37726 13082
rect 37738 13030 37790 13082
rect 37802 13030 37854 13082
rect 37866 13030 37918 13082
rect 23296 12971 23348 12980
rect 23296 12937 23305 12971
rect 23305 12937 23339 12971
rect 23339 12937 23348 12971
rect 23296 12928 23348 12937
rect 38752 12928 38804 12980
rect 21456 12792 21508 12844
rect 23388 12835 23440 12844
rect 23388 12801 23397 12835
rect 23397 12801 23431 12835
rect 23431 12801 23440 12835
rect 23388 12792 23440 12801
rect 30288 12724 30340 12776
rect 1950 12486 2002 12538
rect 2014 12486 2066 12538
rect 2078 12486 2130 12538
rect 2142 12486 2194 12538
rect 2206 12486 2258 12538
rect 6950 12486 7002 12538
rect 7014 12486 7066 12538
rect 7078 12486 7130 12538
rect 7142 12486 7194 12538
rect 7206 12486 7258 12538
rect 11950 12486 12002 12538
rect 12014 12486 12066 12538
rect 12078 12486 12130 12538
rect 12142 12486 12194 12538
rect 12206 12486 12258 12538
rect 16950 12486 17002 12538
rect 17014 12486 17066 12538
rect 17078 12486 17130 12538
rect 17142 12486 17194 12538
rect 17206 12486 17258 12538
rect 21950 12486 22002 12538
rect 22014 12486 22066 12538
rect 22078 12486 22130 12538
rect 22142 12486 22194 12538
rect 22206 12486 22258 12538
rect 26950 12486 27002 12538
rect 27014 12486 27066 12538
rect 27078 12486 27130 12538
rect 27142 12486 27194 12538
rect 27206 12486 27258 12538
rect 31950 12486 32002 12538
rect 32014 12486 32066 12538
rect 32078 12486 32130 12538
rect 32142 12486 32194 12538
rect 32206 12486 32258 12538
rect 36950 12486 37002 12538
rect 37014 12486 37066 12538
rect 37078 12486 37130 12538
rect 37142 12486 37194 12538
rect 37206 12486 37258 12538
rect 16488 12223 16540 12232
rect 16488 12189 16497 12223
rect 16497 12189 16531 12223
rect 16531 12189 16540 12223
rect 16488 12180 16540 12189
rect 21548 12248 21600 12300
rect 21364 12180 21416 12232
rect 31760 12112 31812 12164
rect 2610 11942 2662 11994
rect 2674 11942 2726 11994
rect 2738 11942 2790 11994
rect 2802 11942 2854 11994
rect 2866 11942 2918 11994
rect 7610 11942 7662 11994
rect 7674 11942 7726 11994
rect 7738 11942 7790 11994
rect 7802 11942 7854 11994
rect 7866 11942 7918 11994
rect 12610 11942 12662 11994
rect 12674 11942 12726 11994
rect 12738 11942 12790 11994
rect 12802 11942 12854 11994
rect 12866 11942 12918 11994
rect 17610 11942 17662 11994
rect 17674 11942 17726 11994
rect 17738 11942 17790 11994
rect 17802 11942 17854 11994
rect 17866 11942 17918 11994
rect 22610 11942 22662 11994
rect 22674 11942 22726 11994
rect 22738 11942 22790 11994
rect 22802 11942 22854 11994
rect 22866 11942 22918 11994
rect 27610 11942 27662 11994
rect 27674 11942 27726 11994
rect 27738 11942 27790 11994
rect 27802 11942 27854 11994
rect 27866 11942 27918 11994
rect 32610 11942 32662 11994
rect 32674 11942 32726 11994
rect 32738 11942 32790 11994
rect 32802 11942 32854 11994
rect 32866 11942 32918 11994
rect 37610 11942 37662 11994
rect 37674 11942 37726 11994
rect 37738 11942 37790 11994
rect 37802 11942 37854 11994
rect 37866 11942 37918 11994
rect 3148 11704 3200 11756
rect 29644 11704 29696 11756
rect 1950 11398 2002 11450
rect 2014 11398 2066 11450
rect 2078 11398 2130 11450
rect 2142 11398 2194 11450
rect 2206 11398 2258 11450
rect 6950 11398 7002 11450
rect 7014 11398 7066 11450
rect 7078 11398 7130 11450
rect 7142 11398 7194 11450
rect 7206 11398 7258 11450
rect 11950 11398 12002 11450
rect 12014 11398 12066 11450
rect 12078 11398 12130 11450
rect 12142 11398 12194 11450
rect 12206 11398 12258 11450
rect 16950 11398 17002 11450
rect 17014 11398 17066 11450
rect 17078 11398 17130 11450
rect 17142 11398 17194 11450
rect 17206 11398 17258 11450
rect 21950 11398 22002 11450
rect 22014 11398 22066 11450
rect 22078 11398 22130 11450
rect 22142 11398 22194 11450
rect 22206 11398 22258 11450
rect 26950 11398 27002 11450
rect 27014 11398 27066 11450
rect 27078 11398 27130 11450
rect 27142 11398 27194 11450
rect 27206 11398 27258 11450
rect 31950 11398 32002 11450
rect 32014 11398 32066 11450
rect 32078 11398 32130 11450
rect 32142 11398 32194 11450
rect 32206 11398 32258 11450
rect 36950 11398 37002 11450
rect 37014 11398 37066 11450
rect 37078 11398 37130 11450
rect 37142 11398 37194 11450
rect 37206 11398 37258 11450
rect 13268 11228 13320 11280
rect 2412 11135 2464 11144
rect 2412 11101 2421 11135
rect 2421 11101 2455 11135
rect 2455 11101 2464 11135
rect 2412 11092 2464 11101
rect 21088 11160 21140 11212
rect 23572 11160 23624 11212
rect 15108 11135 15160 11144
rect 15108 11101 15117 11135
rect 15117 11101 15151 11135
rect 15151 11101 15160 11135
rect 15108 11092 15160 11101
rect 16580 11092 16632 11144
rect 6092 11024 6144 11076
rect 18420 11024 18472 11076
rect 32404 11135 32456 11144
rect 32404 11101 32413 11135
rect 32413 11101 32447 11135
rect 32447 11101 32456 11135
rect 32404 11092 32456 11101
rect 33600 11135 33652 11144
rect 33600 11101 33609 11135
rect 33609 11101 33643 11135
rect 33643 11101 33652 11135
rect 33600 11092 33652 11101
rect 34612 11092 34664 11144
rect 21180 10956 21232 11008
rect 28172 10956 28224 11008
rect 2610 10854 2662 10906
rect 2674 10854 2726 10906
rect 2738 10854 2790 10906
rect 2802 10854 2854 10906
rect 2866 10854 2918 10906
rect 7610 10854 7662 10906
rect 7674 10854 7726 10906
rect 7738 10854 7790 10906
rect 7802 10854 7854 10906
rect 7866 10854 7918 10906
rect 12610 10854 12662 10906
rect 12674 10854 12726 10906
rect 12738 10854 12790 10906
rect 12802 10854 12854 10906
rect 12866 10854 12918 10906
rect 17610 10854 17662 10906
rect 17674 10854 17726 10906
rect 17738 10854 17790 10906
rect 17802 10854 17854 10906
rect 17866 10854 17918 10906
rect 22610 10854 22662 10906
rect 22674 10854 22726 10906
rect 22738 10854 22790 10906
rect 22802 10854 22854 10906
rect 22866 10854 22918 10906
rect 27610 10854 27662 10906
rect 27674 10854 27726 10906
rect 27738 10854 27790 10906
rect 27802 10854 27854 10906
rect 27866 10854 27918 10906
rect 32610 10854 32662 10906
rect 32674 10854 32726 10906
rect 32738 10854 32790 10906
rect 32802 10854 32854 10906
rect 32866 10854 32918 10906
rect 37610 10854 37662 10906
rect 37674 10854 37726 10906
rect 37738 10854 37790 10906
rect 37802 10854 37854 10906
rect 37866 10854 37918 10906
rect 3056 10659 3108 10668
rect 3056 10625 3065 10659
rect 3065 10625 3099 10659
rect 3099 10625 3108 10659
rect 3056 10616 3108 10625
rect 10968 10684 11020 10736
rect 20444 10684 20496 10736
rect 18696 10616 18748 10668
rect 12348 10548 12400 10600
rect 8208 10480 8260 10532
rect 17960 10480 18012 10532
rect 36820 10480 36872 10532
rect 9312 10412 9364 10464
rect 31208 10412 31260 10464
rect 1950 10310 2002 10362
rect 2014 10310 2066 10362
rect 2078 10310 2130 10362
rect 2142 10310 2194 10362
rect 2206 10310 2258 10362
rect 6950 10310 7002 10362
rect 7014 10310 7066 10362
rect 7078 10310 7130 10362
rect 7142 10310 7194 10362
rect 7206 10310 7258 10362
rect 11950 10310 12002 10362
rect 12014 10310 12066 10362
rect 12078 10310 12130 10362
rect 12142 10310 12194 10362
rect 12206 10310 12258 10362
rect 16950 10310 17002 10362
rect 17014 10310 17066 10362
rect 17078 10310 17130 10362
rect 17142 10310 17194 10362
rect 17206 10310 17258 10362
rect 21950 10310 22002 10362
rect 22014 10310 22066 10362
rect 22078 10310 22130 10362
rect 22142 10310 22194 10362
rect 22206 10310 22258 10362
rect 26950 10310 27002 10362
rect 27014 10310 27066 10362
rect 27078 10310 27130 10362
rect 27142 10310 27194 10362
rect 27206 10310 27258 10362
rect 31950 10310 32002 10362
rect 32014 10310 32066 10362
rect 32078 10310 32130 10362
rect 32142 10310 32194 10362
rect 32206 10310 32258 10362
rect 36950 10310 37002 10362
rect 37014 10310 37066 10362
rect 37078 10310 37130 10362
rect 37142 10310 37194 10362
rect 37206 10310 37258 10362
rect 2610 9766 2662 9818
rect 2674 9766 2726 9818
rect 2738 9766 2790 9818
rect 2802 9766 2854 9818
rect 2866 9766 2918 9818
rect 7610 9766 7662 9818
rect 7674 9766 7726 9818
rect 7738 9766 7790 9818
rect 7802 9766 7854 9818
rect 7866 9766 7918 9818
rect 12610 9766 12662 9818
rect 12674 9766 12726 9818
rect 12738 9766 12790 9818
rect 12802 9766 12854 9818
rect 12866 9766 12918 9818
rect 17610 9766 17662 9818
rect 17674 9766 17726 9818
rect 17738 9766 17790 9818
rect 17802 9766 17854 9818
rect 17866 9766 17918 9818
rect 22610 9766 22662 9818
rect 22674 9766 22726 9818
rect 22738 9766 22790 9818
rect 22802 9766 22854 9818
rect 22866 9766 22918 9818
rect 27610 9766 27662 9818
rect 27674 9766 27726 9818
rect 27738 9766 27790 9818
rect 27802 9766 27854 9818
rect 27866 9766 27918 9818
rect 32610 9766 32662 9818
rect 32674 9766 32726 9818
rect 32738 9766 32790 9818
rect 32802 9766 32854 9818
rect 32866 9766 32918 9818
rect 37610 9766 37662 9818
rect 37674 9766 37726 9818
rect 37738 9766 37790 9818
rect 37802 9766 37854 9818
rect 37866 9766 37918 9818
rect 12992 9596 13044 9648
rect 14188 9639 14240 9648
rect 14188 9605 14197 9639
rect 14197 9605 14231 9639
rect 14231 9605 14240 9639
rect 14188 9596 14240 9605
rect 13636 9571 13688 9580
rect 13636 9537 13645 9571
rect 13645 9537 13679 9571
rect 13679 9537 13688 9571
rect 13636 9528 13688 9537
rect 13820 9571 13872 9580
rect 13820 9537 13829 9571
rect 13829 9537 13863 9571
rect 13863 9537 13872 9571
rect 13820 9528 13872 9537
rect 2504 9460 2556 9512
rect 15660 9460 15712 9512
rect 16028 9460 16080 9512
rect 16580 9528 16632 9580
rect 16856 9639 16908 9648
rect 16856 9605 16865 9639
rect 16865 9605 16899 9639
rect 16899 9605 16908 9639
rect 16856 9596 16908 9605
rect 32404 9596 32456 9648
rect 17960 9528 18012 9580
rect 23480 9460 23532 9512
rect 17408 9392 17460 9444
rect 16672 9324 16724 9376
rect 1950 9222 2002 9274
rect 2014 9222 2066 9274
rect 2078 9222 2130 9274
rect 2142 9222 2194 9274
rect 2206 9222 2258 9274
rect 6950 9222 7002 9274
rect 7014 9222 7066 9274
rect 7078 9222 7130 9274
rect 7142 9222 7194 9274
rect 7206 9222 7258 9274
rect 11950 9222 12002 9274
rect 12014 9222 12066 9274
rect 12078 9222 12130 9274
rect 12142 9222 12194 9274
rect 12206 9222 12258 9274
rect 16950 9222 17002 9274
rect 17014 9222 17066 9274
rect 17078 9222 17130 9274
rect 17142 9222 17194 9274
rect 17206 9222 17258 9274
rect 21950 9222 22002 9274
rect 22014 9222 22066 9274
rect 22078 9222 22130 9274
rect 22142 9222 22194 9274
rect 22206 9222 22258 9274
rect 26950 9222 27002 9274
rect 27014 9222 27066 9274
rect 27078 9222 27130 9274
rect 27142 9222 27194 9274
rect 27206 9222 27258 9274
rect 31950 9222 32002 9274
rect 32014 9222 32066 9274
rect 32078 9222 32130 9274
rect 32142 9222 32194 9274
rect 32206 9222 32258 9274
rect 36950 9222 37002 9274
rect 37014 9222 37066 9274
rect 37078 9222 37130 9274
rect 37142 9222 37194 9274
rect 37206 9222 37258 9274
rect 35164 9163 35216 9172
rect 35164 9129 35173 9163
rect 35173 9129 35207 9163
rect 35207 9129 35216 9163
rect 35164 9120 35216 9129
rect 1860 9027 1912 9036
rect 1860 8993 1869 9027
rect 1869 8993 1903 9027
rect 1903 8993 1912 9027
rect 1860 8984 1912 8993
rect 3608 9052 3660 9104
rect 8208 9052 8260 9104
rect 19156 9052 19208 9104
rect 23388 9052 23440 9104
rect 2504 8916 2556 8968
rect 4896 8984 4948 9036
rect 30288 8984 30340 9036
rect 26700 8916 26752 8968
rect 27344 8916 27396 8968
rect 27528 8959 27580 8968
rect 27528 8925 27537 8959
rect 27537 8925 27571 8959
rect 27571 8925 27580 8959
rect 27528 8916 27580 8925
rect 35072 8916 35124 8968
rect 16580 8848 16632 8900
rect 20260 8848 20312 8900
rect 26424 8848 26476 8900
rect 2610 8678 2662 8730
rect 2674 8678 2726 8730
rect 2738 8678 2790 8730
rect 2802 8678 2854 8730
rect 2866 8678 2918 8730
rect 7610 8678 7662 8730
rect 7674 8678 7726 8730
rect 7738 8678 7790 8730
rect 7802 8678 7854 8730
rect 7866 8678 7918 8730
rect 12610 8678 12662 8730
rect 12674 8678 12726 8730
rect 12738 8678 12790 8730
rect 12802 8678 12854 8730
rect 12866 8678 12918 8730
rect 17610 8678 17662 8730
rect 17674 8678 17726 8730
rect 17738 8678 17790 8730
rect 17802 8678 17854 8730
rect 17866 8678 17918 8730
rect 22610 8678 22662 8730
rect 22674 8678 22726 8730
rect 22738 8678 22790 8730
rect 22802 8678 22854 8730
rect 22866 8678 22918 8730
rect 27610 8678 27662 8730
rect 27674 8678 27726 8730
rect 27738 8678 27790 8730
rect 27802 8678 27854 8730
rect 27866 8678 27918 8730
rect 32610 8678 32662 8730
rect 32674 8678 32726 8730
rect 32738 8678 32790 8730
rect 32802 8678 32854 8730
rect 32866 8678 32918 8730
rect 37610 8678 37662 8730
rect 37674 8678 37726 8730
rect 37738 8678 37790 8730
rect 37802 8678 37854 8730
rect 37866 8678 37918 8730
rect 16212 8304 16264 8356
rect 16672 8304 16724 8356
rect 34612 8304 34664 8356
rect 36268 8304 36320 8356
rect 1950 8134 2002 8186
rect 2014 8134 2066 8186
rect 2078 8134 2130 8186
rect 2142 8134 2194 8186
rect 2206 8134 2258 8186
rect 6950 8134 7002 8186
rect 7014 8134 7066 8186
rect 7078 8134 7130 8186
rect 7142 8134 7194 8186
rect 7206 8134 7258 8186
rect 11950 8134 12002 8186
rect 12014 8134 12066 8186
rect 12078 8134 12130 8186
rect 12142 8134 12194 8186
rect 12206 8134 12258 8186
rect 16950 8134 17002 8186
rect 17014 8134 17066 8186
rect 17078 8134 17130 8186
rect 17142 8134 17194 8186
rect 17206 8134 17258 8186
rect 21950 8134 22002 8186
rect 22014 8134 22066 8186
rect 22078 8134 22130 8186
rect 22142 8134 22194 8186
rect 22206 8134 22258 8186
rect 26950 8134 27002 8186
rect 27014 8134 27066 8186
rect 27078 8134 27130 8186
rect 27142 8134 27194 8186
rect 27206 8134 27258 8186
rect 31950 8134 32002 8186
rect 32014 8134 32066 8186
rect 32078 8134 32130 8186
rect 32142 8134 32194 8186
rect 32206 8134 32258 8186
rect 36950 8134 37002 8186
rect 37014 8134 37066 8186
rect 37078 8134 37130 8186
rect 37142 8134 37194 8186
rect 37206 8134 37258 8186
rect 26792 8032 26844 8084
rect 14648 7964 14700 8016
rect 15660 7871 15712 7880
rect 15660 7837 15669 7871
rect 15669 7837 15703 7871
rect 15703 7837 15712 7871
rect 15660 7828 15712 7837
rect 16396 7896 16448 7948
rect 30932 7964 30984 8016
rect 22468 7896 22520 7948
rect 36544 7896 36596 7948
rect 13636 7760 13688 7812
rect 22376 7760 22428 7812
rect 24860 7692 24912 7744
rect 2610 7590 2662 7642
rect 2674 7590 2726 7642
rect 2738 7590 2790 7642
rect 2802 7590 2854 7642
rect 2866 7590 2918 7642
rect 7610 7590 7662 7642
rect 7674 7590 7726 7642
rect 7738 7590 7790 7642
rect 7802 7590 7854 7642
rect 7866 7590 7918 7642
rect 12610 7590 12662 7642
rect 12674 7590 12726 7642
rect 12738 7590 12790 7642
rect 12802 7590 12854 7642
rect 12866 7590 12918 7642
rect 17610 7590 17662 7642
rect 17674 7590 17726 7642
rect 17738 7590 17790 7642
rect 17802 7590 17854 7642
rect 17866 7590 17918 7642
rect 22610 7590 22662 7642
rect 22674 7590 22726 7642
rect 22738 7590 22790 7642
rect 22802 7590 22854 7642
rect 22866 7590 22918 7642
rect 27610 7590 27662 7642
rect 27674 7590 27726 7642
rect 27738 7590 27790 7642
rect 27802 7590 27854 7642
rect 27866 7590 27918 7642
rect 32610 7590 32662 7642
rect 32674 7590 32726 7642
rect 32738 7590 32790 7642
rect 32802 7590 32854 7642
rect 32866 7590 32918 7642
rect 37610 7590 37662 7642
rect 37674 7590 37726 7642
rect 37738 7590 37790 7642
rect 37802 7590 37854 7642
rect 37866 7590 37918 7642
rect 8944 7488 8996 7540
rect 15752 7352 15804 7404
rect 19800 7395 19852 7404
rect 19800 7361 19809 7395
rect 19809 7361 19843 7395
rect 19843 7361 19852 7395
rect 19800 7352 19852 7361
rect 20076 7352 20128 7404
rect 6092 7284 6144 7336
rect 19892 7327 19944 7336
rect 19892 7293 19901 7327
rect 19901 7293 19935 7327
rect 19935 7293 19944 7327
rect 19892 7284 19944 7293
rect 24952 7284 25004 7336
rect 1950 7046 2002 7098
rect 2014 7046 2066 7098
rect 2078 7046 2130 7098
rect 2142 7046 2194 7098
rect 2206 7046 2258 7098
rect 6950 7046 7002 7098
rect 7014 7046 7066 7098
rect 7078 7046 7130 7098
rect 7142 7046 7194 7098
rect 7206 7046 7258 7098
rect 11950 7046 12002 7098
rect 12014 7046 12066 7098
rect 12078 7046 12130 7098
rect 12142 7046 12194 7098
rect 12206 7046 12258 7098
rect 16950 7046 17002 7098
rect 17014 7046 17066 7098
rect 17078 7046 17130 7098
rect 17142 7046 17194 7098
rect 17206 7046 17258 7098
rect 21950 7046 22002 7098
rect 22014 7046 22066 7098
rect 22078 7046 22130 7098
rect 22142 7046 22194 7098
rect 22206 7046 22258 7098
rect 26950 7046 27002 7098
rect 27014 7046 27066 7098
rect 27078 7046 27130 7098
rect 27142 7046 27194 7098
rect 27206 7046 27258 7098
rect 31950 7046 32002 7098
rect 32014 7046 32066 7098
rect 32078 7046 32130 7098
rect 32142 7046 32194 7098
rect 32206 7046 32258 7098
rect 36950 7046 37002 7098
rect 37014 7046 37066 7098
rect 37078 7046 37130 7098
rect 37142 7046 37194 7098
rect 37206 7046 37258 7098
rect 34520 6808 34572 6860
rect 6828 6740 6880 6792
rect 16948 6672 17000 6724
rect 21732 6672 21784 6724
rect 29644 6672 29696 6724
rect 6184 6604 6236 6656
rect 30196 6604 30248 6656
rect 34704 6715 34756 6724
rect 34704 6681 34713 6715
rect 34713 6681 34747 6715
rect 34747 6681 34756 6715
rect 34704 6672 34756 6681
rect 35532 6783 35584 6792
rect 35532 6749 35541 6783
rect 35541 6749 35575 6783
rect 35575 6749 35584 6783
rect 35532 6740 35584 6749
rect 35624 6783 35676 6792
rect 35624 6749 35633 6783
rect 35633 6749 35667 6783
rect 35667 6749 35676 6783
rect 35624 6740 35676 6749
rect 37280 6672 37332 6724
rect 35624 6604 35676 6656
rect 2610 6502 2662 6554
rect 2674 6502 2726 6554
rect 2738 6502 2790 6554
rect 2802 6502 2854 6554
rect 2866 6502 2918 6554
rect 7610 6502 7662 6554
rect 7674 6502 7726 6554
rect 7738 6502 7790 6554
rect 7802 6502 7854 6554
rect 7866 6502 7918 6554
rect 12610 6502 12662 6554
rect 12674 6502 12726 6554
rect 12738 6502 12790 6554
rect 12802 6502 12854 6554
rect 12866 6502 12918 6554
rect 17610 6502 17662 6554
rect 17674 6502 17726 6554
rect 17738 6502 17790 6554
rect 17802 6502 17854 6554
rect 17866 6502 17918 6554
rect 22610 6502 22662 6554
rect 22674 6502 22726 6554
rect 22738 6502 22790 6554
rect 22802 6502 22854 6554
rect 22866 6502 22918 6554
rect 27610 6502 27662 6554
rect 27674 6502 27726 6554
rect 27738 6502 27790 6554
rect 27802 6502 27854 6554
rect 27866 6502 27918 6554
rect 32610 6502 32662 6554
rect 32674 6502 32726 6554
rect 32738 6502 32790 6554
rect 32802 6502 32854 6554
rect 32866 6502 32918 6554
rect 37610 6502 37662 6554
rect 37674 6502 37726 6554
rect 37738 6502 37790 6554
rect 37802 6502 37854 6554
rect 37866 6502 37918 6554
rect 5724 6443 5776 6452
rect 5724 6409 5733 6443
rect 5733 6409 5767 6443
rect 5767 6409 5776 6443
rect 5724 6400 5776 6409
rect 1400 6332 1452 6384
rect 37372 6400 37424 6452
rect 6184 6307 6236 6316
rect 6184 6273 6193 6307
rect 6193 6273 6227 6307
rect 6227 6273 6236 6307
rect 6184 6264 6236 6273
rect 17500 6332 17552 6384
rect 16672 6307 16724 6316
rect 16672 6273 16681 6307
rect 16681 6273 16715 6307
rect 16715 6273 16724 6307
rect 16672 6264 16724 6273
rect 16764 6307 16816 6316
rect 16764 6273 16773 6307
rect 16773 6273 16807 6307
rect 16807 6273 16816 6307
rect 16764 6264 16816 6273
rect 16948 6307 17000 6316
rect 16948 6273 16957 6307
rect 16957 6273 16991 6307
rect 16991 6273 17000 6307
rect 16948 6264 17000 6273
rect 25228 6264 25280 6316
rect 31208 6307 31260 6316
rect 31208 6273 31217 6307
rect 31217 6273 31251 6307
rect 31251 6273 31260 6307
rect 31208 6264 31260 6273
rect 31668 6264 31720 6316
rect 31852 6307 31904 6316
rect 31852 6273 31861 6307
rect 31861 6273 31895 6307
rect 31895 6273 31904 6307
rect 31852 6264 31904 6273
rect 18788 6196 18840 6248
rect 34152 6196 34204 6248
rect 29552 6128 29604 6180
rect 1950 5958 2002 6010
rect 2014 5958 2066 6010
rect 2078 5958 2130 6010
rect 2142 5958 2194 6010
rect 2206 5958 2258 6010
rect 6950 5958 7002 6010
rect 7014 5958 7066 6010
rect 7078 5958 7130 6010
rect 7142 5958 7194 6010
rect 7206 5958 7258 6010
rect 11950 5958 12002 6010
rect 12014 5958 12066 6010
rect 12078 5958 12130 6010
rect 12142 5958 12194 6010
rect 12206 5958 12258 6010
rect 16950 5958 17002 6010
rect 17014 5958 17066 6010
rect 17078 5958 17130 6010
rect 17142 5958 17194 6010
rect 17206 5958 17258 6010
rect 21950 5958 22002 6010
rect 22014 5958 22066 6010
rect 22078 5958 22130 6010
rect 22142 5958 22194 6010
rect 22206 5958 22258 6010
rect 26950 5958 27002 6010
rect 27014 5958 27066 6010
rect 27078 5958 27130 6010
rect 27142 5958 27194 6010
rect 27206 5958 27258 6010
rect 31950 5958 32002 6010
rect 32014 5958 32066 6010
rect 32078 5958 32130 6010
rect 32142 5958 32194 6010
rect 32206 5958 32258 6010
rect 36950 5958 37002 6010
rect 37014 5958 37066 6010
rect 37078 5958 37130 6010
rect 37142 5958 37194 6010
rect 37206 5958 37258 6010
rect 2610 5414 2662 5466
rect 2674 5414 2726 5466
rect 2738 5414 2790 5466
rect 2802 5414 2854 5466
rect 2866 5414 2918 5466
rect 7610 5414 7662 5466
rect 7674 5414 7726 5466
rect 7738 5414 7790 5466
rect 7802 5414 7854 5466
rect 7866 5414 7918 5466
rect 12610 5414 12662 5466
rect 12674 5414 12726 5466
rect 12738 5414 12790 5466
rect 12802 5414 12854 5466
rect 12866 5414 12918 5466
rect 17610 5414 17662 5466
rect 17674 5414 17726 5466
rect 17738 5414 17790 5466
rect 17802 5414 17854 5466
rect 17866 5414 17918 5466
rect 22610 5414 22662 5466
rect 22674 5414 22726 5466
rect 22738 5414 22790 5466
rect 22802 5414 22854 5466
rect 22866 5414 22918 5466
rect 27610 5414 27662 5466
rect 27674 5414 27726 5466
rect 27738 5414 27790 5466
rect 27802 5414 27854 5466
rect 27866 5414 27918 5466
rect 32610 5414 32662 5466
rect 32674 5414 32726 5466
rect 32738 5414 32790 5466
rect 32802 5414 32854 5466
rect 32866 5414 32918 5466
rect 37610 5414 37662 5466
rect 37674 5414 37726 5466
rect 37738 5414 37790 5466
rect 37802 5414 37854 5466
rect 37866 5414 37918 5466
rect 3700 5312 3752 5364
rect 12532 5312 12584 5364
rect 12992 5312 13044 5364
rect 8392 5287 8444 5296
rect 8392 5253 8401 5287
rect 8401 5253 8435 5287
rect 8435 5253 8444 5287
rect 8392 5244 8444 5253
rect 8208 5219 8260 5228
rect 8208 5185 8217 5219
rect 8217 5185 8251 5219
rect 8251 5185 8260 5219
rect 8208 5176 8260 5185
rect 8484 5219 8536 5228
rect 8484 5185 8493 5219
rect 8493 5185 8527 5219
rect 8527 5185 8536 5219
rect 8484 5176 8536 5185
rect 7288 5108 7340 5160
rect 22468 5176 22520 5228
rect 8760 5083 8812 5092
rect 8760 5049 8769 5083
rect 8769 5049 8803 5083
rect 8803 5049 8812 5083
rect 8760 5040 8812 5049
rect 4344 4972 4396 5024
rect 8116 4972 8168 5024
rect 19616 5040 19668 5092
rect 31024 4972 31076 5024
rect 37464 4972 37516 5024
rect 38568 4972 38620 5024
rect 1950 4870 2002 4922
rect 2014 4870 2066 4922
rect 2078 4870 2130 4922
rect 2142 4870 2194 4922
rect 2206 4870 2258 4922
rect 6950 4870 7002 4922
rect 7014 4870 7066 4922
rect 7078 4870 7130 4922
rect 7142 4870 7194 4922
rect 7206 4870 7258 4922
rect 11950 4870 12002 4922
rect 12014 4870 12066 4922
rect 12078 4870 12130 4922
rect 12142 4870 12194 4922
rect 12206 4870 12258 4922
rect 16950 4870 17002 4922
rect 17014 4870 17066 4922
rect 17078 4870 17130 4922
rect 17142 4870 17194 4922
rect 17206 4870 17258 4922
rect 21950 4870 22002 4922
rect 22014 4870 22066 4922
rect 22078 4870 22130 4922
rect 22142 4870 22194 4922
rect 22206 4870 22258 4922
rect 26950 4870 27002 4922
rect 27014 4870 27066 4922
rect 27078 4870 27130 4922
rect 27142 4870 27194 4922
rect 27206 4870 27258 4922
rect 31950 4870 32002 4922
rect 32014 4870 32066 4922
rect 32078 4870 32130 4922
rect 32142 4870 32194 4922
rect 32206 4870 32258 4922
rect 36950 4870 37002 4922
rect 37014 4870 37066 4922
rect 37078 4870 37130 4922
rect 37142 4870 37194 4922
rect 37206 4870 37258 4922
rect 7380 4768 7432 4820
rect 3700 4632 3752 4684
rect 3792 4675 3844 4684
rect 3792 4641 3801 4675
rect 3801 4641 3835 4675
rect 3835 4641 3844 4675
rect 3792 4632 3844 4641
rect 8392 4700 8444 4752
rect 31024 4768 31076 4820
rect 35624 4768 35676 4820
rect 848 4564 900 4616
rect 4344 4607 4396 4616
rect 4344 4573 4353 4607
rect 4353 4573 4387 4607
rect 4387 4573 4396 4607
rect 4344 4564 4396 4573
rect 6092 4564 6144 4616
rect 7472 4632 7524 4684
rect 14096 4675 14148 4684
rect 14096 4641 14105 4675
rect 14105 4641 14139 4675
rect 14139 4641 14148 4675
rect 14096 4632 14148 4641
rect 7012 4607 7064 4616
rect 7012 4573 7021 4607
rect 7021 4573 7055 4607
rect 7055 4573 7064 4607
rect 7012 4564 7064 4573
rect 8208 4564 8260 4616
rect 14280 4607 14332 4616
rect 14280 4573 14289 4607
rect 14289 4573 14323 4607
rect 14323 4573 14332 4607
rect 14280 4564 14332 4573
rect 6276 4496 6328 4548
rect 18604 4564 18656 4616
rect 19524 4607 19576 4616
rect 19524 4573 19533 4607
rect 19533 4573 19567 4607
rect 19567 4573 19576 4607
rect 19524 4564 19576 4573
rect 19984 4675 20036 4684
rect 19984 4641 19993 4675
rect 19993 4641 20027 4675
rect 20027 4641 20036 4675
rect 19984 4632 20036 4641
rect 26424 4632 26476 4684
rect 34704 4564 34756 4616
rect 37372 4675 37424 4684
rect 37372 4641 37381 4675
rect 37381 4641 37415 4675
rect 37415 4641 37424 4675
rect 37372 4632 37424 4641
rect 38108 4632 38160 4684
rect 38568 4743 38620 4752
rect 38568 4709 38577 4743
rect 38577 4709 38611 4743
rect 38611 4709 38620 4743
rect 38568 4700 38620 4709
rect 18236 4496 18288 4548
rect 19616 4539 19668 4548
rect 19616 4505 19625 4539
rect 19625 4505 19659 4539
rect 19659 4505 19668 4539
rect 19616 4496 19668 4505
rect 37280 4496 37332 4548
rect 7288 4428 7340 4480
rect 35532 4428 35584 4480
rect 2610 4326 2662 4378
rect 2674 4326 2726 4378
rect 2738 4326 2790 4378
rect 2802 4326 2854 4378
rect 2866 4326 2918 4378
rect 7610 4326 7662 4378
rect 7674 4326 7726 4378
rect 7738 4326 7790 4378
rect 7802 4326 7854 4378
rect 7866 4326 7918 4378
rect 12610 4326 12662 4378
rect 12674 4326 12726 4378
rect 12738 4326 12790 4378
rect 12802 4326 12854 4378
rect 12866 4326 12918 4378
rect 17610 4326 17662 4378
rect 17674 4326 17726 4378
rect 17738 4326 17790 4378
rect 17802 4326 17854 4378
rect 17866 4326 17918 4378
rect 22610 4326 22662 4378
rect 22674 4326 22726 4378
rect 22738 4326 22790 4378
rect 22802 4326 22854 4378
rect 22866 4326 22918 4378
rect 27610 4326 27662 4378
rect 27674 4326 27726 4378
rect 27738 4326 27790 4378
rect 27802 4326 27854 4378
rect 27866 4326 27918 4378
rect 32610 4326 32662 4378
rect 32674 4326 32726 4378
rect 32738 4326 32790 4378
rect 32802 4326 32854 4378
rect 32866 4326 32918 4378
rect 37610 4326 37662 4378
rect 37674 4326 37726 4378
rect 37738 4326 37790 4378
rect 37802 4326 37854 4378
rect 37866 4326 37918 4378
rect 40500 4199 40552 4208
rect 40500 4165 40509 4199
rect 40509 4165 40543 4199
rect 40543 4165 40552 4199
rect 40500 4156 40552 4165
rect 6460 4131 6512 4140
rect 6460 4097 6469 4131
rect 6469 4097 6503 4131
rect 6503 4097 6512 4131
rect 6460 4088 6512 4097
rect 9220 4088 9272 4140
rect 34152 4131 34204 4140
rect 34152 4097 34161 4131
rect 34161 4097 34195 4131
rect 34195 4097 34204 4131
rect 34152 4088 34204 4097
rect 8852 4020 8904 4072
rect 36820 4020 36872 4072
rect 1950 3782 2002 3834
rect 2014 3782 2066 3834
rect 2078 3782 2130 3834
rect 2142 3782 2194 3834
rect 2206 3782 2258 3834
rect 6950 3782 7002 3834
rect 7014 3782 7066 3834
rect 7078 3782 7130 3834
rect 7142 3782 7194 3834
rect 7206 3782 7258 3834
rect 11950 3782 12002 3834
rect 12014 3782 12066 3834
rect 12078 3782 12130 3834
rect 12142 3782 12194 3834
rect 12206 3782 12258 3834
rect 16950 3782 17002 3834
rect 17014 3782 17066 3834
rect 17078 3782 17130 3834
rect 17142 3782 17194 3834
rect 17206 3782 17258 3834
rect 21950 3782 22002 3834
rect 22014 3782 22066 3834
rect 22078 3782 22130 3834
rect 22142 3782 22194 3834
rect 22206 3782 22258 3834
rect 26950 3782 27002 3834
rect 27014 3782 27066 3834
rect 27078 3782 27130 3834
rect 27142 3782 27194 3834
rect 27206 3782 27258 3834
rect 31950 3782 32002 3834
rect 32014 3782 32066 3834
rect 32078 3782 32130 3834
rect 32142 3782 32194 3834
rect 32206 3782 32258 3834
rect 36950 3782 37002 3834
rect 37014 3782 37066 3834
rect 37078 3782 37130 3834
rect 37142 3782 37194 3834
rect 37206 3782 37258 3834
rect 4804 3476 4856 3528
rect 10968 3655 11020 3664
rect 10968 3621 10977 3655
rect 10977 3621 11011 3655
rect 11011 3621 11020 3655
rect 10968 3612 11020 3621
rect 34152 3723 34204 3732
rect 34152 3689 34161 3723
rect 34161 3689 34195 3723
rect 34195 3689 34204 3723
rect 34152 3680 34204 3689
rect 33692 3612 33744 3664
rect 10876 3544 10928 3596
rect 8024 3408 8076 3460
rect 11152 3519 11204 3528
rect 11152 3485 11161 3519
rect 11161 3485 11195 3519
rect 11195 3485 11204 3519
rect 11152 3476 11204 3485
rect 12532 3476 12584 3528
rect 35900 3544 35952 3596
rect 36820 3544 36872 3596
rect 8208 3383 8260 3392
rect 8208 3349 8217 3383
rect 8217 3349 8251 3383
rect 8251 3349 8260 3383
rect 14464 3476 14516 3528
rect 8208 3340 8260 3349
rect 26056 3340 26108 3392
rect 29644 3340 29696 3392
rect 2610 3238 2662 3290
rect 2674 3238 2726 3290
rect 2738 3238 2790 3290
rect 2802 3238 2854 3290
rect 2866 3238 2918 3290
rect 7610 3238 7662 3290
rect 7674 3238 7726 3290
rect 7738 3238 7790 3290
rect 7802 3238 7854 3290
rect 7866 3238 7918 3290
rect 12610 3238 12662 3290
rect 12674 3238 12726 3290
rect 12738 3238 12790 3290
rect 12802 3238 12854 3290
rect 12866 3238 12918 3290
rect 17610 3238 17662 3290
rect 17674 3238 17726 3290
rect 17738 3238 17790 3290
rect 17802 3238 17854 3290
rect 17866 3238 17918 3290
rect 22610 3238 22662 3290
rect 22674 3238 22726 3290
rect 22738 3238 22790 3290
rect 22802 3238 22854 3290
rect 22866 3238 22918 3290
rect 27610 3238 27662 3290
rect 27674 3238 27726 3290
rect 27738 3238 27790 3290
rect 27802 3238 27854 3290
rect 27866 3238 27918 3290
rect 32610 3238 32662 3290
rect 32674 3238 32726 3290
rect 32738 3238 32790 3290
rect 32802 3238 32854 3290
rect 32866 3238 32918 3290
rect 37610 3238 37662 3290
rect 37674 3238 37726 3290
rect 37738 3238 37790 3290
rect 37802 3238 37854 3290
rect 37866 3238 37918 3290
rect 8484 3136 8536 3188
rect 27528 3136 27580 3188
rect 34152 3179 34204 3188
rect 34152 3145 34161 3179
rect 34161 3145 34195 3179
rect 34195 3145 34204 3179
rect 34152 3136 34204 3145
rect 28172 3043 28224 3052
rect 28172 3009 28181 3043
rect 28181 3009 28215 3043
rect 28215 3009 28224 3043
rect 28172 3000 28224 3009
rect 20076 2932 20128 2984
rect 27988 2932 28040 2984
rect 29644 3111 29696 3120
rect 29644 3077 29653 3111
rect 29653 3077 29687 3111
rect 29687 3077 29696 3111
rect 29644 3068 29696 3077
rect 28632 3043 28684 3052
rect 28632 3009 28641 3043
rect 28641 3009 28675 3043
rect 28675 3009 28684 3043
rect 28632 3000 28684 3009
rect 33232 3000 33284 3052
rect 26332 2864 26384 2916
rect 17316 2796 17368 2848
rect 1950 2694 2002 2746
rect 2014 2694 2066 2746
rect 2078 2694 2130 2746
rect 2142 2694 2194 2746
rect 2206 2694 2258 2746
rect 6950 2694 7002 2746
rect 7014 2694 7066 2746
rect 7078 2694 7130 2746
rect 7142 2694 7194 2746
rect 7206 2694 7258 2746
rect 11950 2694 12002 2746
rect 12014 2694 12066 2746
rect 12078 2694 12130 2746
rect 12142 2694 12194 2746
rect 12206 2694 12258 2746
rect 16950 2694 17002 2746
rect 17014 2694 17066 2746
rect 17078 2694 17130 2746
rect 17142 2694 17194 2746
rect 17206 2694 17258 2746
rect 21950 2694 22002 2746
rect 22014 2694 22066 2746
rect 22078 2694 22130 2746
rect 22142 2694 22194 2746
rect 22206 2694 22258 2746
rect 26950 2694 27002 2746
rect 27014 2694 27066 2746
rect 27078 2694 27130 2746
rect 27142 2694 27194 2746
rect 27206 2694 27258 2746
rect 31950 2694 32002 2746
rect 32014 2694 32066 2746
rect 32078 2694 32130 2746
rect 32142 2694 32194 2746
rect 32206 2694 32258 2746
rect 36950 2694 37002 2746
rect 37014 2694 37066 2746
rect 37078 2694 37130 2746
rect 37142 2694 37194 2746
rect 37206 2694 37258 2746
rect 2504 2499 2556 2508
rect 2504 2465 2513 2499
rect 2513 2465 2547 2499
rect 2547 2465 2556 2499
rect 2504 2456 2556 2465
rect 11704 2456 11756 2508
rect 10140 2388 10192 2440
rect 24584 2592 24636 2644
rect 14372 2524 14424 2576
rect 34612 2456 34664 2508
rect 8024 2320 8076 2372
rect 34152 2431 34204 2440
rect 34152 2397 34161 2431
rect 34161 2397 34195 2431
rect 34195 2397 34204 2431
rect 34152 2388 34204 2397
rect 2320 2252 2372 2304
rect 28632 2363 28684 2372
rect 28632 2329 28641 2363
rect 28641 2329 28675 2363
rect 28675 2329 28684 2363
rect 28632 2320 28684 2329
rect 13084 2252 13136 2304
rect 18328 2252 18380 2304
rect 23572 2252 23624 2304
rect 28816 2252 28868 2304
rect 34060 2252 34112 2304
rect 39304 2252 39356 2304
rect 2610 2150 2662 2202
rect 2674 2150 2726 2202
rect 2738 2150 2790 2202
rect 2802 2150 2854 2202
rect 2866 2150 2918 2202
rect 7610 2150 7662 2202
rect 7674 2150 7726 2202
rect 7738 2150 7790 2202
rect 7802 2150 7854 2202
rect 7866 2150 7918 2202
rect 12610 2150 12662 2202
rect 12674 2150 12726 2202
rect 12738 2150 12790 2202
rect 12802 2150 12854 2202
rect 12866 2150 12918 2202
rect 17610 2150 17662 2202
rect 17674 2150 17726 2202
rect 17738 2150 17790 2202
rect 17802 2150 17854 2202
rect 17866 2150 17918 2202
rect 22610 2150 22662 2202
rect 22674 2150 22726 2202
rect 22738 2150 22790 2202
rect 22802 2150 22854 2202
rect 22866 2150 22918 2202
rect 27610 2150 27662 2202
rect 27674 2150 27726 2202
rect 27738 2150 27790 2202
rect 27802 2150 27854 2202
rect 27866 2150 27918 2202
rect 32610 2150 32662 2202
rect 32674 2150 32726 2202
rect 32738 2150 32790 2202
rect 32802 2150 32854 2202
rect 32866 2150 32918 2202
rect 37610 2150 37662 2202
rect 37674 2150 37726 2202
rect 37738 2150 37790 2202
rect 37802 2150 37854 2202
rect 37866 2150 37918 2202
<< metal2 >>
rect 6918 71346 6974 72000
rect 6918 71318 7144 71346
rect 6918 71200 6974 71318
rect 2610 69660 2918 69669
rect 2610 69658 2616 69660
rect 2672 69658 2696 69660
rect 2752 69658 2776 69660
rect 2832 69658 2856 69660
rect 2912 69658 2918 69660
rect 2672 69606 2674 69658
rect 2854 69606 2856 69658
rect 2610 69604 2616 69606
rect 2672 69604 2696 69606
rect 2752 69604 2776 69606
rect 2832 69604 2856 69606
rect 2912 69604 2918 69606
rect 2610 69595 2918 69604
rect 7116 69426 7144 71318
rect 20902 71200 20958 72000
rect 34886 71346 34942 72000
rect 34886 71318 35020 71346
rect 34886 71200 34942 71318
rect 7610 69660 7918 69669
rect 7610 69658 7616 69660
rect 7672 69658 7696 69660
rect 7752 69658 7776 69660
rect 7832 69658 7856 69660
rect 7912 69658 7918 69660
rect 7672 69606 7674 69658
rect 7854 69606 7856 69658
rect 7610 69604 7616 69606
rect 7672 69604 7696 69606
rect 7752 69604 7776 69606
rect 7832 69604 7856 69606
rect 7912 69604 7918 69606
rect 7610 69595 7918 69604
rect 12610 69660 12918 69669
rect 12610 69658 12616 69660
rect 12672 69658 12696 69660
rect 12752 69658 12776 69660
rect 12832 69658 12856 69660
rect 12912 69658 12918 69660
rect 12672 69606 12674 69658
rect 12854 69606 12856 69658
rect 12610 69604 12616 69606
rect 12672 69604 12696 69606
rect 12752 69604 12776 69606
rect 12832 69604 12856 69606
rect 12912 69604 12918 69606
rect 12610 69595 12918 69604
rect 17610 69660 17918 69669
rect 17610 69658 17616 69660
rect 17672 69658 17696 69660
rect 17752 69658 17776 69660
rect 17832 69658 17856 69660
rect 17912 69658 17918 69660
rect 17672 69606 17674 69658
rect 17854 69606 17856 69658
rect 17610 69604 17616 69606
rect 17672 69604 17696 69606
rect 17752 69604 17776 69606
rect 17832 69604 17856 69606
rect 17912 69604 17918 69606
rect 17610 69595 17918 69604
rect 20916 69426 20944 71200
rect 22610 69660 22918 69669
rect 22610 69658 22616 69660
rect 22672 69658 22696 69660
rect 22752 69658 22776 69660
rect 22832 69658 22856 69660
rect 22912 69658 22918 69660
rect 22672 69606 22674 69658
rect 22854 69606 22856 69658
rect 22610 69604 22616 69606
rect 22672 69604 22696 69606
rect 22752 69604 22776 69606
rect 22832 69604 22856 69606
rect 22912 69604 22918 69606
rect 22610 69595 22918 69604
rect 27610 69660 27918 69669
rect 27610 69658 27616 69660
rect 27672 69658 27696 69660
rect 27752 69658 27776 69660
rect 27832 69658 27856 69660
rect 27912 69658 27918 69660
rect 27672 69606 27674 69658
rect 27854 69606 27856 69658
rect 27610 69604 27616 69606
rect 27672 69604 27696 69606
rect 27752 69604 27776 69606
rect 27832 69604 27856 69606
rect 27912 69604 27918 69606
rect 27610 69595 27918 69604
rect 32610 69660 32918 69669
rect 32610 69658 32616 69660
rect 32672 69658 32696 69660
rect 32752 69658 32776 69660
rect 32832 69658 32856 69660
rect 32912 69658 32918 69660
rect 32672 69606 32674 69658
rect 32854 69606 32856 69658
rect 32610 69604 32616 69606
rect 32672 69604 32696 69606
rect 32752 69604 32776 69606
rect 32832 69604 32856 69606
rect 32912 69604 32918 69606
rect 32610 69595 32918 69604
rect 34992 69494 35020 71318
rect 37610 69660 37918 69669
rect 37610 69658 37616 69660
rect 37672 69658 37696 69660
rect 37752 69658 37776 69660
rect 37832 69658 37856 69660
rect 37912 69658 37918 69660
rect 37672 69606 37674 69658
rect 37854 69606 37856 69658
rect 37610 69604 37616 69606
rect 37672 69604 37696 69606
rect 37752 69604 37776 69606
rect 37832 69604 37856 69606
rect 37912 69604 37918 69606
rect 37610 69595 37918 69604
rect 34980 69488 35032 69494
rect 34980 69430 35032 69436
rect 7104 69420 7156 69426
rect 7104 69362 7156 69368
rect 20904 69420 20956 69426
rect 20904 69362 20956 69368
rect 9588 69352 9640 69358
rect 9588 69294 9640 69300
rect 22376 69352 22428 69358
rect 22376 69294 22428 69300
rect 35440 69352 35492 69358
rect 35440 69294 35492 69300
rect 1950 69116 2258 69125
rect 1950 69114 1956 69116
rect 2012 69114 2036 69116
rect 2092 69114 2116 69116
rect 2172 69114 2196 69116
rect 2252 69114 2258 69116
rect 2012 69062 2014 69114
rect 2194 69062 2196 69114
rect 1950 69060 1956 69062
rect 2012 69060 2036 69062
rect 2092 69060 2116 69062
rect 2172 69060 2196 69062
rect 2252 69060 2258 69062
rect 1950 69051 2258 69060
rect 6950 69116 7258 69125
rect 6950 69114 6956 69116
rect 7012 69114 7036 69116
rect 7092 69114 7116 69116
rect 7172 69114 7196 69116
rect 7252 69114 7258 69116
rect 7012 69062 7014 69114
rect 7194 69062 7196 69114
rect 6950 69060 6956 69062
rect 7012 69060 7036 69062
rect 7092 69060 7116 69062
rect 7172 69060 7196 69062
rect 7252 69060 7258 69062
rect 6950 69051 7258 69060
rect 2610 68572 2918 68581
rect 2610 68570 2616 68572
rect 2672 68570 2696 68572
rect 2752 68570 2776 68572
rect 2832 68570 2856 68572
rect 2912 68570 2918 68572
rect 2672 68518 2674 68570
rect 2854 68518 2856 68570
rect 2610 68516 2616 68518
rect 2672 68516 2696 68518
rect 2752 68516 2776 68518
rect 2832 68516 2856 68518
rect 2912 68516 2918 68518
rect 2610 68507 2918 68516
rect 7610 68572 7918 68581
rect 7610 68570 7616 68572
rect 7672 68570 7696 68572
rect 7752 68570 7776 68572
rect 7832 68570 7856 68572
rect 7912 68570 7918 68572
rect 7672 68518 7674 68570
rect 7854 68518 7856 68570
rect 7610 68516 7616 68518
rect 7672 68516 7696 68518
rect 7752 68516 7776 68518
rect 7832 68516 7856 68518
rect 7912 68516 7918 68518
rect 7610 68507 7918 68516
rect 1950 68028 2258 68037
rect 1950 68026 1956 68028
rect 2012 68026 2036 68028
rect 2092 68026 2116 68028
rect 2172 68026 2196 68028
rect 2252 68026 2258 68028
rect 2012 67974 2014 68026
rect 2194 67974 2196 68026
rect 1950 67972 1956 67974
rect 2012 67972 2036 67974
rect 2092 67972 2116 67974
rect 2172 67972 2196 67974
rect 2252 67972 2258 67974
rect 1950 67963 2258 67972
rect 6950 68028 7258 68037
rect 6950 68026 6956 68028
rect 7012 68026 7036 68028
rect 7092 68026 7116 68028
rect 7172 68026 7196 68028
rect 7252 68026 7258 68028
rect 7012 67974 7014 68026
rect 7194 67974 7196 68026
rect 6950 67972 6956 67974
rect 7012 67972 7036 67974
rect 7092 67972 7116 67974
rect 7172 67972 7196 67974
rect 7252 67972 7258 67974
rect 6950 67963 7258 67972
rect 8944 67924 8996 67930
rect 8944 67866 8996 67872
rect 1400 67720 1452 67726
rect 1400 67662 1452 67668
rect 1412 67289 1440 67662
rect 6552 67652 6604 67658
rect 6552 67594 6604 67600
rect 2610 67484 2918 67493
rect 2610 67482 2616 67484
rect 2672 67482 2696 67484
rect 2752 67482 2776 67484
rect 2832 67482 2856 67484
rect 2912 67482 2918 67484
rect 2672 67430 2674 67482
rect 2854 67430 2856 67482
rect 2610 67428 2616 67430
rect 2672 67428 2696 67430
rect 2752 67428 2776 67430
rect 2832 67428 2856 67430
rect 2912 67428 2918 67430
rect 2610 67419 2918 67428
rect 1398 67280 1454 67289
rect 1398 67215 1454 67224
rect 1950 66940 2258 66949
rect 1950 66938 1956 66940
rect 2012 66938 2036 66940
rect 2092 66938 2116 66940
rect 2172 66938 2196 66940
rect 2252 66938 2258 66940
rect 2012 66886 2014 66938
rect 2194 66886 2196 66938
rect 1950 66884 1956 66886
rect 2012 66884 2036 66886
rect 2092 66884 2116 66886
rect 2172 66884 2196 66886
rect 2252 66884 2258 66886
rect 1950 66875 2258 66884
rect 2610 66396 2918 66405
rect 2610 66394 2616 66396
rect 2672 66394 2696 66396
rect 2752 66394 2776 66396
rect 2832 66394 2856 66396
rect 2912 66394 2918 66396
rect 2672 66342 2674 66394
rect 2854 66342 2856 66394
rect 2610 66340 2616 66342
rect 2672 66340 2696 66342
rect 2752 66340 2776 66342
rect 2832 66340 2856 66342
rect 2912 66340 2918 66342
rect 2610 66331 2918 66340
rect 4528 66156 4580 66162
rect 4528 66098 4580 66104
rect 6460 66156 6512 66162
rect 6460 66098 6512 66104
rect 1950 65852 2258 65861
rect 1950 65850 1956 65852
rect 2012 65850 2036 65852
rect 2092 65850 2116 65852
rect 2172 65850 2196 65852
rect 2252 65850 2258 65852
rect 2012 65798 2014 65850
rect 2194 65798 2196 65850
rect 1950 65796 1956 65798
rect 2012 65796 2036 65798
rect 2092 65796 2116 65798
rect 2172 65796 2196 65798
rect 2252 65796 2258 65798
rect 1950 65787 2258 65796
rect 2964 65612 3016 65618
rect 2964 65554 3016 65560
rect 1584 65476 1636 65482
rect 1584 65418 1636 65424
rect 848 58540 900 58546
rect 848 58482 900 58488
rect 860 58449 888 58482
rect 846 58440 902 58449
rect 846 58375 902 58384
rect 1400 49836 1452 49842
rect 1400 49778 1452 49784
rect 1412 49337 1440 49778
rect 1398 49328 1454 49337
rect 1398 49263 1454 49272
rect 846 40216 902 40225
rect 846 40151 902 40160
rect 860 40118 888 40151
rect 848 40112 900 40118
rect 848 40054 900 40060
rect 1400 31816 1452 31822
rect 1400 31758 1452 31764
rect 1412 31385 1440 31758
rect 1398 31376 1454 31385
rect 1398 31311 1454 31320
rect 1492 30660 1544 30666
rect 1492 30602 1544 30608
rect 848 22636 900 22642
rect 848 22578 900 22584
rect 860 22545 888 22578
rect 846 22536 902 22545
rect 846 22471 902 22480
rect 1400 13932 1452 13938
rect 1400 13874 1452 13880
rect 1412 13433 1440 13874
rect 1398 13424 1454 13433
rect 1398 13359 1454 13368
rect 1504 6914 1532 30602
rect 1596 20534 1624 65418
rect 2610 65308 2918 65317
rect 2610 65306 2616 65308
rect 2672 65306 2696 65308
rect 2752 65306 2776 65308
rect 2832 65306 2856 65308
rect 2912 65306 2918 65308
rect 2672 65254 2674 65306
rect 2854 65254 2856 65306
rect 2610 65252 2616 65254
rect 2672 65252 2696 65254
rect 2752 65252 2776 65254
rect 2832 65252 2856 65254
rect 2912 65252 2918 65254
rect 2610 65243 2918 65252
rect 1950 64764 2258 64773
rect 1950 64762 1956 64764
rect 2012 64762 2036 64764
rect 2092 64762 2116 64764
rect 2172 64762 2196 64764
rect 2252 64762 2258 64764
rect 2012 64710 2014 64762
rect 2194 64710 2196 64762
rect 1950 64708 1956 64710
rect 2012 64708 2036 64710
rect 2092 64708 2116 64710
rect 2172 64708 2196 64710
rect 2252 64708 2258 64710
rect 1950 64699 2258 64708
rect 2610 64220 2918 64229
rect 2610 64218 2616 64220
rect 2672 64218 2696 64220
rect 2752 64218 2776 64220
rect 2832 64218 2856 64220
rect 2912 64218 2918 64220
rect 2672 64166 2674 64218
rect 2854 64166 2856 64218
rect 2610 64164 2616 64166
rect 2672 64164 2696 64166
rect 2752 64164 2776 64166
rect 2832 64164 2856 64166
rect 2912 64164 2918 64166
rect 2610 64155 2918 64164
rect 1950 63676 2258 63685
rect 1950 63674 1956 63676
rect 2012 63674 2036 63676
rect 2092 63674 2116 63676
rect 2172 63674 2196 63676
rect 2252 63674 2258 63676
rect 2012 63622 2014 63674
rect 2194 63622 2196 63674
rect 1950 63620 1956 63622
rect 2012 63620 2036 63622
rect 2092 63620 2116 63622
rect 2172 63620 2196 63622
rect 2252 63620 2258 63622
rect 1950 63611 2258 63620
rect 2610 63132 2918 63141
rect 2610 63130 2616 63132
rect 2672 63130 2696 63132
rect 2752 63130 2776 63132
rect 2832 63130 2856 63132
rect 2912 63130 2918 63132
rect 2672 63078 2674 63130
rect 2854 63078 2856 63130
rect 2610 63076 2616 63078
rect 2672 63076 2696 63078
rect 2752 63076 2776 63078
rect 2832 63076 2856 63078
rect 2912 63076 2918 63078
rect 2610 63067 2918 63076
rect 1860 62824 1912 62830
rect 1860 62766 1912 62772
rect 1676 60716 1728 60722
rect 1676 60658 1728 60664
rect 1688 31822 1716 60658
rect 1768 40520 1820 40526
rect 1768 40462 1820 40468
rect 1780 33998 1808 40462
rect 1768 33992 1820 33998
rect 1768 33934 1820 33940
rect 1676 31816 1728 31822
rect 1676 31758 1728 31764
rect 1688 25974 1716 31758
rect 1676 25968 1728 25974
rect 1676 25910 1728 25916
rect 1676 24336 1728 24342
rect 1676 24278 1728 24284
rect 1688 20602 1716 24278
rect 1780 24274 1808 33934
rect 1872 30734 1900 62766
rect 1950 62588 2258 62597
rect 1950 62586 1956 62588
rect 2012 62586 2036 62588
rect 2092 62586 2116 62588
rect 2172 62586 2196 62588
rect 2252 62586 2258 62588
rect 2012 62534 2014 62586
rect 2194 62534 2196 62586
rect 1950 62532 1956 62534
rect 2012 62532 2036 62534
rect 2092 62532 2116 62534
rect 2172 62532 2196 62534
rect 2252 62532 2258 62534
rect 1950 62523 2258 62532
rect 2610 62044 2918 62053
rect 2610 62042 2616 62044
rect 2672 62042 2696 62044
rect 2752 62042 2776 62044
rect 2832 62042 2856 62044
rect 2912 62042 2918 62044
rect 2672 61990 2674 62042
rect 2854 61990 2856 62042
rect 2610 61988 2616 61990
rect 2672 61988 2696 61990
rect 2752 61988 2776 61990
rect 2832 61988 2856 61990
rect 2912 61988 2918 61990
rect 2610 61979 2918 61988
rect 1950 61500 2258 61509
rect 1950 61498 1956 61500
rect 2012 61498 2036 61500
rect 2092 61498 2116 61500
rect 2172 61498 2196 61500
rect 2252 61498 2258 61500
rect 2012 61446 2014 61498
rect 2194 61446 2196 61498
rect 1950 61444 1956 61446
rect 2012 61444 2036 61446
rect 2092 61444 2116 61446
rect 2172 61444 2196 61446
rect 2252 61444 2258 61446
rect 1950 61435 2258 61444
rect 2504 61192 2556 61198
rect 2504 61134 2556 61140
rect 2320 61124 2372 61130
rect 2320 61066 2372 61072
rect 1950 60412 2258 60421
rect 1950 60410 1956 60412
rect 2012 60410 2036 60412
rect 2092 60410 2116 60412
rect 2172 60410 2196 60412
rect 2252 60410 2258 60412
rect 2012 60358 2014 60410
rect 2194 60358 2196 60410
rect 1950 60356 1956 60358
rect 2012 60356 2036 60358
rect 2092 60356 2116 60358
rect 2172 60356 2196 60358
rect 2252 60356 2258 60358
rect 1950 60347 2258 60356
rect 1950 59324 2258 59333
rect 1950 59322 1956 59324
rect 2012 59322 2036 59324
rect 2092 59322 2116 59324
rect 2172 59322 2196 59324
rect 2252 59322 2258 59324
rect 2012 59270 2014 59322
rect 2194 59270 2196 59322
rect 1950 59268 1956 59270
rect 2012 59268 2036 59270
rect 2092 59268 2116 59270
rect 2172 59268 2196 59270
rect 2252 59268 2258 59270
rect 1950 59259 2258 59268
rect 1950 58236 2258 58245
rect 1950 58234 1956 58236
rect 2012 58234 2036 58236
rect 2092 58234 2116 58236
rect 2172 58234 2196 58236
rect 2252 58234 2258 58236
rect 2012 58182 2014 58234
rect 2194 58182 2196 58234
rect 1950 58180 1956 58182
rect 2012 58180 2036 58182
rect 2092 58180 2116 58182
rect 2172 58180 2196 58182
rect 2252 58180 2258 58182
rect 1950 58171 2258 58180
rect 2332 57254 2360 61066
rect 2320 57248 2372 57254
rect 2320 57190 2372 57196
rect 1950 57148 2258 57157
rect 1950 57146 1956 57148
rect 2012 57146 2036 57148
rect 2092 57146 2116 57148
rect 2172 57146 2196 57148
rect 2252 57146 2258 57148
rect 2012 57094 2014 57146
rect 2194 57094 2196 57146
rect 1950 57092 1956 57094
rect 2012 57092 2036 57094
rect 2092 57092 2116 57094
rect 2172 57092 2196 57094
rect 2252 57092 2258 57094
rect 1950 57083 2258 57092
rect 1950 56060 2258 56069
rect 1950 56058 1956 56060
rect 2012 56058 2036 56060
rect 2092 56058 2116 56060
rect 2172 56058 2196 56060
rect 2252 56058 2258 56060
rect 2012 56006 2014 56058
rect 2194 56006 2196 56058
rect 1950 56004 1956 56006
rect 2012 56004 2036 56006
rect 2092 56004 2116 56006
rect 2172 56004 2196 56006
rect 2252 56004 2258 56006
rect 1950 55995 2258 56004
rect 1950 54972 2258 54981
rect 1950 54970 1956 54972
rect 2012 54970 2036 54972
rect 2092 54970 2116 54972
rect 2172 54970 2196 54972
rect 2252 54970 2258 54972
rect 2012 54918 2014 54970
rect 2194 54918 2196 54970
rect 1950 54916 1956 54918
rect 2012 54916 2036 54918
rect 2092 54916 2116 54918
rect 2172 54916 2196 54918
rect 2252 54916 2258 54918
rect 1950 54907 2258 54916
rect 1950 53884 2258 53893
rect 1950 53882 1956 53884
rect 2012 53882 2036 53884
rect 2092 53882 2116 53884
rect 2172 53882 2196 53884
rect 2252 53882 2258 53884
rect 2012 53830 2014 53882
rect 2194 53830 2196 53882
rect 1950 53828 1956 53830
rect 2012 53828 2036 53830
rect 2092 53828 2116 53830
rect 2172 53828 2196 53830
rect 2252 53828 2258 53830
rect 1950 53819 2258 53828
rect 2516 53174 2544 61134
rect 2610 60956 2918 60965
rect 2610 60954 2616 60956
rect 2672 60954 2696 60956
rect 2752 60954 2776 60956
rect 2832 60954 2856 60956
rect 2912 60954 2918 60956
rect 2672 60902 2674 60954
rect 2854 60902 2856 60954
rect 2610 60900 2616 60902
rect 2672 60900 2696 60902
rect 2752 60900 2776 60902
rect 2832 60900 2856 60902
rect 2912 60900 2918 60902
rect 2610 60891 2918 60900
rect 2610 59868 2918 59877
rect 2610 59866 2616 59868
rect 2672 59866 2696 59868
rect 2752 59866 2776 59868
rect 2832 59866 2856 59868
rect 2912 59866 2918 59868
rect 2672 59814 2674 59866
rect 2854 59814 2856 59866
rect 2610 59812 2616 59814
rect 2672 59812 2696 59814
rect 2752 59812 2776 59814
rect 2832 59812 2856 59814
rect 2912 59812 2918 59814
rect 2610 59803 2918 59812
rect 2610 58780 2918 58789
rect 2610 58778 2616 58780
rect 2672 58778 2696 58780
rect 2752 58778 2776 58780
rect 2832 58778 2856 58780
rect 2912 58778 2918 58780
rect 2672 58726 2674 58778
rect 2854 58726 2856 58778
rect 2610 58724 2616 58726
rect 2672 58724 2696 58726
rect 2752 58724 2776 58726
rect 2832 58724 2856 58726
rect 2912 58724 2918 58726
rect 2610 58715 2918 58724
rect 2610 57692 2918 57701
rect 2610 57690 2616 57692
rect 2672 57690 2696 57692
rect 2752 57690 2776 57692
rect 2832 57690 2856 57692
rect 2912 57690 2918 57692
rect 2672 57638 2674 57690
rect 2854 57638 2856 57690
rect 2610 57636 2616 57638
rect 2672 57636 2696 57638
rect 2752 57636 2776 57638
rect 2832 57636 2856 57638
rect 2912 57636 2918 57638
rect 2610 57627 2918 57636
rect 2610 56604 2918 56613
rect 2610 56602 2616 56604
rect 2672 56602 2696 56604
rect 2752 56602 2776 56604
rect 2832 56602 2856 56604
rect 2912 56602 2918 56604
rect 2672 56550 2674 56602
rect 2854 56550 2856 56602
rect 2610 56548 2616 56550
rect 2672 56548 2696 56550
rect 2752 56548 2776 56550
rect 2832 56548 2856 56550
rect 2912 56548 2918 56550
rect 2610 56539 2918 56548
rect 2610 55516 2918 55525
rect 2610 55514 2616 55516
rect 2672 55514 2696 55516
rect 2752 55514 2776 55516
rect 2832 55514 2856 55516
rect 2912 55514 2918 55516
rect 2672 55462 2674 55514
rect 2854 55462 2856 55514
rect 2610 55460 2616 55462
rect 2672 55460 2696 55462
rect 2752 55460 2776 55462
rect 2832 55460 2856 55462
rect 2912 55460 2918 55462
rect 2610 55451 2918 55460
rect 2610 54428 2918 54437
rect 2610 54426 2616 54428
rect 2672 54426 2696 54428
rect 2752 54426 2776 54428
rect 2832 54426 2856 54428
rect 2912 54426 2918 54428
rect 2672 54374 2674 54426
rect 2854 54374 2856 54426
rect 2610 54372 2616 54374
rect 2672 54372 2696 54374
rect 2752 54372 2776 54374
rect 2832 54372 2856 54374
rect 2912 54372 2918 54374
rect 2610 54363 2918 54372
rect 2610 53340 2918 53349
rect 2610 53338 2616 53340
rect 2672 53338 2696 53340
rect 2752 53338 2776 53340
rect 2832 53338 2856 53340
rect 2912 53338 2918 53340
rect 2672 53286 2674 53338
rect 2854 53286 2856 53338
rect 2610 53284 2616 53286
rect 2672 53284 2696 53286
rect 2752 53284 2776 53286
rect 2832 53284 2856 53286
rect 2912 53284 2918 53286
rect 2610 53275 2918 53284
rect 2504 53168 2556 53174
rect 2504 53110 2556 53116
rect 1950 52796 2258 52805
rect 1950 52794 1956 52796
rect 2012 52794 2036 52796
rect 2092 52794 2116 52796
rect 2172 52794 2196 52796
rect 2252 52794 2258 52796
rect 2012 52742 2014 52794
rect 2194 52742 2196 52794
rect 1950 52740 1956 52742
rect 2012 52740 2036 52742
rect 2092 52740 2116 52742
rect 2172 52740 2196 52742
rect 2252 52740 2258 52742
rect 1950 52731 2258 52740
rect 2610 52252 2918 52261
rect 2610 52250 2616 52252
rect 2672 52250 2696 52252
rect 2752 52250 2776 52252
rect 2832 52250 2856 52252
rect 2912 52250 2918 52252
rect 2672 52198 2674 52250
rect 2854 52198 2856 52250
rect 2610 52196 2616 52198
rect 2672 52196 2696 52198
rect 2752 52196 2776 52198
rect 2832 52196 2856 52198
rect 2912 52196 2918 52198
rect 2610 52187 2918 52196
rect 1950 51708 2258 51717
rect 1950 51706 1956 51708
rect 2012 51706 2036 51708
rect 2092 51706 2116 51708
rect 2172 51706 2196 51708
rect 2252 51706 2258 51708
rect 2012 51654 2014 51706
rect 2194 51654 2196 51706
rect 1950 51652 1956 51654
rect 2012 51652 2036 51654
rect 2092 51652 2116 51654
rect 2172 51652 2196 51654
rect 2252 51652 2258 51654
rect 1950 51643 2258 51652
rect 2610 51164 2918 51173
rect 2610 51162 2616 51164
rect 2672 51162 2696 51164
rect 2752 51162 2776 51164
rect 2832 51162 2856 51164
rect 2912 51162 2918 51164
rect 2672 51110 2674 51162
rect 2854 51110 2856 51162
rect 2610 51108 2616 51110
rect 2672 51108 2696 51110
rect 2752 51108 2776 51110
rect 2832 51108 2856 51110
rect 2912 51108 2918 51110
rect 2610 51099 2918 51108
rect 1950 50620 2258 50629
rect 1950 50618 1956 50620
rect 2012 50618 2036 50620
rect 2092 50618 2116 50620
rect 2172 50618 2196 50620
rect 2252 50618 2258 50620
rect 2012 50566 2014 50618
rect 2194 50566 2196 50618
rect 1950 50564 1956 50566
rect 2012 50564 2036 50566
rect 2092 50564 2116 50566
rect 2172 50564 2196 50566
rect 2252 50564 2258 50566
rect 1950 50555 2258 50564
rect 2610 50076 2918 50085
rect 2610 50074 2616 50076
rect 2672 50074 2696 50076
rect 2752 50074 2776 50076
rect 2832 50074 2856 50076
rect 2912 50074 2918 50076
rect 2672 50022 2674 50074
rect 2854 50022 2856 50074
rect 2610 50020 2616 50022
rect 2672 50020 2696 50022
rect 2752 50020 2776 50022
rect 2832 50020 2856 50022
rect 2912 50020 2918 50022
rect 2610 50011 2918 50020
rect 1950 49532 2258 49541
rect 1950 49530 1956 49532
rect 2012 49530 2036 49532
rect 2092 49530 2116 49532
rect 2172 49530 2196 49532
rect 2252 49530 2258 49532
rect 2012 49478 2014 49530
rect 2194 49478 2196 49530
rect 1950 49476 1956 49478
rect 2012 49476 2036 49478
rect 2092 49476 2116 49478
rect 2172 49476 2196 49478
rect 2252 49476 2258 49478
rect 1950 49467 2258 49476
rect 2610 48988 2918 48997
rect 2610 48986 2616 48988
rect 2672 48986 2696 48988
rect 2752 48986 2776 48988
rect 2832 48986 2856 48988
rect 2912 48986 2918 48988
rect 2672 48934 2674 48986
rect 2854 48934 2856 48986
rect 2610 48932 2616 48934
rect 2672 48932 2696 48934
rect 2752 48932 2776 48934
rect 2832 48932 2856 48934
rect 2912 48932 2918 48934
rect 2610 48923 2918 48932
rect 1950 48444 2258 48453
rect 1950 48442 1956 48444
rect 2012 48442 2036 48444
rect 2092 48442 2116 48444
rect 2172 48442 2196 48444
rect 2252 48442 2258 48444
rect 2012 48390 2014 48442
rect 2194 48390 2196 48442
rect 1950 48388 1956 48390
rect 2012 48388 2036 48390
rect 2092 48388 2116 48390
rect 2172 48388 2196 48390
rect 2252 48388 2258 48390
rect 1950 48379 2258 48388
rect 2610 47900 2918 47909
rect 2610 47898 2616 47900
rect 2672 47898 2696 47900
rect 2752 47898 2776 47900
rect 2832 47898 2856 47900
rect 2912 47898 2918 47900
rect 2672 47846 2674 47898
rect 2854 47846 2856 47898
rect 2610 47844 2616 47846
rect 2672 47844 2696 47846
rect 2752 47844 2776 47846
rect 2832 47844 2856 47846
rect 2912 47844 2918 47846
rect 2610 47835 2918 47844
rect 2320 47592 2372 47598
rect 2320 47534 2372 47540
rect 1950 47356 2258 47365
rect 1950 47354 1956 47356
rect 2012 47354 2036 47356
rect 2092 47354 2116 47356
rect 2172 47354 2196 47356
rect 2252 47354 2258 47356
rect 2012 47302 2014 47354
rect 2194 47302 2196 47354
rect 1950 47300 1956 47302
rect 2012 47300 2036 47302
rect 2092 47300 2116 47302
rect 2172 47300 2196 47302
rect 2252 47300 2258 47302
rect 1950 47291 2258 47300
rect 1950 46268 2258 46277
rect 1950 46266 1956 46268
rect 2012 46266 2036 46268
rect 2092 46266 2116 46268
rect 2172 46266 2196 46268
rect 2252 46266 2258 46268
rect 2012 46214 2014 46266
rect 2194 46214 2196 46266
rect 1950 46212 1956 46214
rect 2012 46212 2036 46214
rect 2092 46212 2116 46214
rect 2172 46212 2196 46214
rect 2252 46212 2258 46214
rect 1950 46203 2258 46212
rect 1950 45180 2258 45189
rect 1950 45178 1956 45180
rect 2012 45178 2036 45180
rect 2092 45178 2116 45180
rect 2172 45178 2196 45180
rect 2252 45178 2258 45180
rect 2012 45126 2014 45178
rect 2194 45126 2196 45178
rect 1950 45124 1956 45126
rect 2012 45124 2036 45126
rect 2092 45124 2116 45126
rect 2172 45124 2196 45126
rect 2252 45124 2258 45126
rect 1950 45115 2258 45124
rect 1950 44092 2258 44101
rect 1950 44090 1956 44092
rect 2012 44090 2036 44092
rect 2092 44090 2116 44092
rect 2172 44090 2196 44092
rect 2252 44090 2258 44092
rect 2012 44038 2014 44090
rect 2194 44038 2196 44090
rect 1950 44036 1956 44038
rect 2012 44036 2036 44038
rect 2092 44036 2116 44038
rect 2172 44036 2196 44038
rect 2252 44036 2258 44038
rect 1950 44027 2258 44036
rect 1950 43004 2258 43013
rect 1950 43002 1956 43004
rect 2012 43002 2036 43004
rect 2092 43002 2116 43004
rect 2172 43002 2196 43004
rect 2252 43002 2258 43004
rect 2012 42950 2014 43002
rect 2194 42950 2196 43002
rect 1950 42948 1956 42950
rect 2012 42948 2036 42950
rect 2092 42948 2116 42950
rect 2172 42948 2196 42950
rect 2252 42948 2258 42950
rect 1950 42939 2258 42948
rect 1950 41916 2258 41925
rect 1950 41914 1956 41916
rect 2012 41914 2036 41916
rect 2092 41914 2116 41916
rect 2172 41914 2196 41916
rect 2252 41914 2258 41916
rect 2012 41862 2014 41914
rect 2194 41862 2196 41914
rect 1950 41860 1956 41862
rect 2012 41860 2036 41862
rect 2092 41860 2116 41862
rect 2172 41860 2196 41862
rect 2252 41860 2258 41862
rect 1950 41851 2258 41860
rect 1950 40828 2258 40837
rect 1950 40826 1956 40828
rect 2012 40826 2036 40828
rect 2092 40826 2116 40828
rect 2172 40826 2196 40828
rect 2252 40826 2258 40828
rect 2012 40774 2014 40826
rect 2194 40774 2196 40826
rect 1950 40772 1956 40774
rect 2012 40772 2036 40774
rect 2092 40772 2116 40774
rect 2172 40772 2196 40774
rect 2252 40772 2258 40774
rect 1950 40763 2258 40772
rect 1950 39740 2258 39749
rect 1950 39738 1956 39740
rect 2012 39738 2036 39740
rect 2092 39738 2116 39740
rect 2172 39738 2196 39740
rect 2252 39738 2258 39740
rect 2012 39686 2014 39738
rect 2194 39686 2196 39738
rect 1950 39684 1956 39686
rect 2012 39684 2036 39686
rect 2092 39684 2116 39686
rect 2172 39684 2196 39686
rect 2252 39684 2258 39686
rect 1950 39675 2258 39684
rect 1950 38652 2258 38661
rect 1950 38650 1956 38652
rect 2012 38650 2036 38652
rect 2092 38650 2116 38652
rect 2172 38650 2196 38652
rect 2252 38650 2258 38652
rect 2012 38598 2014 38650
rect 2194 38598 2196 38650
rect 1950 38596 1956 38598
rect 2012 38596 2036 38598
rect 2092 38596 2116 38598
rect 2172 38596 2196 38598
rect 2252 38596 2258 38598
rect 1950 38587 2258 38596
rect 1950 37564 2258 37573
rect 1950 37562 1956 37564
rect 2012 37562 2036 37564
rect 2092 37562 2116 37564
rect 2172 37562 2196 37564
rect 2252 37562 2258 37564
rect 2012 37510 2014 37562
rect 2194 37510 2196 37562
rect 1950 37508 1956 37510
rect 2012 37508 2036 37510
rect 2092 37508 2116 37510
rect 2172 37508 2196 37510
rect 2252 37508 2258 37510
rect 1950 37499 2258 37508
rect 1950 36476 2258 36485
rect 1950 36474 1956 36476
rect 2012 36474 2036 36476
rect 2092 36474 2116 36476
rect 2172 36474 2196 36476
rect 2252 36474 2258 36476
rect 2012 36422 2014 36474
rect 2194 36422 2196 36474
rect 1950 36420 1956 36422
rect 2012 36420 2036 36422
rect 2092 36420 2116 36422
rect 2172 36420 2196 36422
rect 2252 36420 2258 36422
rect 1950 36411 2258 36420
rect 1950 35388 2258 35397
rect 1950 35386 1956 35388
rect 2012 35386 2036 35388
rect 2092 35386 2116 35388
rect 2172 35386 2196 35388
rect 2252 35386 2258 35388
rect 2012 35334 2014 35386
rect 2194 35334 2196 35386
rect 1950 35332 1956 35334
rect 2012 35332 2036 35334
rect 2092 35332 2116 35334
rect 2172 35332 2196 35334
rect 2252 35332 2258 35334
rect 1950 35323 2258 35332
rect 1950 34300 2258 34309
rect 1950 34298 1956 34300
rect 2012 34298 2036 34300
rect 2092 34298 2116 34300
rect 2172 34298 2196 34300
rect 2252 34298 2258 34300
rect 2012 34246 2014 34298
rect 2194 34246 2196 34298
rect 1950 34244 1956 34246
rect 2012 34244 2036 34246
rect 2092 34244 2116 34246
rect 2172 34244 2196 34246
rect 2252 34244 2258 34246
rect 1950 34235 2258 34244
rect 1950 33212 2258 33221
rect 1950 33210 1956 33212
rect 2012 33210 2036 33212
rect 2092 33210 2116 33212
rect 2172 33210 2196 33212
rect 2252 33210 2258 33212
rect 2012 33158 2014 33210
rect 2194 33158 2196 33210
rect 1950 33156 1956 33158
rect 2012 33156 2036 33158
rect 2092 33156 2116 33158
rect 2172 33156 2196 33158
rect 2252 33156 2258 33158
rect 1950 33147 2258 33156
rect 1950 32124 2258 32133
rect 1950 32122 1956 32124
rect 2012 32122 2036 32124
rect 2092 32122 2116 32124
rect 2172 32122 2196 32124
rect 2252 32122 2258 32124
rect 2012 32070 2014 32122
rect 2194 32070 2196 32122
rect 1950 32068 1956 32070
rect 2012 32068 2036 32070
rect 2092 32068 2116 32070
rect 2172 32068 2196 32070
rect 2252 32068 2258 32070
rect 1950 32059 2258 32068
rect 1950 31036 2258 31045
rect 1950 31034 1956 31036
rect 2012 31034 2036 31036
rect 2092 31034 2116 31036
rect 2172 31034 2196 31036
rect 2252 31034 2258 31036
rect 2012 30982 2014 31034
rect 2194 30982 2196 31034
rect 1950 30980 1956 30982
rect 2012 30980 2036 30982
rect 2092 30980 2116 30982
rect 2172 30980 2196 30982
rect 2252 30980 2258 30982
rect 1950 30971 2258 30980
rect 1860 30728 1912 30734
rect 1860 30670 1912 30676
rect 1950 29948 2258 29957
rect 1950 29946 1956 29948
rect 2012 29946 2036 29948
rect 2092 29946 2116 29948
rect 2172 29946 2196 29948
rect 2252 29946 2258 29948
rect 2012 29894 2014 29946
rect 2194 29894 2196 29946
rect 1950 29892 1956 29894
rect 2012 29892 2036 29894
rect 2092 29892 2116 29894
rect 2172 29892 2196 29894
rect 2252 29892 2258 29894
rect 1950 29883 2258 29892
rect 1950 28860 2258 28869
rect 1950 28858 1956 28860
rect 2012 28858 2036 28860
rect 2092 28858 2116 28860
rect 2172 28858 2196 28860
rect 2252 28858 2258 28860
rect 2012 28806 2014 28858
rect 2194 28806 2196 28858
rect 1950 28804 1956 28806
rect 2012 28804 2036 28806
rect 2092 28804 2116 28806
rect 2172 28804 2196 28806
rect 2252 28804 2258 28806
rect 1950 28795 2258 28804
rect 1950 27772 2258 27781
rect 1950 27770 1956 27772
rect 2012 27770 2036 27772
rect 2092 27770 2116 27772
rect 2172 27770 2196 27772
rect 2252 27770 2258 27772
rect 2012 27718 2014 27770
rect 2194 27718 2196 27770
rect 1950 27716 1956 27718
rect 2012 27716 2036 27718
rect 2092 27716 2116 27718
rect 2172 27716 2196 27718
rect 2252 27716 2258 27718
rect 1950 27707 2258 27716
rect 1950 26684 2258 26693
rect 1950 26682 1956 26684
rect 2012 26682 2036 26684
rect 2092 26682 2116 26684
rect 2172 26682 2196 26684
rect 2252 26682 2258 26684
rect 2012 26630 2014 26682
rect 2194 26630 2196 26682
rect 1950 26628 1956 26630
rect 2012 26628 2036 26630
rect 2092 26628 2116 26630
rect 2172 26628 2196 26630
rect 2252 26628 2258 26630
rect 1950 26619 2258 26628
rect 1950 25596 2258 25605
rect 1950 25594 1956 25596
rect 2012 25594 2036 25596
rect 2092 25594 2116 25596
rect 2172 25594 2196 25596
rect 2252 25594 2258 25596
rect 2012 25542 2014 25594
rect 2194 25542 2196 25594
rect 1950 25540 1956 25542
rect 2012 25540 2036 25542
rect 2092 25540 2116 25542
rect 2172 25540 2196 25542
rect 2252 25540 2258 25542
rect 1950 25531 2258 25540
rect 1950 24508 2258 24517
rect 1950 24506 1956 24508
rect 2012 24506 2036 24508
rect 2092 24506 2116 24508
rect 2172 24506 2196 24508
rect 2252 24506 2258 24508
rect 2012 24454 2014 24506
rect 2194 24454 2196 24506
rect 1950 24452 1956 24454
rect 2012 24452 2036 24454
rect 2092 24452 2116 24454
rect 2172 24452 2196 24454
rect 2252 24452 2258 24454
rect 1950 24443 2258 24452
rect 1768 24268 1820 24274
rect 1768 24210 1820 24216
rect 1950 23420 2258 23429
rect 1950 23418 1956 23420
rect 2012 23418 2036 23420
rect 2092 23418 2116 23420
rect 2172 23418 2196 23420
rect 2252 23418 2258 23420
rect 2012 23366 2014 23418
rect 2194 23366 2196 23418
rect 1950 23364 1956 23366
rect 2012 23364 2036 23366
rect 2092 23364 2116 23366
rect 2172 23364 2196 23366
rect 2252 23364 2258 23366
rect 1950 23355 2258 23364
rect 1950 22332 2258 22341
rect 1950 22330 1956 22332
rect 2012 22330 2036 22332
rect 2092 22330 2116 22332
rect 2172 22330 2196 22332
rect 2252 22330 2258 22332
rect 2012 22278 2014 22330
rect 2194 22278 2196 22330
rect 1950 22276 1956 22278
rect 2012 22276 2036 22278
rect 2092 22276 2116 22278
rect 2172 22276 2196 22278
rect 2252 22276 2258 22278
rect 1950 22267 2258 22276
rect 1950 21244 2258 21253
rect 1950 21242 1956 21244
rect 2012 21242 2036 21244
rect 2092 21242 2116 21244
rect 2172 21242 2196 21244
rect 2252 21242 2258 21244
rect 2012 21190 2014 21242
rect 2194 21190 2196 21242
rect 1950 21188 1956 21190
rect 2012 21188 2036 21190
rect 2092 21188 2116 21190
rect 2172 21188 2196 21190
rect 2252 21188 2258 21190
rect 1950 21179 2258 21188
rect 1676 20596 1728 20602
rect 1676 20538 1728 20544
rect 1584 20528 1636 20534
rect 1584 20470 1636 20476
rect 1950 20156 2258 20165
rect 1950 20154 1956 20156
rect 2012 20154 2036 20156
rect 2092 20154 2116 20156
rect 2172 20154 2196 20156
rect 2252 20154 2258 20156
rect 2012 20102 2014 20154
rect 2194 20102 2196 20154
rect 1950 20100 1956 20102
rect 2012 20100 2036 20102
rect 2092 20100 2116 20102
rect 2172 20100 2196 20102
rect 2252 20100 2258 20102
rect 1950 20091 2258 20100
rect 1950 19068 2258 19077
rect 1950 19066 1956 19068
rect 2012 19066 2036 19068
rect 2092 19066 2116 19068
rect 2172 19066 2196 19068
rect 2252 19066 2258 19068
rect 2012 19014 2014 19066
rect 2194 19014 2196 19066
rect 1950 19012 1956 19014
rect 2012 19012 2036 19014
rect 2092 19012 2116 19014
rect 2172 19012 2196 19014
rect 2252 19012 2258 19014
rect 1950 19003 2258 19012
rect 1950 17980 2258 17989
rect 1950 17978 1956 17980
rect 2012 17978 2036 17980
rect 2092 17978 2116 17980
rect 2172 17978 2196 17980
rect 2252 17978 2258 17980
rect 2012 17926 2014 17978
rect 2194 17926 2196 17978
rect 1950 17924 1956 17926
rect 2012 17924 2036 17926
rect 2092 17924 2116 17926
rect 2172 17924 2196 17926
rect 2252 17924 2258 17926
rect 1950 17915 2258 17924
rect 1950 16892 2258 16901
rect 1950 16890 1956 16892
rect 2012 16890 2036 16892
rect 2092 16890 2116 16892
rect 2172 16890 2196 16892
rect 2252 16890 2258 16892
rect 2012 16838 2014 16890
rect 2194 16838 2196 16890
rect 1950 16836 1956 16838
rect 2012 16836 2036 16838
rect 2092 16836 2116 16838
rect 2172 16836 2196 16838
rect 2252 16836 2258 16838
rect 1950 16827 2258 16836
rect 2332 16114 2360 47534
rect 2610 46812 2918 46821
rect 2610 46810 2616 46812
rect 2672 46810 2696 46812
rect 2752 46810 2776 46812
rect 2832 46810 2856 46812
rect 2912 46810 2918 46812
rect 2672 46758 2674 46810
rect 2854 46758 2856 46810
rect 2610 46756 2616 46758
rect 2672 46756 2696 46758
rect 2752 46756 2776 46758
rect 2832 46756 2856 46758
rect 2912 46756 2918 46758
rect 2610 46747 2918 46756
rect 2610 45724 2918 45733
rect 2610 45722 2616 45724
rect 2672 45722 2696 45724
rect 2752 45722 2776 45724
rect 2832 45722 2856 45724
rect 2912 45722 2918 45724
rect 2672 45670 2674 45722
rect 2854 45670 2856 45722
rect 2610 45668 2616 45670
rect 2672 45668 2696 45670
rect 2752 45668 2776 45670
rect 2832 45668 2856 45670
rect 2912 45668 2918 45670
rect 2610 45659 2918 45668
rect 2610 44636 2918 44645
rect 2610 44634 2616 44636
rect 2672 44634 2696 44636
rect 2752 44634 2776 44636
rect 2832 44634 2856 44636
rect 2912 44634 2918 44636
rect 2672 44582 2674 44634
rect 2854 44582 2856 44634
rect 2610 44580 2616 44582
rect 2672 44580 2696 44582
rect 2752 44580 2776 44582
rect 2832 44580 2856 44582
rect 2912 44580 2918 44582
rect 2610 44571 2918 44580
rect 2610 43548 2918 43557
rect 2610 43546 2616 43548
rect 2672 43546 2696 43548
rect 2752 43546 2776 43548
rect 2832 43546 2856 43548
rect 2912 43546 2918 43548
rect 2672 43494 2674 43546
rect 2854 43494 2856 43546
rect 2610 43492 2616 43494
rect 2672 43492 2696 43494
rect 2752 43492 2776 43494
rect 2832 43492 2856 43494
rect 2912 43492 2918 43494
rect 2610 43483 2918 43492
rect 2610 42460 2918 42469
rect 2610 42458 2616 42460
rect 2672 42458 2696 42460
rect 2752 42458 2776 42460
rect 2832 42458 2856 42460
rect 2912 42458 2918 42460
rect 2672 42406 2674 42458
rect 2854 42406 2856 42458
rect 2610 42404 2616 42406
rect 2672 42404 2696 42406
rect 2752 42404 2776 42406
rect 2832 42404 2856 42406
rect 2912 42404 2918 42406
rect 2610 42395 2918 42404
rect 2976 41414 3004 65554
rect 4436 62144 4488 62150
rect 4436 62086 4488 62092
rect 3700 61124 3752 61130
rect 3700 61066 3752 61072
rect 3056 50448 3108 50454
rect 3056 50390 3108 50396
rect 3068 42770 3096 50390
rect 3424 45484 3476 45490
rect 3424 45426 3476 45432
rect 3056 42764 3108 42770
rect 3056 42706 3108 42712
rect 2976 41386 3188 41414
rect 2610 41372 2918 41381
rect 2610 41370 2616 41372
rect 2672 41370 2696 41372
rect 2752 41370 2776 41372
rect 2832 41370 2856 41372
rect 2912 41370 2918 41372
rect 2672 41318 2674 41370
rect 2854 41318 2856 41370
rect 2610 41316 2616 41318
rect 2672 41316 2696 41318
rect 2752 41316 2776 41318
rect 2832 41316 2856 41318
rect 2912 41316 2918 41318
rect 2610 41307 2918 41316
rect 2964 40520 3016 40526
rect 2964 40462 3016 40468
rect 2610 40284 2918 40293
rect 2610 40282 2616 40284
rect 2672 40282 2696 40284
rect 2752 40282 2776 40284
rect 2832 40282 2856 40284
rect 2912 40282 2918 40284
rect 2672 40230 2674 40282
rect 2854 40230 2856 40282
rect 2610 40228 2616 40230
rect 2672 40228 2696 40230
rect 2752 40228 2776 40230
rect 2832 40228 2856 40230
rect 2912 40228 2918 40230
rect 2610 40219 2918 40228
rect 2504 39840 2556 39846
rect 2504 39782 2556 39788
rect 2516 30802 2544 39782
rect 2610 39196 2918 39205
rect 2610 39194 2616 39196
rect 2672 39194 2696 39196
rect 2752 39194 2776 39196
rect 2832 39194 2856 39196
rect 2912 39194 2918 39196
rect 2672 39142 2674 39194
rect 2854 39142 2856 39194
rect 2610 39140 2616 39142
rect 2672 39140 2696 39142
rect 2752 39140 2776 39142
rect 2832 39140 2856 39142
rect 2912 39140 2918 39142
rect 2610 39131 2918 39140
rect 2610 38108 2918 38117
rect 2610 38106 2616 38108
rect 2672 38106 2696 38108
rect 2752 38106 2776 38108
rect 2832 38106 2856 38108
rect 2912 38106 2918 38108
rect 2672 38054 2674 38106
rect 2854 38054 2856 38106
rect 2610 38052 2616 38054
rect 2672 38052 2696 38054
rect 2752 38052 2776 38054
rect 2832 38052 2856 38054
rect 2912 38052 2918 38054
rect 2610 38043 2918 38052
rect 2610 37020 2918 37029
rect 2610 37018 2616 37020
rect 2672 37018 2696 37020
rect 2752 37018 2776 37020
rect 2832 37018 2856 37020
rect 2912 37018 2918 37020
rect 2672 36966 2674 37018
rect 2854 36966 2856 37018
rect 2610 36964 2616 36966
rect 2672 36964 2696 36966
rect 2752 36964 2776 36966
rect 2832 36964 2856 36966
rect 2912 36964 2918 36966
rect 2610 36955 2918 36964
rect 2610 35932 2918 35941
rect 2610 35930 2616 35932
rect 2672 35930 2696 35932
rect 2752 35930 2776 35932
rect 2832 35930 2856 35932
rect 2912 35930 2918 35932
rect 2672 35878 2674 35930
rect 2854 35878 2856 35930
rect 2610 35876 2616 35878
rect 2672 35876 2696 35878
rect 2752 35876 2776 35878
rect 2832 35876 2856 35878
rect 2912 35876 2918 35878
rect 2610 35867 2918 35876
rect 2610 34844 2918 34853
rect 2610 34842 2616 34844
rect 2672 34842 2696 34844
rect 2752 34842 2776 34844
rect 2832 34842 2856 34844
rect 2912 34842 2918 34844
rect 2672 34790 2674 34842
rect 2854 34790 2856 34842
rect 2610 34788 2616 34790
rect 2672 34788 2696 34790
rect 2752 34788 2776 34790
rect 2832 34788 2856 34790
rect 2912 34788 2918 34790
rect 2610 34779 2918 34788
rect 2976 34134 3004 40462
rect 3056 40452 3108 40458
rect 3056 40394 3108 40400
rect 2964 34128 3016 34134
rect 2964 34070 3016 34076
rect 2610 33756 2918 33765
rect 2610 33754 2616 33756
rect 2672 33754 2696 33756
rect 2752 33754 2776 33756
rect 2832 33754 2856 33756
rect 2912 33754 2918 33756
rect 2672 33702 2674 33754
rect 2854 33702 2856 33754
rect 2610 33700 2616 33702
rect 2672 33700 2696 33702
rect 2752 33700 2776 33702
rect 2832 33700 2856 33702
rect 2912 33700 2918 33702
rect 2610 33691 2918 33700
rect 2610 32668 2918 32677
rect 2610 32666 2616 32668
rect 2672 32666 2696 32668
rect 2752 32666 2776 32668
rect 2832 32666 2856 32668
rect 2912 32666 2918 32668
rect 2672 32614 2674 32666
rect 2854 32614 2856 32666
rect 2610 32612 2616 32614
rect 2672 32612 2696 32614
rect 2752 32612 2776 32614
rect 2832 32612 2856 32614
rect 2912 32612 2918 32614
rect 2610 32603 2918 32612
rect 3068 31754 3096 40394
rect 3160 33046 3188 41386
rect 3436 41070 3464 45426
rect 3424 41064 3476 41070
rect 3424 41006 3476 41012
rect 3516 40520 3568 40526
rect 3516 40462 3568 40468
rect 3528 33930 3556 40462
rect 3516 33924 3568 33930
rect 3516 33866 3568 33872
rect 3148 33040 3200 33046
rect 3148 32982 3200 32988
rect 3068 31726 3188 31754
rect 2610 31580 2918 31589
rect 2610 31578 2616 31580
rect 2672 31578 2696 31580
rect 2752 31578 2776 31580
rect 2832 31578 2856 31580
rect 2912 31578 2918 31580
rect 2672 31526 2674 31578
rect 2854 31526 2856 31578
rect 2610 31524 2616 31526
rect 2672 31524 2696 31526
rect 2752 31524 2776 31526
rect 2832 31524 2856 31526
rect 2912 31524 2918 31526
rect 2610 31515 2918 31524
rect 2504 30796 2556 30802
rect 2504 30738 2556 30744
rect 2610 30492 2918 30501
rect 2610 30490 2616 30492
rect 2672 30490 2696 30492
rect 2752 30490 2776 30492
rect 2832 30490 2856 30492
rect 2912 30490 2918 30492
rect 2672 30438 2674 30490
rect 2854 30438 2856 30490
rect 2610 30436 2616 30438
rect 2672 30436 2696 30438
rect 2752 30436 2776 30438
rect 2832 30436 2856 30438
rect 2912 30436 2918 30438
rect 2610 30427 2918 30436
rect 2610 29404 2918 29413
rect 2610 29402 2616 29404
rect 2672 29402 2696 29404
rect 2752 29402 2776 29404
rect 2832 29402 2856 29404
rect 2912 29402 2918 29404
rect 2672 29350 2674 29402
rect 2854 29350 2856 29402
rect 2610 29348 2616 29350
rect 2672 29348 2696 29350
rect 2752 29348 2776 29350
rect 2832 29348 2856 29350
rect 2912 29348 2918 29350
rect 2610 29339 2918 29348
rect 2610 28316 2918 28325
rect 2610 28314 2616 28316
rect 2672 28314 2696 28316
rect 2752 28314 2776 28316
rect 2832 28314 2856 28316
rect 2912 28314 2918 28316
rect 2672 28262 2674 28314
rect 2854 28262 2856 28314
rect 2610 28260 2616 28262
rect 2672 28260 2696 28262
rect 2752 28260 2776 28262
rect 2832 28260 2856 28262
rect 2912 28260 2918 28262
rect 2610 28251 2918 28260
rect 2610 27228 2918 27237
rect 2610 27226 2616 27228
rect 2672 27226 2696 27228
rect 2752 27226 2776 27228
rect 2832 27226 2856 27228
rect 2912 27226 2918 27228
rect 2672 27174 2674 27226
rect 2854 27174 2856 27226
rect 2610 27172 2616 27174
rect 2672 27172 2696 27174
rect 2752 27172 2776 27174
rect 2832 27172 2856 27174
rect 2912 27172 2918 27174
rect 2610 27163 2918 27172
rect 2610 26140 2918 26149
rect 2610 26138 2616 26140
rect 2672 26138 2696 26140
rect 2752 26138 2776 26140
rect 2832 26138 2856 26140
rect 2912 26138 2918 26140
rect 2672 26086 2674 26138
rect 2854 26086 2856 26138
rect 2610 26084 2616 26086
rect 2672 26084 2696 26086
rect 2752 26084 2776 26086
rect 2832 26084 2856 26086
rect 2912 26084 2918 26086
rect 2610 26075 2918 26084
rect 2412 25968 2464 25974
rect 2412 25910 2464 25916
rect 2320 16108 2372 16114
rect 2320 16050 2372 16056
rect 2320 15904 2372 15910
rect 2320 15846 2372 15852
rect 1950 15804 2258 15813
rect 1950 15802 1956 15804
rect 2012 15802 2036 15804
rect 2092 15802 2116 15804
rect 2172 15802 2196 15804
rect 2252 15802 2258 15804
rect 2012 15750 2014 15802
rect 2194 15750 2196 15802
rect 1950 15748 1956 15750
rect 2012 15748 2036 15750
rect 2092 15748 2116 15750
rect 2172 15748 2196 15750
rect 2252 15748 2258 15750
rect 1950 15739 2258 15748
rect 1950 14716 2258 14725
rect 1950 14714 1956 14716
rect 2012 14714 2036 14716
rect 2092 14714 2116 14716
rect 2172 14714 2196 14716
rect 2252 14714 2258 14716
rect 2012 14662 2014 14714
rect 2194 14662 2196 14714
rect 1950 14660 1956 14662
rect 2012 14660 2036 14662
rect 2092 14660 2116 14662
rect 2172 14660 2196 14662
rect 2252 14660 2258 14662
rect 1950 14651 2258 14660
rect 1950 13628 2258 13637
rect 1950 13626 1956 13628
rect 2012 13626 2036 13628
rect 2092 13626 2116 13628
rect 2172 13626 2196 13628
rect 2252 13626 2258 13628
rect 2012 13574 2014 13626
rect 2194 13574 2196 13626
rect 1950 13572 1956 13574
rect 2012 13572 2036 13574
rect 2092 13572 2116 13574
rect 2172 13572 2196 13574
rect 2252 13572 2258 13574
rect 1950 13563 2258 13572
rect 1950 12540 2258 12549
rect 1950 12538 1956 12540
rect 2012 12538 2036 12540
rect 2092 12538 2116 12540
rect 2172 12538 2196 12540
rect 2252 12538 2258 12540
rect 2012 12486 2014 12538
rect 2194 12486 2196 12538
rect 1950 12484 1956 12486
rect 2012 12484 2036 12486
rect 2092 12484 2116 12486
rect 2172 12484 2196 12486
rect 2252 12484 2258 12486
rect 1950 12475 2258 12484
rect 1950 11452 2258 11461
rect 1950 11450 1956 11452
rect 2012 11450 2036 11452
rect 2092 11450 2116 11452
rect 2172 11450 2196 11452
rect 2252 11450 2258 11452
rect 2012 11398 2014 11450
rect 2194 11398 2196 11450
rect 1950 11396 1956 11398
rect 2012 11396 2036 11398
rect 2092 11396 2116 11398
rect 2172 11396 2196 11398
rect 2252 11396 2258 11398
rect 1950 11387 2258 11396
rect 1858 11112 1914 11121
rect 1858 11047 1914 11056
rect 1872 9042 1900 11047
rect 1950 10364 2258 10373
rect 1950 10362 1956 10364
rect 2012 10362 2036 10364
rect 2092 10362 2116 10364
rect 2172 10362 2196 10364
rect 2252 10362 2258 10364
rect 2012 10310 2014 10362
rect 2194 10310 2196 10362
rect 1950 10308 1956 10310
rect 2012 10308 2036 10310
rect 2092 10308 2116 10310
rect 2172 10308 2196 10310
rect 2252 10308 2258 10310
rect 1950 10299 2258 10308
rect 1950 9276 2258 9285
rect 1950 9274 1956 9276
rect 2012 9274 2036 9276
rect 2092 9274 2116 9276
rect 2172 9274 2196 9276
rect 2252 9274 2258 9276
rect 2012 9222 2014 9274
rect 2194 9222 2196 9274
rect 1950 9220 1956 9222
rect 2012 9220 2036 9222
rect 2092 9220 2116 9222
rect 2172 9220 2196 9222
rect 2252 9220 2258 9222
rect 1950 9211 2258 9220
rect 1860 9036 1912 9042
rect 1860 8978 1912 8984
rect 1950 8188 2258 8197
rect 1950 8186 1956 8188
rect 2012 8186 2036 8188
rect 2092 8186 2116 8188
rect 2172 8186 2196 8188
rect 2252 8186 2258 8188
rect 2012 8134 2014 8186
rect 2194 8134 2196 8186
rect 1950 8132 1956 8134
rect 2012 8132 2036 8134
rect 2092 8132 2116 8134
rect 2172 8132 2196 8134
rect 2252 8132 2258 8134
rect 1950 8123 2258 8132
rect 1950 7100 2258 7109
rect 1950 7098 1956 7100
rect 2012 7098 2036 7100
rect 2092 7098 2116 7100
rect 2172 7098 2196 7100
rect 2252 7098 2258 7100
rect 2012 7046 2014 7098
rect 2194 7046 2196 7098
rect 1950 7044 1956 7046
rect 2012 7044 2036 7046
rect 2092 7044 2116 7046
rect 2172 7044 2196 7046
rect 2252 7044 2258 7046
rect 1950 7035 2258 7044
rect 1412 6886 1532 6914
rect 1412 6390 1440 6886
rect 1400 6384 1452 6390
rect 1400 6326 1452 6332
rect 1950 6012 2258 6021
rect 1950 6010 1956 6012
rect 2012 6010 2036 6012
rect 2092 6010 2116 6012
rect 2172 6010 2196 6012
rect 2252 6010 2258 6012
rect 2012 5958 2014 6010
rect 2194 5958 2196 6010
rect 1950 5956 1956 5958
rect 2012 5956 2036 5958
rect 2092 5956 2116 5958
rect 2172 5956 2196 5958
rect 2252 5956 2258 5958
rect 1950 5947 2258 5956
rect 1950 4924 2258 4933
rect 1950 4922 1956 4924
rect 2012 4922 2036 4924
rect 2092 4922 2116 4924
rect 2172 4922 2196 4924
rect 2252 4922 2258 4924
rect 2012 4870 2014 4922
rect 2194 4870 2196 4922
rect 1950 4868 1956 4870
rect 2012 4868 2036 4870
rect 2092 4868 2116 4870
rect 2172 4868 2196 4870
rect 2252 4868 2258 4870
rect 1950 4859 2258 4868
rect 848 4616 900 4622
rect 846 4584 848 4593
rect 900 4584 902 4593
rect 846 4519 902 4528
rect 1950 3836 2258 3845
rect 1950 3834 1956 3836
rect 2012 3834 2036 3836
rect 2092 3834 2116 3836
rect 2172 3834 2196 3836
rect 2252 3834 2258 3836
rect 2012 3782 2014 3834
rect 2194 3782 2196 3834
rect 1950 3780 1956 3782
rect 2012 3780 2036 3782
rect 2092 3780 2116 3782
rect 2172 3780 2196 3782
rect 2252 3780 2258 3782
rect 1950 3771 2258 3780
rect 1950 2748 2258 2757
rect 1950 2746 1956 2748
rect 2012 2746 2036 2748
rect 2092 2746 2116 2748
rect 2172 2746 2196 2748
rect 2252 2746 2258 2748
rect 2012 2694 2014 2746
rect 2194 2694 2196 2746
rect 1950 2692 1956 2694
rect 2012 2692 2036 2694
rect 2092 2692 2116 2694
rect 2172 2692 2196 2694
rect 2252 2692 2258 2694
rect 1950 2683 2258 2692
rect 2332 2310 2360 15846
rect 2424 11150 2452 25910
rect 2610 25052 2918 25061
rect 2610 25050 2616 25052
rect 2672 25050 2696 25052
rect 2752 25050 2776 25052
rect 2832 25050 2856 25052
rect 2912 25050 2918 25052
rect 2672 24998 2674 25050
rect 2854 24998 2856 25050
rect 2610 24996 2616 24998
rect 2672 24996 2696 24998
rect 2752 24996 2776 24998
rect 2832 24996 2856 24998
rect 2912 24996 2918 24998
rect 2610 24987 2918 24996
rect 2610 23964 2918 23973
rect 2610 23962 2616 23964
rect 2672 23962 2696 23964
rect 2752 23962 2776 23964
rect 2832 23962 2856 23964
rect 2912 23962 2918 23964
rect 2672 23910 2674 23962
rect 2854 23910 2856 23962
rect 2610 23908 2616 23910
rect 2672 23908 2696 23910
rect 2752 23908 2776 23910
rect 2832 23908 2856 23910
rect 2912 23908 2918 23910
rect 2610 23899 2918 23908
rect 2610 22876 2918 22885
rect 2610 22874 2616 22876
rect 2672 22874 2696 22876
rect 2752 22874 2776 22876
rect 2832 22874 2856 22876
rect 2912 22874 2918 22876
rect 2672 22822 2674 22874
rect 2854 22822 2856 22874
rect 2610 22820 2616 22822
rect 2672 22820 2696 22822
rect 2752 22820 2776 22822
rect 2832 22820 2856 22822
rect 2912 22820 2918 22822
rect 2610 22811 2918 22820
rect 2610 21788 2918 21797
rect 2610 21786 2616 21788
rect 2672 21786 2696 21788
rect 2752 21786 2776 21788
rect 2832 21786 2856 21788
rect 2912 21786 2918 21788
rect 2672 21734 2674 21786
rect 2854 21734 2856 21786
rect 2610 21732 2616 21734
rect 2672 21732 2696 21734
rect 2752 21732 2776 21734
rect 2832 21732 2856 21734
rect 2912 21732 2918 21734
rect 2610 21723 2918 21732
rect 2610 20700 2918 20709
rect 2610 20698 2616 20700
rect 2672 20698 2696 20700
rect 2752 20698 2776 20700
rect 2832 20698 2856 20700
rect 2912 20698 2918 20700
rect 2672 20646 2674 20698
rect 2854 20646 2856 20698
rect 2610 20644 2616 20646
rect 2672 20644 2696 20646
rect 2752 20644 2776 20646
rect 2832 20644 2856 20646
rect 2912 20644 2918 20646
rect 2610 20635 2918 20644
rect 2610 19612 2918 19621
rect 2610 19610 2616 19612
rect 2672 19610 2696 19612
rect 2752 19610 2776 19612
rect 2832 19610 2856 19612
rect 2912 19610 2918 19612
rect 2672 19558 2674 19610
rect 2854 19558 2856 19610
rect 2610 19556 2616 19558
rect 2672 19556 2696 19558
rect 2752 19556 2776 19558
rect 2832 19556 2856 19558
rect 2912 19556 2918 19558
rect 2610 19547 2918 19556
rect 2610 18524 2918 18533
rect 2610 18522 2616 18524
rect 2672 18522 2696 18524
rect 2752 18522 2776 18524
rect 2832 18522 2856 18524
rect 2912 18522 2918 18524
rect 2672 18470 2674 18522
rect 2854 18470 2856 18522
rect 2610 18468 2616 18470
rect 2672 18468 2696 18470
rect 2752 18468 2776 18470
rect 2832 18468 2856 18470
rect 2912 18468 2918 18470
rect 2610 18459 2918 18468
rect 2610 17436 2918 17445
rect 2610 17434 2616 17436
rect 2672 17434 2696 17436
rect 2752 17434 2776 17436
rect 2832 17434 2856 17436
rect 2912 17434 2918 17436
rect 2672 17382 2674 17434
rect 2854 17382 2856 17434
rect 2610 17380 2616 17382
rect 2672 17380 2696 17382
rect 2752 17380 2776 17382
rect 2832 17380 2856 17382
rect 2912 17380 2918 17382
rect 2610 17371 2918 17380
rect 3056 17332 3108 17338
rect 3056 17274 3108 17280
rect 2610 16348 2918 16357
rect 2610 16346 2616 16348
rect 2672 16346 2696 16348
rect 2752 16346 2776 16348
rect 2832 16346 2856 16348
rect 2912 16346 2918 16348
rect 2672 16294 2674 16346
rect 2854 16294 2856 16346
rect 2610 16292 2616 16294
rect 2672 16292 2696 16294
rect 2752 16292 2776 16294
rect 2832 16292 2856 16294
rect 2912 16292 2918 16294
rect 2610 16283 2918 16292
rect 2610 15260 2918 15269
rect 2610 15258 2616 15260
rect 2672 15258 2696 15260
rect 2752 15258 2776 15260
rect 2832 15258 2856 15260
rect 2912 15258 2918 15260
rect 2672 15206 2674 15258
rect 2854 15206 2856 15258
rect 2610 15204 2616 15206
rect 2672 15204 2696 15206
rect 2752 15204 2776 15206
rect 2832 15204 2856 15206
rect 2912 15204 2918 15206
rect 2610 15195 2918 15204
rect 2610 14172 2918 14181
rect 2610 14170 2616 14172
rect 2672 14170 2696 14172
rect 2752 14170 2776 14172
rect 2832 14170 2856 14172
rect 2912 14170 2918 14172
rect 2672 14118 2674 14170
rect 2854 14118 2856 14170
rect 2610 14116 2616 14118
rect 2672 14116 2696 14118
rect 2752 14116 2776 14118
rect 2832 14116 2856 14118
rect 2912 14116 2918 14118
rect 2610 14107 2918 14116
rect 2610 13084 2918 13093
rect 2610 13082 2616 13084
rect 2672 13082 2696 13084
rect 2752 13082 2776 13084
rect 2832 13082 2856 13084
rect 2912 13082 2918 13084
rect 2672 13030 2674 13082
rect 2854 13030 2856 13082
rect 2610 13028 2616 13030
rect 2672 13028 2696 13030
rect 2752 13028 2776 13030
rect 2832 13028 2856 13030
rect 2912 13028 2918 13030
rect 2610 13019 2918 13028
rect 2610 11996 2918 12005
rect 2610 11994 2616 11996
rect 2672 11994 2696 11996
rect 2752 11994 2776 11996
rect 2832 11994 2856 11996
rect 2912 11994 2918 11996
rect 2672 11942 2674 11994
rect 2854 11942 2856 11994
rect 2610 11940 2616 11942
rect 2672 11940 2696 11942
rect 2752 11940 2776 11942
rect 2832 11940 2856 11942
rect 2912 11940 2918 11942
rect 2610 11931 2918 11940
rect 2412 11144 2464 11150
rect 2412 11086 2464 11092
rect 2610 10908 2918 10917
rect 2610 10906 2616 10908
rect 2672 10906 2696 10908
rect 2752 10906 2776 10908
rect 2832 10906 2856 10908
rect 2912 10906 2918 10908
rect 2672 10854 2674 10906
rect 2854 10854 2856 10906
rect 2610 10852 2616 10854
rect 2672 10852 2696 10854
rect 2752 10852 2776 10854
rect 2832 10852 2856 10854
rect 2912 10852 2918 10854
rect 2610 10843 2918 10852
rect 3068 10674 3096 17274
rect 3160 11762 3188 31726
rect 3516 30728 3568 30734
rect 3516 30670 3568 30676
rect 3424 24812 3476 24818
rect 3424 24754 3476 24760
rect 3436 20942 3464 24754
rect 3528 20942 3556 30670
rect 3608 23316 3660 23322
rect 3608 23258 3660 23264
rect 3620 22438 3648 23258
rect 3608 22432 3660 22438
rect 3608 22374 3660 22380
rect 3424 20936 3476 20942
rect 3424 20878 3476 20884
rect 3516 20936 3568 20942
rect 3516 20878 3568 20884
rect 3528 16250 3556 20878
rect 3516 16244 3568 16250
rect 3516 16186 3568 16192
rect 3148 11756 3200 11762
rect 3148 11698 3200 11704
rect 3056 10668 3108 10674
rect 3056 10610 3108 10616
rect 2610 9820 2918 9829
rect 2610 9818 2616 9820
rect 2672 9818 2696 9820
rect 2752 9818 2776 9820
rect 2832 9818 2856 9820
rect 2912 9818 2918 9820
rect 2672 9766 2674 9818
rect 2854 9766 2856 9818
rect 2610 9764 2616 9766
rect 2672 9764 2696 9766
rect 2752 9764 2776 9766
rect 2832 9764 2856 9766
rect 2912 9764 2918 9766
rect 2610 9755 2918 9764
rect 2504 9512 2556 9518
rect 2504 9454 2556 9460
rect 2516 8974 2544 9454
rect 3620 9110 3648 22374
rect 3608 9104 3660 9110
rect 3608 9046 3660 9052
rect 2504 8968 2556 8974
rect 2504 8910 2556 8916
rect 2610 8732 2918 8741
rect 2610 8730 2616 8732
rect 2672 8730 2696 8732
rect 2752 8730 2776 8732
rect 2832 8730 2856 8732
rect 2912 8730 2918 8732
rect 2672 8678 2674 8730
rect 2854 8678 2856 8730
rect 2610 8676 2616 8678
rect 2672 8676 2696 8678
rect 2752 8676 2776 8678
rect 2832 8676 2856 8678
rect 2912 8676 2918 8678
rect 2610 8667 2918 8676
rect 2610 7644 2918 7653
rect 2610 7642 2616 7644
rect 2672 7642 2696 7644
rect 2752 7642 2776 7644
rect 2832 7642 2856 7644
rect 2912 7642 2918 7644
rect 2672 7590 2674 7642
rect 2854 7590 2856 7642
rect 2610 7588 2616 7590
rect 2672 7588 2696 7590
rect 2752 7588 2776 7590
rect 2832 7588 2856 7590
rect 2912 7588 2918 7590
rect 2610 7579 2918 7588
rect 2610 6556 2918 6565
rect 2610 6554 2616 6556
rect 2672 6554 2696 6556
rect 2752 6554 2776 6556
rect 2832 6554 2856 6556
rect 2912 6554 2918 6556
rect 2672 6502 2674 6554
rect 2854 6502 2856 6554
rect 2610 6500 2616 6502
rect 2672 6500 2696 6502
rect 2752 6500 2776 6502
rect 2832 6500 2856 6502
rect 2912 6500 2918 6502
rect 2610 6491 2918 6500
rect 2610 5468 2918 5477
rect 2610 5466 2616 5468
rect 2672 5466 2696 5468
rect 2752 5466 2776 5468
rect 2832 5466 2856 5468
rect 2912 5466 2918 5468
rect 2672 5414 2674 5466
rect 2854 5414 2856 5466
rect 2610 5412 2616 5414
rect 2672 5412 2696 5414
rect 2752 5412 2776 5414
rect 2832 5412 2856 5414
rect 2912 5412 2918 5414
rect 2610 5403 2918 5412
rect 3712 5370 3740 61066
rect 3884 61056 3936 61062
rect 3884 60998 3936 61004
rect 3792 55888 3844 55894
rect 3792 55830 3844 55836
rect 3804 35290 3832 55830
rect 3896 49978 3924 60998
rect 4344 59016 4396 59022
rect 4344 58958 4396 58964
rect 4252 54528 4304 54534
rect 4252 54470 4304 54476
rect 3884 49972 3936 49978
rect 3884 49914 3936 49920
rect 3976 47660 4028 47666
rect 3976 47602 4028 47608
rect 3884 41064 3936 41070
rect 3884 41006 3936 41012
rect 3896 35714 3924 41006
rect 3988 35834 4016 47602
rect 4264 39574 4292 54470
rect 4252 39568 4304 39574
rect 4252 39510 4304 39516
rect 4158 36680 4214 36689
rect 4158 36615 4214 36624
rect 3976 35828 4028 35834
rect 3976 35770 4028 35776
rect 3896 35686 4016 35714
rect 4172 35698 4200 36615
rect 3988 35562 4016 35686
rect 4160 35692 4212 35698
rect 4160 35634 4212 35640
rect 3976 35556 4028 35562
rect 3976 35498 4028 35504
rect 3792 35284 3844 35290
rect 3792 35226 3844 35232
rect 3988 23322 4016 35498
rect 4068 34944 4120 34950
rect 4068 34886 4120 34892
rect 4080 26858 4108 34886
rect 4068 26852 4120 26858
rect 4068 26794 4120 26800
rect 3976 23316 4028 23322
rect 3976 23258 4028 23264
rect 4356 19854 4384 58958
rect 4448 53582 4476 62086
rect 4436 53576 4488 53582
rect 4436 53518 4488 53524
rect 4344 19848 4396 19854
rect 4344 19790 4396 19796
rect 4540 17542 4568 66098
rect 4988 66020 5040 66026
rect 4988 65962 5040 65968
rect 4896 62756 4948 62762
rect 4896 62698 4948 62704
rect 4712 61124 4764 61130
rect 4712 61066 4764 61072
rect 4620 58948 4672 58954
rect 4620 58890 4672 58896
rect 4632 19990 4660 58890
rect 4724 54534 4752 61066
rect 4804 61056 4856 61062
rect 4804 60998 4856 61004
rect 4816 60790 4844 60998
rect 4804 60784 4856 60790
rect 4804 60726 4856 60732
rect 4908 55214 4936 62698
rect 4816 55186 4936 55214
rect 4712 54528 4764 54534
rect 4712 54470 4764 54476
rect 4712 29096 4764 29102
rect 4712 29038 4764 29044
rect 4724 26382 4752 29038
rect 4712 26376 4764 26382
rect 4712 26318 4764 26324
rect 4816 20806 4844 55186
rect 4896 52012 4948 52018
rect 4896 51954 4948 51960
rect 4908 44198 4936 51954
rect 5000 51814 5028 65962
rect 6368 65612 6420 65618
rect 6368 65554 6420 65560
rect 5540 61192 5592 61198
rect 5540 61134 5592 61140
rect 5552 60654 5580 61134
rect 5540 60648 5592 60654
rect 5540 60590 5592 60596
rect 5540 60512 5592 60518
rect 5540 60454 5592 60460
rect 5080 56840 5132 56846
rect 5080 56782 5132 56788
rect 4988 51808 5040 51814
rect 4988 51750 5040 51756
rect 5092 45554 5120 56782
rect 5552 54602 5580 60454
rect 6000 60104 6052 60110
rect 6000 60046 6052 60052
rect 5540 54596 5592 54602
rect 5540 54538 5592 54544
rect 5908 54596 5960 54602
rect 5908 54538 5960 54544
rect 5000 45526 5120 45554
rect 4896 44192 4948 44198
rect 4896 44134 4948 44140
rect 4896 33108 4948 33114
rect 4896 33050 4948 33056
rect 4804 20800 4856 20806
rect 4804 20742 4856 20748
rect 4620 19984 4672 19990
rect 4620 19926 4672 19932
rect 4528 17536 4580 17542
rect 4528 17478 4580 17484
rect 4632 16574 4660 19926
rect 4632 16546 4844 16574
rect 3790 11656 3846 11665
rect 3790 11591 3846 11600
rect 3700 5364 3752 5370
rect 3700 5306 3752 5312
rect 3712 4690 3740 5306
rect 3804 4690 3832 11591
rect 4344 5024 4396 5030
rect 4344 4966 4396 4972
rect 3700 4684 3752 4690
rect 3700 4626 3752 4632
rect 3792 4684 3844 4690
rect 3792 4626 3844 4632
rect 4356 4622 4384 4966
rect 4344 4616 4396 4622
rect 4344 4558 4396 4564
rect 2610 4380 2918 4389
rect 2610 4378 2616 4380
rect 2672 4378 2696 4380
rect 2752 4378 2776 4380
rect 2832 4378 2856 4380
rect 2912 4378 2918 4380
rect 2672 4326 2674 4378
rect 2854 4326 2856 4378
rect 2610 4324 2616 4326
rect 2672 4324 2696 4326
rect 2752 4324 2776 4326
rect 2832 4324 2856 4326
rect 2912 4324 2918 4326
rect 2610 4315 2918 4324
rect 4816 3534 4844 16546
rect 4908 9042 4936 33050
rect 5000 24342 5028 45526
rect 5080 44192 5132 44198
rect 5080 44134 5132 44140
rect 5092 43382 5120 44134
rect 5080 43376 5132 43382
rect 5080 43318 5132 43324
rect 5172 42560 5224 42566
rect 5172 42502 5224 42508
rect 5080 38752 5132 38758
rect 5080 38694 5132 38700
rect 4988 24336 5040 24342
rect 4988 24278 5040 24284
rect 4988 22976 5040 22982
rect 4988 22918 5040 22924
rect 5000 20874 5028 22918
rect 4988 20868 5040 20874
rect 4988 20810 5040 20816
rect 5092 20466 5120 38694
rect 5184 24818 5212 42502
rect 5540 42084 5592 42090
rect 5540 42026 5592 42032
rect 5552 41138 5580 42026
rect 5540 41132 5592 41138
rect 5540 41074 5592 41080
rect 5540 34128 5592 34134
rect 5540 34070 5592 34076
rect 5552 28150 5580 34070
rect 5724 32972 5776 32978
rect 5724 32914 5776 32920
rect 5540 28144 5592 28150
rect 5540 28086 5592 28092
rect 5552 25838 5580 28086
rect 5540 25832 5592 25838
rect 5540 25774 5592 25780
rect 5172 24812 5224 24818
rect 5172 24754 5224 24760
rect 5080 20460 5132 20466
rect 5080 20402 5132 20408
rect 4896 9036 4948 9042
rect 4896 8978 4948 8984
rect 5736 6458 5764 32914
rect 5920 25906 5948 54538
rect 6012 53650 6040 60046
rect 6380 59090 6408 65554
rect 6368 59084 6420 59090
rect 6368 59026 6420 59032
rect 6184 55276 6236 55282
rect 6184 55218 6236 55224
rect 6092 53984 6144 53990
rect 6092 53926 6144 53932
rect 6000 53644 6052 53650
rect 6000 53586 6052 53592
rect 6012 52698 6040 53586
rect 6000 52692 6052 52698
rect 6000 52634 6052 52640
rect 6104 42090 6132 53926
rect 6092 42084 6144 42090
rect 6092 42026 6144 42032
rect 6092 35624 6144 35630
rect 6092 35566 6144 35572
rect 6000 35148 6052 35154
rect 6000 35090 6052 35096
rect 6012 32434 6040 35090
rect 6104 32502 6132 35566
rect 6092 32496 6144 32502
rect 6092 32438 6144 32444
rect 6000 32428 6052 32434
rect 6000 32370 6052 32376
rect 5908 25900 5960 25906
rect 5908 25842 5960 25848
rect 6196 15978 6224 55218
rect 6276 55072 6328 55078
rect 6276 55014 6328 55020
rect 6288 26246 6316 55014
rect 6380 33590 6408 59026
rect 6472 48006 6500 66098
rect 6564 54602 6592 67594
rect 7610 67484 7918 67493
rect 7610 67482 7616 67484
rect 7672 67482 7696 67484
rect 7752 67482 7776 67484
rect 7832 67482 7856 67484
rect 7912 67482 7918 67484
rect 7672 67430 7674 67482
rect 7854 67430 7856 67482
rect 7610 67428 7616 67430
rect 7672 67428 7696 67430
rect 7752 67428 7776 67430
rect 7832 67428 7856 67430
rect 7912 67428 7918 67430
rect 7610 67419 7918 67428
rect 6950 66940 7258 66949
rect 6950 66938 6956 66940
rect 7012 66938 7036 66940
rect 7092 66938 7116 66940
rect 7172 66938 7196 66940
rect 7252 66938 7258 66940
rect 7012 66886 7014 66938
rect 7194 66886 7196 66938
rect 6950 66884 6956 66886
rect 7012 66884 7036 66886
rect 7092 66884 7116 66886
rect 7172 66884 7196 66886
rect 7252 66884 7258 66886
rect 6950 66875 7258 66884
rect 8116 66768 8168 66774
rect 8116 66710 8168 66716
rect 7472 66632 7524 66638
rect 7472 66574 7524 66580
rect 6950 65852 7258 65861
rect 6950 65850 6956 65852
rect 7012 65850 7036 65852
rect 7092 65850 7116 65852
rect 7172 65850 7196 65852
rect 7252 65850 7258 65852
rect 7012 65798 7014 65850
rect 7194 65798 7196 65850
rect 6950 65796 6956 65798
rect 7012 65796 7036 65798
rect 7092 65796 7116 65798
rect 7172 65796 7196 65798
rect 7252 65796 7258 65798
rect 6950 65787 7258 65796
rect 6950 64764 7258 64773
rect 6950 64762 6956 64764
rect 7012 64762 7036 64764
rect 7092 64762 7116 64764
rect 7172 64762 7196 64764
rect 7252 64762 7258 64764
rect 7012 64710 7014 64762
rect 7194 64710 7196 64762
rect 6950 64708 6956 64710
rect 7012 64708 7036 64710
rect 7092 64708 7116 64710
rect 7172 64708 7196 64710
rect 7252 64708 7258 64710
rect 6950 64699 7258 64708
rect 6950 63676 7258 63685
rect 6950 63674 6956 63676
rect 7012 63674 7036 63676
rect 7092 63674 7116 63676
rect 7172 63674 7196 63676
rect 7252 63674 7258 63676
rect 7012 63622 7014 63674
rect 7194 63622 7196 63674
rect 6950 63620 6956 63622
rect 7012 63620 7036 63622
rect 7092 63620 7116 63622
rect 7172 63620 7196 63622
rect 7252 63620 7258 63622
rect 6950 63611 7258 63620
rect 6828 62892 6880 62898
rect 6828 62834 6880 62840
rect 6736 59016 6788 59022
rect 6736 58958 6788 58964
rect 6748 58614 6776 58958
rect 6736 58608 6788 58614
rect 6736 58550 6788 58556
rect 6748 54738 6776 58550
rect 6736 54732 6788 54738
rect 6736 54674 6788 54680
rect 6552 54596 6604 54602
rect 6552 54538 6604 54544
rect 6564 53990 6592 54538
rect 6748 54534 6776 54674
rect 6736 54528 6788 54534
rect 6736 54470 6788 54476
rect 6552 53984 6604 53990
rect 6552 53926 6604 53932
rect 6552 52692 6604 52698
rect 6552 52634 6604 52640
rect 6460 48000 6512 48006
rect 6460 47942 6512 47948
rect 6460 45280 6512 45286
rect 6460 45222 6512 45228
rect 6472 44878 6500 45222
rect 6460 44872 6512 44878
rect 6460 44814 6512 44820
rect 6460 38480 6512 38486
rect 6460 38422 6512 38428
rect 6472 35086 6500 38422
rect 6460 35080 6512 35086
rect 6460 35022 6512 35028
rect 6460 34944 6512 34950
rect 6460 34886 6512 34892
rect 6368 33584 6420 33590
rect 6368 33526 6420 33532
rect 6380 33386 6408 33526
rect 6368 33380 6420 33386
rect 6368 33322 6420 33328
rect 6368 32428 6420 32434
rect 6368 32370 6420 32376
rect 6276 26240 6328 26246
rect 6276 26182 6328 26188
rect 6276 19712 6328 19718
rect 6276 19654 6328 19660
rect 6184 15972 6236 15978
rect 6184 15914 6236 15920
rect 6092 11076 6144 11082
rect 6092 11018 6144 11024
rect 6104 7342 6132 11018
rect 6092 7336 6144 7342
rect 6092 7278 6144 7284
rect 5724 6452 5776 6458
rect 5724 6394 5776 6400
rect 6104 4622 6132 7278
rect 6184 6656 6236 6662
rect 6184 6598 6236 6604
rect 6196 6322 6224 6598
rect 6184 6316 6236 6322
rect 6184 6258 6236 6264
rect 6092 4616 6144 4622
rect 6092 4558 6144 4564
rect 6288 4554 6316 19654
rect 6380 16114 6408 32370
rect 6472 32366 6500 34886
rect 6460 32360 6512 32366
rect 6460 32302 6512 32308
rect 6460 26240 6512 26246
rect 6460 26182 6512 26188
rect 6472 26042 6500 26182
rect 6460 26036 6512 26042
rect 6460 25978 6512 25984
rect 6368 16108 6420 16114
rect 6368 16050 6420 16056
rect 6276 4548 6328 4554
rect 6276 4490 6328 4496
rect 6472 4146 6500 25978
rect 6564 16658 6592 52634
rect 6840 51338 6868 62834
rect 6950 62588 7258 62597
rect 6950 62586 6956 62588
rect 7012 62586 7036 62588
rect 7092 62586 7116 62588
rect 7172 62586 7196 62588
rect 7252 62586 7258 62588
rect 7012 62534 7014 62586
rect 7194 62534 7196 62586
rect 6950 62532 6956 62534
rect 7012 62532 7036 62534
rect 7092 62532 7116 62534
rect 7172 62532 7196 62534
rect 7252 62532 7258 62534
rect 6950 62523 7258 62532
rect 7380 62280 7432 62286
rect 7380 62222 7432 62228
rect 6950 61500 7258 61509
rect 6950 61498 6956 61500
rect 7012 61498 7036 61500
rect 7092 61498 7116 61500
rect 7172 61498 7196 61500
rect 7252 61498 7258 61500
rect 7012 61446 7014 61498
rect 7194 61446 7196 61498
rect 6950 61444 6956 61446
rect 7012 61444 7036 61446
rect 7092 61444 7116 61446
rect 7172 61444 7196 61446
rect 7252 61444 7258 61446
rect 6950 61435 7258 61444
rect 6950 60412 7258 60421
rect 6950 60410 6956 60412
rect 7012 60410 7036 60412
rect 7092 60410 7116 60412
rect 7172 60410 7196 60412
rect 7252 60410 7258 60412
rect 7012 60358 7014 60410
rect 7194 60358 7196 60410
rect 6950 60356 6956 60358
rect 7012 60356 7036 60358
rect 7092 60356 7116 60358
rect 7172 60356 7196 60358
rect 7252 60356 7258 60358
rect 6950 60347 7258 60356
rect 6950 59324 7258 59333
rect 6950 59322 6956 59324
rect 7012 59322 7036 59324
rect 7092 59322 7116 59324
rect 7172 59322 7196 59324
rect 7252 59322 7258 59324
rect 7012 59270 7014 59322
rect 7194 59270 7196 59322
rect 6950 59268 6956 59270
rect 7012 59268 7036 59270
rect 7092 59268 7116 59270
rect 7172 59268 7196 59270
rect 7252 59268 7258 59270
rect 6950 59259 7258 59268
rect 6950 58236 7258 58245
rect 6950 58234 6956 58236
rect 7012 58234 7036 58236
rect 7092 58234 7116 58236
rect 7172 58234 7196 58236
rect 7252 58234 7258 58236
rect 7012 58182 7014 58234
rect 7194 58182 7196 58234
rect 6950 58180 6956 58182
rect 7012 58180 7036 58182
rect 7092 58180 7116 58182
rect 7172 58180 7196 58182
rect 7252 58180 7258 58182
rect 6950 58171 7258 58180
rect 6950 57148 7258 57157
rect 6950 57146 6956 57148
rect 7012 57146 7036 57148
rect 7092 57146 7116 57148
rect 7172 57146 7196 57148
rect 7252 57146 7258 57148
rect 7012 57094 7014 57146
rect 7194 57094 7196 57146
rect 6950 57092 6956 57094
rect 7012 57092 7036 57094
rect 7092 57092 7116 57094
rect 7172 57092 7196 57094
rect 7252 57092 7258 57094
rect 6950 57083 7258 57092
rect 6950 56060 7258 56069
rect 6950 56058 6956 56060
rect 7012 56058 7036 56060
rect 7092 56058 7116 56060
rect 7172 56058 7196 56060
rect 7252 56058 7258 56060
rect 7012 56006 7014 56058
rect 7194 56006 7196 56058
rect 6950 56004 6956 56006
rect 7012 56004 7036 56006
rect 7092 56004 7116 56006
rect 7172 56004 7196 56006
rect 7252 56004 7258 56006
rect 6950 55995 7258 56004
rect 6950 54972 7258 54981
rect 6950 54970 6956 54972
rect 7012 54970 7036 54972
rect 7092 54970 7116 54972
rect 7172 54970 7196 54972
rect 7252 54970 7258 54972
rect 7012 54918 7014 54970
rect 7194 54918 7196 54970
rect 6950 54916 6956 54918
rect 7012 54916 7036 54918
rect 7092 54916 7116 54918
rect 7172 54916 7196 54918
rect 7252 54916 7258 54918
rect 6950 54907 7258 54916
rect 7104 54528 7156 54534
rect 7104 54470 7156 54476
rect 7116 54330 7144 54470
rect 7104 54324 7156 54330
rect 7104 54266 7156 54272
rect 6950 53884 7258 53893
rect 6950 53882 6956 53884
rect 7012 53882 7036 53884
rect 7092 53882 7116 53884
rect 7172 53882 7196 53884
rect 7252 53882 7258 53884
rect 7012 53830 7014 53882
rect 7194 53830 7196 53882
rect 6950 53828 6956 53830
rect 7012 53828 7036 53830
rect 7092 53828 7116 53830
rect 7172 53828 7196 53830
rect 7252 53828 7258 53830
rect 6950 53819 7258 53828
rect 7288 53440 7340 53446
rect 7288 53382 7340 53388
rect 6950 52796 7258 52805
rect 6950 52794 6956 52796
rect 7012 52794 7036 52796
rect 7092 52794 7116 52796
rect 7172 52794 7196 52796
rect 7252 52794 7258 52796
rect 7012 52742 7014 52794
rect 7194 52742 7196 52794
rect 6950 52740 6956 52742
rect 7012 52740 7036 52742
rect 7092 52740 7116 52742
rect 7172 52740 7196 52742
rect 7252 52740 7258 52742
rect 6950 52731 7258 52740
rect 6950 51708 7258 51717
rect 6950 51706 6956 51708
rect 7012 51706 7036 51708
rect 7092 51706 7116 51708
rect 7172 51706 7196 51708
rect 7252 51706 7258 51708
rect 7012 51654 7014 51706
rect 7194 51654 7196 51706
rect 6950 51652 6956 51654
rect 7012 51652 7036 51654
rect 7092 51652 7116 51654
rect 7172 51652 7196 51654
rect 7252 51652 7258 51654
rect 6950 51643 7258 51652
rect 6828 51332 6880 51338
rect 6828 51274 6880 51280
rect 6736 50244 6788 50250
rect 6736 50186 6788 50192
rect 6748 44878 6776 50186
rect 6736 44872 6788 44878
rect 6736 44814 6788 44820
rect 6736 35284 6788 35290
rect 6736 35226 6788 35232
rect 6644 35216 6696 35222
rect 6748 35193 6776 35226
rect 6644 35158 6696 35164
rect 6734 35184 6790 35193
rect 6656 32434 6684 35158
rect 6734 35119 6790 35128
rect 6644 32428 6696 32434
rect 6644 32370 6696 32376
rect 6736 32428 6788 32434
rect 6736 32370 6788 32376
rect 6644 25900 6696 25906
rect 6644 25842 6696 25848
rect 6656 22574 6684 25842
rect 6644 22568 6696 22574
rect 6644 22510 6696 22516
rect 6552 16652 6604 16658
rect 6552 16594 6604 16600
rect 6748 5794 6776 32370
rect 6840 29102 6868 51274
rect 6950 50620 7258 50629
rect 6950 50618 6956 50620
rect 7012 50618 7036 50620
rect 7092 50618 7116 50620
rect 7172 50618 7196 50620
rect 7252 50618 7258 50620
rect 7012 50566 7014 50618
rect 7194 50566 7196 50618
rect 6950 50564 6956 50566
rect 7012 50564 7036 50566
rect 7092 50564 7116 50566
rect 7172 50564 7196 50566
rect 7252 50564 7258 50566
rect 6950 50555 7258 50564
rect 7300 49910 7328 53382
rect 7288 49904 7340 49910
rect 7288 49846 7340 49852
rect 6950 49532 7258 49541
rect 6950 49530 6956 49532
rect 7012 49530 7036 49532
rect 7092 49530 7116 49532
rect 7172 49530 7196 49532
rect 7252 49530 7258 49532
rect 7012 49478 7014 49530
rect 7194 49478 7196 49530
rect 6950 49476 6956 49478
rect 7012 49476 7036 49478
rect 7092 49476 7116 49478
rect 7172 49476 7196 49478
rect 7252 49476 7258 49478
rect 6950 49467 7258 49476
rect 6950 48444 7258 48453
rect 6950 48442 6956 48444
rect 7012 48442 7036 48444
rect 7092 48442 7116 48444
rect 7172 48442 7196 48444
rect 7252 48442 7258 48444
rect 7012 48390 7014 48442
rect 7194 48390 7196 48442
rect 6950 48388 6956 48390
rect 7012 48388 7036 48390
rect 7092 48388 7116 48390
rect 7172 48388 7196 48390
rect 7252 48388 7258 48390
rect 6950 48379 7258 48388
rect 6950 47356 7258 47365
rect 6950 47354 6956 47356
rect 7012 47354 7036 47356
rect 7092 47354 7116 47356
rect 7172 47354 7196 47356
rect 7252 47354 7258 47356
rect 7012 47302 7014 47354
rect 7194 47302 7196 47354
rect 6950 47300 6956 47302
rect 7012 47300 7036 47302
rect 7092 47300 7116 47302
rect 7172 47300 7196 47302
rect 7252 47300 7258 47302
rect 6950 47291 7258 47300
rect 6950 46268 7258 46277
rect 6950 46266 6956 46268
rect 7012 46266 7036 46268
rect 7092 46266 7116 46268
rect 7172 46266 7196 46268
rect 7252 46266 7258 46268
rect 7012 46214 7014 46266
rect 7194 46214 7196 46266
rect 6950 46212 6956 46214
rect 7012 46212 7036 46214
rect 7092 46212 7116 46214
rect 7172 46212 7196 46214
rect 7252 46212 7258 46214
rect 6950 46203 7258 46212
rect 6950 45180 7258 45189
rect 6950 45178 6956 45180
rect 7012 45178 7036 45180
rect 7092 45178 7116 45180
rect 7172 45178 7196 45180
rect 7252 45178 7258 45180
rect 7012 45126 7014 45178
rect 7194 45126 7196 45178
rect 6950 45124 6956 45126
rect 7012 45124 7036 45126
rect 7092 45124 7116 45126
rect 7172 45124 7196 45126
rect 7252 45124 7258 45126
rect 6950 45115 7258 45124
rect 6950 44092 7258 44101
rect 6950 44090 6956 44092
rect 7012 44090 7036 44092
rect 7092 44090 7116 44092
rect 7172 44090 7196 44092
rect 7252 44090 7258 44092
rect 7012 44038 7014 44090
rect 7194 44038 7196 44090
rect 6950 44036 6956 44038
rect 7012 44036 7036 44038
rect 7092 44036 7116 44038
rect 7172 44036 7196 44038
rect 7252 44036 7258 44038
rect 6950 44027 7258 44036
rect 6950 43004 7258 43013
rect 6950 43002 6956 43004
rect 7012 43002 7036 43004
rect 7092 43002 7116 43004
rect 7172 43002 7196 43004
rect 7252 43002 7258 43004
rect 7012 42950 7014 43002
rect 7194 42950 7196 43002
rect 6950 42948 6956 42950
rect 7012 42948 7036 42950
rect 7092 42948 7116 42950
rect 7172 42948 7196 42950
rect 7252 42948 7258 42950
rect 6950 42939 7258 42948
rect 6950 41916 7258 41925
rect 6950 41914 6956 41916
rect 7012 41914 7036 41916
rect 7092 41914 7116 41916
rect 7172 41914 7196 41916
rect 7252 41914 7258 41916
rect 7012 41862 7014 41914
rect 7194 41862 7196 41914
rect 6950 41860 6956 41862
rect 7012 41860 7036 41862
rect 7092 41860 7116 41862
rect 7172 41860 7196 41862
rect 7252 41860 7258 41862
rect 6950 41851 7258 41860
rect 6950 40828 7258 40837
rect 6950 40826 6956 40828
rect 7012 40826 7036 40828
rect 7092 40826 7116 40828
rect 7172 40826 7196 40828
rect 7252 40826 7258 40828
rect 7012 40774 7014 40826
rect 7194 40774 7196 40826
rect 6950 40772 6956 40774
rect 7012 40772 7036 40774
rect 7092 40772 7116 40774
rect 7172 40772 7196 40774
rect 7252 40772 7258 40774
rect 6950 40763 7258 40772
rect 6950 39740 7258 39749
rect 6950 39738 6956 39740
rect 7012 39738 7036 39740
rect 7092 39738 7116 39740
rect 7172 39738 7196 39740
rect 7252 39738 7258 39740
rect 7012 39686 7014 39738
rect 7194 39686 7196 39738
rect 6950 39684 6956 39686
rect 7012 39684 7036 39686
rect 7092 39684 7116 39686
rect 7172 39684 7196 39686
rect 7252 39684 7258 39686
rect 6950 39675 7258 39684
rect 6950 38652 7258 38661
rect 6950 38650 6956 38652
rect 7012 38650 7036 38652
rect 7092 38650 7116 38652
rect 7172 38650 7196 38652
rect 7252 38650 7258 38652
rect 7012 38598 7014 38650
rect 7194 38598 7196 38650
rect 6950 38596 6956 38598
rect 7012 38596 7036 38598
rect 7092 38596 7116 38598
rect 7172 38596 7196 38598
rect 7252 38596 7258 38598
rect 6950 38587 7258 38596
rect 6950 37564 7258 37573
rect 6950 37562 6956 37564
rect 7012 37562 7036 37564
rect 7092 37562 7116 37564
rect 7172 37562 7196 37564
rect 7252 37562 7258 37564
rect 7012 37510 7014 37562
rect 7194 37510 7196 37562
rect 6950 37508 6956 37510
rect 7012 37508 7036 37510
rect 7092 37508 7116 37510
rect 7172 37508 7196 37510
rect 7252 37508 7258 37510
rect 6950 37499 7258 37508
rect 6950 36476 7258 36485
rect 6950 36474 6956 36476
rect 7012 36474 7036 36476
rect 7092 36474 7116 36476
rect 7172 36474 7196 36476
rect 7252 36474 7258 36476
rect 7012 36422 7014 36474
rect 7194 36422 7196 36474
rect 6950 36420 6956 36422
rect 7012 36420 7036 36422
rect 7092 36420 7116 36422
rect 7172 36420 7196 36422
rect 7252 36420 7258 36422
rect 6950 36411 7258 36420
rect 6950 35388 7258 35397
rect 6950 35386 6956 35388
rect 7012 35386 7036 35388
rect 7092 35386 7116 35388
rect 7172 35386 7196 35388
rect 7252 35386 7258 35388
rect 7012 35334 7014 35386
rect 7194 35334 7196 35386
rect 6950 35332 6956 35334
rect 7012 35332 7036 35334
rect 7092 35332 7116 35334
rect 7172 35332 7196 35334
rect 7252 35332 7258 35334
rect 6950 35323 7258 35332
rect 7196 35284 7248 35290
rect 7196 35226 7248 35232
rect 7208 34678 7236 35226
rect 7196 34672 7248 34678
rect 7196 34614 7248 34620
rect 6950 34300 7258 34309
rect 6950 34298 6956 34300
rect 7012 34298 7036 34300
rect 7092 34298 7116 34300
rect 7172 34298 7196 34300
rect 7252 34298 7258 34300
rect 7012 34246 7014 34298
rect 7194 34246 7196 34298
rect 6950 34244 6956 34246
rect 7012 34244 7036 34246
rect 7092 34244 7116 34246
rect 7172 34244 7196 34246
rect 7252 34244 7258 34246
rect 6950 34235 7258 34244
rect 6950 33212 7258 33221
rect 6950 33210 6956 33212
rect 7012 33210 7036 33212
rect 7092 33210 7116 33212
rect 7172 33210 7196 33212
rect 7252 33210 7258 33212
rect 7012 33158 7014 33210
rect 7194 33158 7196 33210
rect 6950 33156 6956 33158
rect 7012 33156 7036 33158
rect 7092 33156 7116 33158
rect 7172 33156 7196 33158
rect 7252 33156 7258 33158
rect 6950 33147 7258 33156
rect 6950 32124 7258 32133
rect 6950 32122 6956 32124
rect 7012 32122 7036 32124
rect 7092 32122 7116 32124
rect 7172 32122 7196 32124
rect 7252 32122 7258 32124
rect 7012 32070 7014 32122
rect 7194 32070 7196 32122
rect 6950 32068 6956 32070
rect 7012 32068 7036 32070
rect 7092 32068 7116 32070
rect 7172 32068 7196 32070
rect 7252 32068 7258 32070
rect 6950 32059 7258 32068
rect 6950 31036 7258 31045
rect 6950 31034 6956 31036
rect 7012 31034 7036 31036
rect 7092 31034 7116 31036
rect 7172 31034 7196 31036
rect 7252 31034 7258 31036
rect 7012 30982 7014 31034
rect 7194 30982 7196 31034
rect 6950 30980 6956 30982
rect 7012 30980 7036 30982
rect 7092 30980 7116 30982
rect 7172 30980 7196 30982
rect 7252 30980 7258 30982
rect 6950 30971 7258 30980
rect 6950 29948 7258 29957
rect 6950 29946 6956 29948
rect 7012 29946 7036 29948
rect 7092 29946 7116 29948
rect 7172 29946 7196 29948
rect 7252 29946 7258 29948
rect 7012 29894 7014 29946
rect 7194 29894 7196 29946
rect 6950 29892 6956 29894
rect 7012 29892 7036 29894
rect 7092 29892 7116 29894
rect 7172 29892 7196 29894
rect 7252 29892 7258 29894
rect 6950 29883 7258 29892
rect 6828 29096 6880 29102
rect 6828 29038 6880 29044
rect 6950 28860 7258 28869
rect 6950 28858 6956 28860
rect 7012 28858 7036 28860
rect 7092 28858 7116 28860
rect 7172 28858 7196 28860
rect 7252 28858 7258 28860
rect 7012 28806 7014 28858
rect 7194 28806 7196 28858
rect 6950 28804 6956 28806
rect 7012 28804 7036 28806
rect 7092 28804 7116 28806
rect 7172 28804 7196 28806
rect 7252 28804 7258 28806
rect 6950 28795 7258 28804
rect 6950 27772 7258 27781
rect 6950 27770 6956 27772
rect 7012 27770 7036 27772
rect 7092 27770 7116 27772
rect 7172 27770 7196 27772
rect 7252 27770 7258 27772
rect 7012 27718 7014 27770
rect 7194 27718 7196 27770
rect 6950 27716 6956 27718
rect 7012 27716 7036 27718
rect 7092 27716 7116 27718
rect 7172 27716 7196 27718
rect 7252 27716 7258 27718
rect 6950 27707 7258 27716
rect 6950 26684 7258 26693
rect 6950 26682 6956 26684
rect 7012 26682 7036 26684
rect 7092 26682 7116 26684
rect 7172 26682 7196 26684
rect 7252 26682 7258 26684
rect 7012 26630 7014 26682
rect 7194 26630 7196 26682
rect 6950 26628 6956 26630
rect 7012 26628 7036 26630
rect 7092 26628 7116 26630
rect 7172 26628 7196 26630
rect 7252 26628 7258 26630
rect 6950 26619 7258 26628
rect 6950 25596 7258 25605
rect 6950 25594 6956 25596
rect 7012 25594 7036 25596
rect 7092 25594 7116 25596
rect 7172 25594 7196 25596
rect 7252 25594 7258 25596
rect 7012 25542 7014 25594
rect 7194 25542 7196 25594
rect 6950 25540 6956 25542
rect 7012 25540 7036 25542
rect 7092 25540 7116 25542
rect 7172 25540 7196 25542
rect 7252 25540 7258 25542
rect 6950 25531 7258 25540
rect 7300 24750 7328 49846
rect 7392 34785 7420 62222
rect 7484 59158 7512 66574
rect 7610 66396 7918 66405
rect 7610 66394 7616 66396
rect 7672 66394 7696 66396
rect 7752 66394 7776 66396
rect 7832 66394 7856 66396
rect 7912 66394 7918 66396
rect 7672 66342 7674 66394
rect 7854 66342 7856 66394
rect 7610 66340 7616 66342
rect 7672 66340 7696 66342
rect 7752 66340 7776 66342
rect 7832 66340 7856 66342
rect 7912 66340 7918 66342
rect 7610 66331 7918 66340
rect 8128 65521 8156 66710
rect 8114 65512 8170 65521
rect 8114 65447 8170 65456
rect 7610 65308 7918 65317
rect 7610 65306 7616 65308
rect 7672 65306 7696 65308
rect 7752 65306 7776 65308
rect 7832 65306 7856 65308
rect 7912 65306 7918 65308
rect 7672 65254 7674 65306
rect 7854 65254 7856 65306
rect 7610 65252 7616 65254
rect 7672 65252 7696 65254
rect 7752 65252 7776 65254
rect 7832 65252 7856 65254
rect 7912 65252 7918 65254
rect 7610 65243 7918 65252
rect 7840 64864 7892 64870
rect 7840 64806 7892 64812
rect 7852 64462 7880 64806
rect 8116 64592 8168 64598
rect 8116 64534 8168 64540
rect 7840 64456 7892 64462
rect 7840 64398 7892 64404
rect 7610 64220 7918 64229
rect 7610 64218 7616 64220
rect 7672 64218 7696 64220
rect 7752 64218 7776 64220
rect 7832 64218 7856 64220
rect 7912 64218 7918 64220
rect 7672 64166 7674 64218
rect 7854 64166 7856 64218
rect 7610 64164 7616 64166
rect 7672 64164 7696 64166
rect 7752 64164 7776 64166
rect 7832 64164 7856 64166
rect 7912 64164 7918 64166
rect 7610 64155 7918 64164
rect 7610 63132 7918 63141
rect 7610 63130 7616 63132
rect 7672 63130 7696 63132
rect 7752 63130 7776 63132
rect 7832 63130 7856 63132
rect 7912 63130 7918 63132
rect 7672 63078 7674 63130
rect 7854 63078 7856 63130
rect 7610 63076 7616 63078
rect 7672 63076 7696 63078
rect 7752 63076 7776 63078
rect 7832 63076 7856 63078
rect 7912 63076 7918 63078
rect 7610 63067 7918 63076
rect 7610 62044 7918 62053
rect 7610 62042 7616 62044
rect 7672 62042 7696 62044
rect 7752 62042 7776 62044
rect 7832 62042 7856 62044
rect 7912 62042 7918 62044
rect 7672 61990 7674 62042
rect 7854 61990 7856 62042
rect 7610 61988 7616 61990
rect 7672 61988 7696 61990
rect 7752 61988 7776 61990
rect 7832 61988 7856 61990
rect 7912 61988 7918 61990
rect 7610 61979 7918 61988
rect 8024 61124 8076 61130
rect 8024 61066 8076 61072
rect 7610 60956 7918 60965
rect 7610 60954 7616 60956
rect 7672 60954 7696 60956
rect 7752 60954 7776 60956
rect 7832 60954 7856 60956
rect 7912 60954 7918 60956
rect 7672 60902 7674 60954
rect 7854 60902 7856 60954
rect 7610 60900 7616 60902
rect 7672 60900 7696 60902
rect 7752 60900 7776 60902
rect 7832 60900 7856 60902
rect 7912 60900 7918 60902
rect 7610 60891 7918 60900
rect 7610 59868 7918 59877
rect 7610 59866 7616 59868
rect 7672 59866 7696 59868
rect 7752 59866 7776 59868
rect 7832 59866 7856 59868
rect 7912 59866 7918 59868
rect 7672 59814 7674 59866
rect 7854 59814 7856 59866
rect 7610 59812 7616 59814
rect 7672 59812 7696 59814
rect 7752 59812 7776 59814
rect 7832 59812 7856 59814
rect 7912 59812 7918 59814
rect 7610 59803 7918 59812
rect 7472 59152 7524 59158
rect 7472 59094 7524 59100
rect 7610 58780 7918 58789
rect 7610 58778 7616 58780
rect 7672 58778 7696 58780
rect 7752 58778 7776 58780
rect 7832 58778 7856 58780
rect 7912 58778 7918 58780
rect 7672 58726 7674 58778
rect 7854 58726 7856 58778
rect 7610 58724 7616 58726
rect 7672 58724 7696 58726
rect 7752 58724 7776 58726
rect 7832 58724 7856 58726
rect 7912 58724 7918 58726
rect 7610 58715 7918 58724
rect 7610 57692 7918 57701
rect 7610 57690 7616 57692
rect 7672 57690 7696 57692
rect 7752 57690 7776 57692
rect 7832 57690 7856 57692
rect 7912 57690 7918 57692
rect 7672 57638 7674 57690
rect 7854 57638 7856 57690
rect 7610 57636 7616 57638
rect 7672 57636 7696 57638
rect 7752 57636 7776 57638
rect 7832 57636 7856 57638
rect 7912 57636 7918 57638
rect 7610 57627 7918 57636
rect 7610 56604 7918 56613
rect 7610 56602 7616 56604
rect 7672 56602 7696 56604
rect 7752 56602 7776 56604
rect 7832 56602 7856 56604
rect 7912 56602 7918 56604
rect 7672 56550 7674 56602
rect 7854 56550 7856 56602
rect 7610 56548 7616 56550
rect 7672 56548 7696 56550
rect 7752 56548 7776 56550
rect 7832 56548 7856 56550
rect 7912 56548 7918 56550
rect 7610 56539 7918 56548
rect 7610 55516 7918 55525
rect 7610 55514 7616 55516
rect 7672 55514 7696 55516
rect 7752 55514 7776 55516
rect 7832 55514 7856 55516
rect 7912 55514 7918 55516
rect 7672 55462 7674 55514
rect 7854 55462 7856 55514
rect 7610 55460 7616 55462
rect 7672 55460 7696 55462
rect 7752 55460 7776 55462
rect 7832 55460 7856 55462
rect 7912 55460 7918 55462
rect 7610 55451 7918 55460
rect 7472 54732 7524 54738
rect 7472 54674 7524 54680
rect 7484 35834 7512 54674
rect 7610 54428 7918 54437
rect 7610 54426 7616 54428
rect 7672 54426 7696 54428
rect 7752 54426 7776 54428
rect 7832 54426 7856 54428
rect 7912 54426 7918 54428
rect 7672 54374 7674 54426
rect 7854 54374 7856 54426
rect 7610 54372 7616 54374
rect 7672 54372 7696 54374
rect 7752 54372 7776 54374
rect 7832 54372 7856 54374
rect 7912 54372 7918 54374
rect 7610 54363 7918 54372
rect 7610 53340 7918 53349
rect 7610 53338 7616 53340
rect 7672 53338 7696 53340
rect 7752 53338 7776 53340
rect 7832 53338 7856 53340
rect 7912 53338 7918 53340
rect 7672 53286 7674 53338
rect 7854 53286 7856 53338
rect 7610 53284 7616 53286
rect 7672 53284 7696 53286
rect 7752 53284 7776 53286
rect 7832 53284 7856 53286
rect 7912 53284 7918 53286
rect 7610 53275 7918 53284
rect 7610 52252 7918 52261
rect 7610 52250 7616 52252
rect 7672 52250 7696 52252
rect 7752 52250 7776 52252
rect 7832 52250 7856 52252
rect 7912 52250 7918 52252
rect 7672 52198 7674 52250
rect 7854 52198 7856 52250
rect 7610 52196 7616 52198
rect 7672 52196 7696 52198
rect 7752 52196 7776 52198
rect 7832 52196 7856 52198
rect 7912 52196 7918 52198
rect 7610 52187 7918 52196
rect 7610 51164 7918 51173
rect 7610 51162 7616 51164
rect 7672 51162 7696 51164
rect 7752 51162 7776 51164
rect 7832 51162 7856 51164
rect 7912 51162 7918 51164
rect 7672 51110 7674 51162
rect 7854 51110 7856 51162
rect 7610 51108 7616 51110
rect 7672 51108 7696 51110
rect 7752 51108 7776 51110
rect 7832 51108 7856 51110
rect 7912 51108 7918 51110
rect 7610 51099 7918 51108
rect 7932 50924 7984 50930
rect 7932 50866 7984 50872
rect 7944 50266 7972 50866
rect 8036 50386 8064 61066
rect 8128 60518 8156 64534
rect 8956 62830 8984 67866
rect 9600 65550 9628 69294
rect 11950 69116 12258 69125
rect 11950 69114 11956 69116
rect 12012 69114 12036 69116
rect 12092 69114 12116 69116
rect 12172 69114 12196 69116
rect 12252 69114 12258 69116
rect 12012 69062 12014 69114
rect 12194 69062 12196 69114
rect 11950 69060 11956 69062
rect 12012 69060 12036 69062
rect 12092 69060 12116 69062
rect 12172 69060 12196 69062
rect 12252 69060 12258 69062
rect 11950 69051 12258 69060
rect 16950 69116 17258 69125
rect 16950 69114 16956 69116
rect 17012 69114 17036 69116
rect 17092 69114 17116 69116
rect 17172 69114 17196 69116
rect 17252 69114 17258 69116
rect 17012 69062 17014 69114
rect 17194 69062 17196 69114
rect 16950 69060 16956 69062
rect 17012 69060 17036 69062
rect 17092 69060 17116 69062
rect 17172 69060 17196 69062
rect 17252 69060 17258 69062
rect 16950 69051 17258 69060
rect 21950 69116 22258 69125
rect 21950 69114 21956 69116
rect 22012 69114 22036 69116
rect 22092 69114 22116 69116
rect 22172 69114 22196 69116
rect 22252 69114 22258 69116
rect 22012 69062 22014 69114
rect 22194 69062 22196 69114
rect 21950 69060 21956 69062
rect 22012 69060 22036 69062
rect 22092 69060 22116 69062
rect 22172 69060 22196 69062
rect 22252 69060 22258 69062
rect 21950 69051 22258 69060
rect 11428 68808 11480 68814
rect 11428 68750 11480 68756
rect 13176 68808 13228 68814
rect 13176 68750 13228 68756
rect 15568 68808 15620 68814
rect 15568 68750 15620 68756
rect 10508 67108 10560 67114
rect 10508 67050 10560 67056
rect 10416 66632 10468 66638
rect 10416 66574 10468 66580
rect 9588 65544 9640 65550
rect 9588 65486 9640 65492
rect 8944 62824 8996 62830
rect 8944 62766 8996 62772
rect 9588 62688 9640 62694
rect 9588 62630 9640 62636
rect 8944 61192 8996 61198
rect 8944 61134 8996 61140
rect 9220 61192 9272 61198
rect 9220 61134 9272 61140
rect 8484 60716 8536 60722
rect 8484 60658 8536 60664
rect 8116 60512 8168 60518
rect 8116 60454 8168 60460
rect 8024 50380 8076 50386
rect 8024 50322 8076 50328
rect 7944 50238 8064 50266
rect 7610 50076 7918 50085
rect 7610 50074 7616 50076
rect 7672 50074 7696 50076
rect 7752 50074 7776 50076
rect 7832 50074 7856 50076
rect 7912 50074 7918 50076
rect 7672 50022 7674 50074
rect 7854 50022 7856 50074
rect 7610 50020 7616 50022
rect 7672 50020 7696 50022
rect 7752 50020 7776 50022
rect 7832 50020 7856 50022
rect 7912 50020 7918 50022
rect 7610 50011 7918 50020
rect 7610 48988 7918 48997
rect 7610 48986 7616 48988
rect 7672 48986 7696 48988
rect 7752 48986 7776 48988
rect 7832 48986 7856 48988
rect 7912 48986 7918 48988
rect 7672 48934 7674 48986
rect 7854 48934 7856 48986
rect 7610 48932 7616 48934
rect 7672 48932 7696 48934
rect 7752 48932 7776 48934
rect 7832 48932 7856 48934
rect 7912 48932 7918 48934
rect 7610 48923 7918 48932
rect 7610 47900 7918 47909
rect 7610 47898 7616 47900
rect 7672 47898 7696 47900
rect 7752 47898 7776 47900
rect 7832 47898 7856 47900
rect 7912 47898 7918 47900
rect 7672 47846 7674 47898
rect 7854 47846 7856 47898
rect 7610 47844 7616 47846
rect 7672 47844 7696 47846
rect 7752 47844 7776 47846
rect 7832 47844 7856 47846
rect 7912 47844 7918 47846
rect 7610 47835 7918 47844
rect 7610 46812 7918 46821
rect 7610 46810 7616 46812
rect 7672 46810 7696 46812
rect 7752 46810 7776 46812
rect 7832 46810 7856 46812
rect 7912 46810 7918 46812
rect 7672 46758 7674 46810
rect 7854 46758 7856 46810
rect 7610 46756 7616 46758
rect 7672 46756 7696 46758
rect 7752 46756 7776 46758
rect 7832 46756 7856 46758
rect 7912 46756 7918 46758
rect 7610 46747 7918 46756
rect 7610 45724 7918 45733
rect 7610 45722 7616 45724
rect 7672 45722 7696 45724
rect 7752 45722 7776 45724
rect 7832 45722 7856 45724
rect 7912 45722 7918 45724
rect 7672 45670 7674 45722
rect 7854 45670 7856 45722
rect 7610 45668 7616 45670
rect 7672 45668 7696 45670
rect 7752 45668 7776 45670
rect 7832 45668 7856 45670
rect 7912 45668 7918 45670
rect 7610 45659 7918 45668
rect 7610 44636 7918 44645
rect 7610 44634 7616 44636
rect 7672 44634 7696 44636
rect 7752 44634 7776 44636
rect 7832 44634 7856 44636
rect 7912 44634 7918 44636
rect 7672 44582 7674 44634
rect 7854 44582 7856 44634
rect 7610 44580 7616 44582
rect 7672 44580 7696 44582
rect 7752 44580 7776 44582
rect 7832 44580 7856 44582
rect 7912 44580 7918 44582
rect 7610 44571 7918 44580
rect 7610 43548 7918 43557
rect 7610 43546 7616 43548
rect 7672 43546 7696 43548
rect 7752 43546 7776 43548
rect 7832 43546 7856 43548
rect 7912 43546 7918 43548
rect 7672 43494 7674 43546
rect 7854 43494 7856 43546
rect 7610 43492 7616 43494
rect 7672 43492 7696 43494
rect 7752 43492 7776 43494
rect 7832 43492 7856 43494
rect 7912 43492 7918 43494
rect 7610 43483 7918 43492
rect 7610 42460 7918 42469
rect 7610 42458 7616 42460
rect 7672 42458 7696 42460
rect 7752 42458 7776 42460
rect 7832 42458 7856 42460
rect 7912 42458 7918 42460
rect 7672 42406 7674 42458
rect 7854 42406 7856 42458
rect 7610 42404 7616 42406
rect 7672 42404 7696 42406
rect 7752 42404 7776 42406
rect 7832 42404 7856 42406
rect 7912 42404 7918 42406
rect 7610 42395 7918 42404
rect 7610 41372 7918 41381
rect 7610 41370 7616 41372
rect 7672 41370 7696 41372
rect 7752 41370 7776 41372
rect 7832 41370 7856 41372
rect 7912 41370 7918 41372
rect 7672 41318 7674 41370
rect 7854 41318 7856 41370
rect 7610 41316 7616 41318
rect 7672 41316 7696 41318
rect 7752 41316 7776 41318
rect 7832 41316 7856 41318
rect 7912 41316 7918 41318
rect 7610 41307 7918 41316
rect 7610 40284 7918 40293
rect 7610 40282 7616 40284
rect 7672 40282 7696 40284
rect 7752 40282 7776 40284
rect 7832 40282 7856 40284
rect 7912 40282 7918 40284
rect 7672 40230 7674 40282
rect 7854 40230 7856 40282
rect 7610 40228 7616 40230
rect 7672 40228 7696 40230
rect 7752 40228 7776 40230
rect 7832 40228 7856 40230
rect 7912 40228 7918 40230
rect 7610 40219 7918 40228
rect 7610 39196 7918 39205
rect 7610 39194 7616 39196
rect 7672 39194 7696 39196
rect 7752 39194 7776 39196
rect 7832 39194 7856 39196
rect 7912 39194 7918 39196
rect 7672 39142 7674 39194
rect 7854 39142 7856 39194
rect 7610 39140 7616 39142
rect 7672 39140 7696 39142
rect 7752 39140 7776 39142
rect 7832 39140 7856 39142
rect 7912 39140 7918 39142
rect 7610 39131 7918 39140
rect 7610 38108 7918 38117
rect 7610 38106 7616 38108
rect 7672 38106 7696 38108
rect 7752 38106 7776 38108
rect 7832 38106 7856 38108
rect 7912 38106 7918 38108
rect 7672 38054 7674 38106
rect 7854 38054 7856 38106
rect 7610 38052 7616 38054
rect 7672 38052 7696 38054
rect 7752 38052 7776 38054
rect 7832 38052 7856 38054
rect 7912 38052 7918 38054
rect 7610 38043 7918 38052
rect 7610 37020 7918 37029
rect 7610 37018 7616 37020
rect 7672 37018 7696 37020
rect 7752 37018 7776 37020
rect 7832 37018 7856 37020
rect 7912 37018 7918 37020
rect 7672 36966 7674 37018
rect 7854 36966 7856 37018
rect 7610 36964 7616 36966
rect 7672 36964 7696 36966
rect 7752 36964 7776 36966
rect 7832 36964 7856 36966
rect 7912 36964 7918 36966
rect 7610 36955 7918 36964
rect 7610 35932 7918 35941
rect 7610 35930 7616 35932
rect 7672 35930 7696 35932
rect 7752 35930 7776 35932
rect 7832 35930 7856 35932
rect 7912 35930 7918 35932
rect 7672 35878 7674 35930
rect 7854 35878 7856 35930
rect 7610 35876 7616 35878
rect 7672 35876 7696 35878
rect 7752 35876 7776 35878
rect 7832 35876 7856 35878
rect 7912 35876 7918 35878
rect 7610 35867 7918 35876
rect 7472 35828 7524 35834
rect 7472 35770 7524 35776
rect 7656 35828 7708 35834
rect 7656 35770 7708 35776
rect 7668 35086 7696 35770
rect 7472 35080 7524 35086
rect 7472 35022 7524 35028
rect 7656 35080 7708 35086
rect 7656 35022 7708 35028
rect 7378 34776 7434 34785
rect 7378 34711 7434 34720
rect 7484 34678 7512 35022
rect 7610 34844 7918 34853
rect 7610 34842 7616 34844
rect 7672 34842 7696 34844
rect 7752 34842 7776 34844
rect 7832 34842 7856 34844
rect 7912 34842 7918 34844
rect 7672 34790 7674 34842
rect 7854 34790 7856 34842
rect 7610 34788 7616 34790
rect 7672 34788 7696 34790
rect 7752 34788 7776 34790
rect 7832 34788 7856 34790
rect 7912 34788 7918 34790
rect 7610 34779 7918 34788
rect 7472 34672 7524 34678
rect 7472 34614 7524 34620
rect 7380 34604 7432 34610
rect 7380 34546 7432 34552
rect 7392 33658 7420 34546
rect 7470 34504 7526 34513
rect 7470 34439 7526 34448
rect 7484 34066 7512 34439
rect 7472 34060 7524 34066
rect 7472 34002 7524 34008
rect 7380 33652 7432 33658
rect 7380 33594 7432 33600
rect 7380 33448 7432 33454
rect 7380 33390 7432 33396
rect 7392 31890 7420 33390
rect 7380 31884 7432 31890
rect 7380 31826 7432 31832
rect 7484 31770 7512 34002
rect 7610 33756 7918 33765
rect 7610 33754 7616 33756
rect 7672 33754 7696 33756
rect 7752 33754 7776 33756
rect 7832 33754 7856 33756
rect 7912 33754 7918 33756
rect 7672 33702 7674 33754
rect 7854 33702 7856 33754
rect 7610 33700 7616 33702
rect 7672 33700 7696 33702
rect 7752 33700 7776 33702
rect 7832 33700 7856 33702
rect 7912 33700 7918 33702
rect 7610 33691 7918 33700
rect 7610 32668 7918 32677
rect 7610 32666 7616 32668
rect 7672 32666 7696 32668
rect 7752 32666 7776 32668
rect 7832 32666 7856 32668
rect 7912 32666 7918 32668
rect 7672 32614 7674 32666
rect 7854 32614 7856 32666
rect 7610 32612 7616 32614
rect 7672 32612 7696 32614
rect 7752 32612 7776 32614
rect 7832 32612 7856 32614
rect 7912 32612 7918 32614
rect 7610 32603 7918 32612
rect 7392 31742 7512 31770
rect 7288 24744 7340 24750
rect 7288 24686 7340 24692
rect 7288 24608 7340 24614
rect 7288 24550 7340 24556
rect 6950 24508 7258 24517
rect 6950 24506 6956 24508
rect 7012 24506 7036 24508
rect 7092 24506 7116 24508
rect 7172 24506 7196 24508
rect 7252 24506 7258 24508
rect 7012 24454 7014 24506
rect 7194 24454 7196 24506
rect 6950 24452 6956 24454
rect 7012 24452 7036 24454
rect 7092 24452 7116 24454
rect 7172 24452 7196 24454
rect 7252 24452 7258 24454
rect 6950 24443 7258 24452
rect 6950 23420 7258 23429
rect 6950 23418 6956 23420
rect 7012 23418 7036 23420
rect 7092 23418 7116 23420
rect 7172 23418 7196 23420
rect 7252 23418 7258 23420
rect 7012 23366 7014 23418
rect 7194 23366 7196 23418
rect 6950 23364 6956 23366
rect 7012 23364 7036 23366
rect 7092 23364 7116 23366
rect 7172 23364 7196 23366
rect 7252 23364 7258 23366
rect 6950 23355 7258 23364
rect 6828 23248 6880 23254
rect 6828 23190 6880 23196
rect 6840 6798 6868 23190
rect 6950 22332 7258 22341
rect 6950 22330 6956 22332
rect 7012 22330 7036 22332
rect 7092 22330 7116 22332
rect 7172 22330 7196 22332
rect 7252 22330 7258 22332
rect 7012 22278 7014 22330
rect 7194 22278 7196 22330
rect 6950 22276 6956 22278
rect 7012 22276 7036 22278
rect 7092 22276 7116 22278
rect 7172 22276 7196 22278
rect 7252 22276 7258 22278
rect 6950 22267 7258 22276
rect 6950 21244 7258 21253
rect 6950 21242 6956 21244
rect 7012 21242 7036 21244
rect 7092 21242 7116 21244
rect 7172 21242 7196 21244
rect 7252 21242 7258 21244
rect 7012 21190 7014 21242
rect 7194 21190 7196 21242
rect 6950 21188 6956 21190
rect 7012 21188 7036 21190
rect 7092 21188 7116 21190
rect 7172 21188 7196 21190
rect 7252 21188 7258 21190
rect 6950 21179 7258 21188
rect 6950 20156 7258 20165
rect 6950 20154 6956 20156
rect 7012 20154 7036 20156
rect 7092 20154 7116 20156
rect 7172 20154 7196 20156
rect 7252 20154 7258 20156
rect 7012 20102 7014 20154
rect 7194 20102 7196 20154
rect 6950 20100 6956 20102
rect 7012 20100 7036 20102
rect 7092 20100 7116 20102
rect 7172 20100 7196 20102
rect 7252 20100 7258 20102
rect 6950 20091 7258 20100
rect 7196 19712 7248 19718
rect 7196 19654 7248 19660
rect 7208 19378 7236 19654
rect 7196 19372 7248 19378
rect 7196 19314 7248 19320
rect 6950 19068 7258 19077
rect 6950 19066 6956 19068
rect 7012 19066 7036 19068
rect 7092 19066 7116 19068
rect 7172 19066 7196 19068
rect 7252 19066 7258 19068
rect 7012 19014 7014 19066
rect 7194 19014 7196 19066
rect 6950 19012 6956 19014
rect 7012 19012 7036 19014
rect 7092 19012 7116 19014
rect 7172 19012 7196 19014
rect 7252 19012 7258 19014
rect 6950 19003 7258 19012
rect 6950 17980 7258 17989
rect 6950 17978 6956 17980
rect 7012 17978 7036 17980
rect 7092 17978 7116 17980
rect 7172 17978 7196 17980
rect 7252 17978 7258 17980
rect 7012 17926 7014 17978
rect 7194 17926 7196 17978
rect 6950 17924 6956 17926
rect 7012 17924 7036 17926
rect 7092 17924 7116 17926
rect 7172 17924 7196 17926
rect 7252 17924 7258 17926
rect 6950 17915 7258 17924
rect 6950 16892 7258 16901
rect 6950 16890 6956 16892
rect 7012 16890 7036 16892
rect 7092 16890 7116 16892
rect 7172 16890 7196 16892
rect 7252 16890 7258 16892
rect 7012 16838 7014 16890
rect 7194 16838 7196 16890
rect 6950 16836 6956 16838
rect 7012 16836 7036 16838
rect 7092 16836 7116 16838
rect 7172 16836 7196 16838
rect 7252 16836 7258 16838
rect 6950 16827 7258 16836
rect 6950 15804 7258 15813
rect 6950 15802 6956 15804
rect 7012 15802 7036 15804
rect 7092 15802 7116 15804
rect 7172 15802 7196 15804
rect 7252 15802 7258 15804
rect 7012 15750 7014 15802
rect 7194 15750 7196 15802
rect 6950 15748 6956 15750
rect 7012 15748 7036 15750
rect 7092 15748 7116 15750
rect 7172 15748 7196 15750
rect 7252 15748 7258 15750
rect 6950 15739 7258 15748
rect 6950 14716 7258 14725
rect 6950 14714 6956 14716
rect 7012 14714 7036 14716
rect 7092 14714 7116 14716
rect 7172 14714 7196 14716
rect 7252 14714 7258 14716
rect 7012 14662 7014 14714
rect 7194 14662 7196 14714
rect 6950 14660 6956 14662
rect 7012 14660 7036 14662
rect 7092 14660 7116 14662
rect 7172 14660 7196 14662
rect 7252 14660 7258 14662
rect 6950 14651 7258 14660
rect 6950 13628 7258 13637
rect 6950 13626 6956 13628
rect 7012 13626 7036 13628
rect 7092 13626 7116 13628
rect 7172 13626 7196 13628
rect 7252 13626 7258 13628
rect 7012 13574 7014 13626
rect 7194 13574 7196 13626
rect 6950 13572 6956 13574
rect 7012 13572 7036 13574
rect 7092 13572 7116 13574
rect 7172 13572 7196 13574
rect 7252 13572 7258 13574
rect 6950 13563 7258 13572
rect 6950 12540 7258 12549
rect 6950 12538 6956 12540
rect 7012 12538 7036 12540
rect 7092 12538 7116 12540
rect 7172 12538 7196 12540
rect 7252 12538 7258 12540
rect 7012 12486 7014 12538
rect 7194 12486 7196 12538
rect 6950 12484 6956 12486
rect 7012 12484 7036 12486
rect 7092 12484 7116 12486
rect 7172 12484 7196 12486
rect 7252 12484 7258 12486
rect 6950 12475 7258 12484
rect 6950 11452 7258 11461
rect 6950 11450 6956 11452
rect 7012 11450 7036 11452
rect 7092 11450 7116 11452
rect 7172 11450 7196 11452
rect 7252 11450 7258 11452
rect 7012 11398 7014 11450
rect 7194 11398 7196 11450
rect 6950 11396 6956 11398
rect 7012 11396 7036 11398
rect 7092 11396 7116 11398
rect 7172 11396 7196 11398
rect 7252 11396 7258 11398
rect 6950 11387 7258 11396
rect 6950 10364 7258 10373
rect 6950 10362 6956 10364
rect 7012 10362 7036 10364
rect 7092 10362 7116 10364
rect 7172 10362 7196 10364
rect 7252 10362 7258 10364
rect 7012 10310 7014 10362
rect 7194 10310 7196 10362
rect 6950 10308 6956 10310
rect 7012 10308 7036 10310
rect 7092 10308 7116 10310
rect 7172 10308 7196 10310
rect 7252 10308 7258 10310
rect 6950 10299 7258 10308
rect 6950 9276 7258 9285
rect 6950 9274 6956 9276
rect 7012 9274 7036 9276
rect 7092 9274 7116 9276
rect 7172 9274 7196 9276
rect 7252 9274 7258 9276
rect 7012 9222 7014 9274
rect 7194 9222 7196 9274
rect 6950 9220 6956 9222
rect 7012 9220 7036 9222
rect 7092 9220 7116 9222
rect 7172 9220 7196 9222
rect 7252 9220 7258 9222
rect 6950 9211 7258 9220
rect 6950 8188 7258 8197
rect 6950 8186 6956 8188
rect 7012 8186 7036 8188
rect 7092 8186 7116 8188
rect 7172 8186 7196 8188
rect 7252 8186 7258 8188
rect 7012 8134 7014 8186
rect 7194 8134 7196 8186
rect 6950 8132 6956 8134
rect 7012 8132 7036 8134
rect 7092 8132 7116 8134
rect 7172 8132 7196 8134
rect 7252 8132 7258 8134
rect 6950 8123 7258 8132
rect 6950 7100 7258 7109
rect 6950 7098 6956 7100
rect 7012 7098 7036 7100
rect 7092 7098 7116 7100
rect 7172 7098 7196 7100
rect 7252 7098 7258 7100
rect 7012 7046 7014 7098
rect 7194 7046 7196 7098
rect 6950 7044 6956 7046
rect 7012 7044 7036 7046
rect 7092 7044 7116 7046
rect 7172 7044 7196 7046
rect 7252 7044 7258 7046
rect 6950 7035 7258 7044
rect 6828 6792 6880 6798
rect 6828 6734 6880 6740
rect 6950 6012 7258 6021
rect 6950 6010 6956 6012
rect 7012 6010 7036 6012
rect 7092 6010 7116 6012
rect 7172 6010 7196 6012
rect 7252 6010 7258 6012
rect 7012 5958 7014 6010
rect 7194 5958 7196 6010
rect 6950 5956 6956 5958
rect 7012 5956 7036 5958
rect 7092 5956 7116 5958
rect 7172 5956 7196 5958
rect 7252 5956 7258 5958
rect 6950 5947 7258 5956
rect 6748 5766 6868 5794
rect 6840 4706 6868 5766
rect 7300 5166 7328 24550
rect 7392 16590 7420 31742
rect 7472 31680 7524 31686
rect 7472 31622 7524 31628
rect 7484 25974 7512 31622
rect 7610 31580 7918 31589
rect 7610 31578 7616 31580
rect 7672 31578 7696 31580
rect 7752 31578 7776 31580
rect 7832 31578 7856 31580
rect 7912 31578 7918 31580
rect 7672 31526 7674 31578
rect 7854 31526 7856 31578
rect 7610 31524 7616 31526
rect 7672 31524 7696 31526
rect 7752 31524 7776 31526
rect 7832 31524 7856 31526
rect 7912 31524 7918 31526
rect 7610 31515 7918 31524
rect 7610 30492 7918 30501
rect 7610 30490 7616 30492
rect 7672 30490 7696 30492
rect 7752 30490 7776 30492
rect 7832 30490 7856 30492
rect 7912 30490 7918 30492
rect 7672 30438 7674 30490
rect 7854 30438 7856 30490
rect 7610 30436 7616 30438
rect 7672 30436 7696 30438
rect 7752 30436 7776 30438
rect 7832 30436 7856 30438
rect 7912 30436 7918 30438
rect 7610 30427 7918 30436
rect 7610 29404 7918 29413
rect 7610 29402 7616 29404
rect 7672 29402 7696 29404
rect 7752 29402 7776 29404
rect 7832 29402 7856 29404
rect 7912 29402 7918 29404
rect 7672 29350 7674 29402
rect 7854 29350 7856 29402
rect 7610 29348 7616 29350
rect 7672 29348 7696 29350
rect 7752 29348 7776 29350
rect 7832 29348 7856 29350
rect 7912 29348 7918 29350
rect 7610 29339 7918 29348
rect 7610 28316 7918 28325
rect 7610 28314 7616 28316
rect 7672 28314 7696 28316
rect 7752 28314 7776 28316
rect 7832 28314 7856 28316
rect 7912 28314 7918 28316
rect 7672 28262 7674 28314
rect 7854 28262 7856 28314
rect 7610 28260 7616 28262
rect 7672 28260 7696 28262
rect 7752 28260 7776 28262
rect 7832 28260 7856 28262
rect 7912 28260 7918 28262
rect 7610 28251 7918 28260
rect 7610 27228 7918 27237
rect 7610 27226 7616 27228
rect 7672 27226 7696 27228
rect 7752 27226 7776 27228
rect 7832 27226 7856 27228
rect 7912 27226 7918 27228
rect 7672 27174 7674 27226
rect 7854 27174 7856 27226
rect 7610 27172 7616 27174
rect 7672 27172 7696 27174
rect 7752 27172 7776 27174
rect 7832 27172 7856 27174
rect 7912 27172 7918 27174
rect 7610 27163 7918 27172
rect 7610 26140 7918 26149
rect 7610 26138 7616 26140
rect 7672 26138 7696 26140
rect 7752 26138 7776 26140
rect 7832 26138 7856 26140
rect 7912 26138 7918 26140
rect 7672 26086 7674 26138
rect 7854 26086 7856 26138
rect 7610 26084 7616 26086
rect 7672 26084 7696 26086
rect 7752 26084 7776 26086
rect 7832 26084 7856 26086
rect 7912 26084 7918 26086
rect 7610 26075 7918 26084
rect 7472 25968 7524 25974
rect 7472 25910 7524 25916
rect 7610 25052 7918 25061
rect 7610 25050 7616 25052
rect 7672 25050 7696 25052
rect 7752 25050 7776 25052
rect 7832 25050 7856 25052
rect 7912 25050 7918 25052
rect 7672 24998 7674 25050
rect 7854 24998 7856 25050
rect 7610 24996 7616 24998
rect 7672 24996 7696 24998
rect 7752 24996 7776 24998
rect 7832 24996 7856 24998
rect 7912 24996 7918 24998
rect 7610 24987 7918 24996
rect 8036 24818 8064 50238
rect 8128 35018 8156 60454
rect 8208 54664 8260 54670
rect 8208 54606 8260 54612
rect 8220 53514 8248 54606
rect 8208 53508 8260 53514
rect 8208 53450 8260 53456
rect 8220 52714 8248 53450
rect 8220 52686 8340 52714
rect 8208 52624 8260 52630
rect 8208 52566 8260 52572
rect 8220 51066 8248 52566
rect 8208 51060 8260 51066
rect 8208 51002 8260 51008
rect 8312 50946 8340 52686
rect 8220 50930 8340 50946
rect 8208 50924 8340 50930
rect 8260 50918 8340 50924
rect 8208 50866 8260 50872
rect 8208 50380 8260 50386
rect 8208 50322 8260 50328
rect 8220 35057 8248 50322
rect 8392 42764 8444 42770
rect 8392 42706 8444 42712
rect 8300 39976 8352 39982
rect 8300 39918 8352 39924
rect 8312 37874 8340 39918
rect 8300 37868 8352 37874
rect 8300 37810 8352 37816
rect 8312 35850 8340 37810
rect 8404 37398 8432 42706
rect 8496 41546 8524 60658
rect 8852 60512 8904 60518
rect 8852 60454 8904 60460
rect 8484 41540 8536 41546
rect 8484 41482 8536 41488
rect 8760 41472 8812 41478
rect 8760 41414 8812 41420
rect 8392 37392 8444 37398
rect 8392 37334 8444 37340
rect 8312 35822 8432 35850
rect 8206 35048 8262 35057
rect 8116 35012 8168 35018
rect 8206 34983 8262 34992
rect 8116 34954 8168 34960
rect 8128 34898 8156 34954
rect 8128 34870 8340 34898
rect 8206 34776 8262 34785
rect 8206 34711 8262 34720
rect 8116 34672 8168 34678
rect 8116 34614 8168 34620
rect 8024 24812 8076 24818
rect 8024 24754 8076 24760
rect 7472 24744 7524 24750
rect 7472 24686 7524 24692
rect 7484 24206 7512 24686
rect 8036 24290 8064 24754
rect 8128 24410 8156 34614
rect 8116 24404 8168 24410
rect 8116 24346 8168 24352
rect 8036 24262 8156 24290
rect 7472 24200 7524 24206
rect 7472 24142 7524 24148
rect 7484 23798 7512 24142
rect 8024 24132 8076 24138
rect 8024 24074 8076 24080
rect 7610 23964 7918 23973
rect 7610 23962 7616 23964
rect 7672 23962 7696 23964
rect 7752 23962 7776 23964
rect 7832 23962 7856 23964
rect 7912 23962 7918 23964
rect 7672 23910 7674 23962
rect 7854 23910 7856 23962
rect 7610 23908 7616 23910
rect 7672 23908 7696 23910
rect 7752 23908 7776 23910
rect 7832 23908 7856 23910
rect 7912 23908 7918 23910
rect 7610 23899 7918 23908
rect 7472 23792 7524 23798
rect 7472 23734 7524 23740
rect 7610 22876 7918 22885
rect 7610 22874 7616 22876
rect 7672 22874 7696 22876
rect 7752 22874 7776 22876
rect 7832 22874 7856 22876
rect 7912 22874 7918 22876
rect 7672 22822 7674 22874
rect 7854 22822 7856 22874
rect 7610 22820 7616 22822
rect 7672 22820 7696 22822
rect 7752 22820 7776 22822
rect 7832 22820 7856 22822
rect 7912 22820 7918 22822
rect 7610 22811 7918 22820
rect 7472 22500 7524 22506
rect 7472 22442 7524 22448
rect 7484 18426 7512 22442
rect 7610 21788 7918 21797
rect 7610 21786 7616 21788
rect 7672 21786 7696 21788
rect 7752 21786 7776 21788
rect 7832 21786 7856 21788
rect 7912 21786 7918 21788
rect 7672 21734 7674 21786
rect 7854 21734 7856 21786
rect 7610 21732 7616 21734
rect 7672 21732 7696 21734
rect 7752 21732 7776 21734
rect 7832 21732 7856 21734
rect 7912 21732 7918 21734
rect 7610 21723 7918 21732
rect 7840 21344 7892 21350
rect 7840 21286 7892 21292
rect 7852 20942 7880 21286
rect 7840 20936 7892 20942
rect 7840 20878 7892 20884
rect 7610 20700 7918 20709
rect 7610 20698 7616 20700
rect 7672 20698 7696 20700
rect 7752 20698 7776 20700
rect 7832 20698 7856 20700
rect 7912 20698 7918 20700
rect 7672 20646 7674 20698
rect 7854 20646 7856 20698
rect 7610 20644 7616 20646
rect 7672 20644 7696 20646
rect 7752 20644 7776 20646
rect 7832 20644 7856 20646
rect 7912 20644 7918 20646
rect 7610 20635 7918 20644
rect 8036 19922 8064 24074
rect 8128 23798 8156 24262
rect 8116 23792 8168 23798
rect 8116 23734 8168 23740
rect 8024 19916 8076 19922
rect 8024 19858 8076 19864
rect 7610 19612 7918 19621
rect 7610 19610 7616 19612
rect 7672 19610 7696 19612
rect 7752 19610 7776 19612
rect 7832 19610 7856 19612
rect 7912 19610 7918 19612
rect 7672 19558 7674 19610
rect 7854 19558 7856 19610
rect 7610 19556 7616 19558
rect 7672 19556 7696 19558
rect 7752 19556 7776 19558
rect 7832 19556 7856 19558
rect 7912 19556 7918 19558
rect 7610 19547 7918 19556
rect 8036 19446 8064 19858
rect 8116 19712 8168 19718
rect 8116 19654 8168 19660
rect 8024 19440 8076 19446
rect 8024 19382 8076 19388
rect 8024 19304 8076 19310
rect 8024 19246 8076 19252
rect 7610 18524 7918 18533
rect 7610 18522 7616 18524
rect 7672 18522 7696 18524
rect 7752 18522 7776 18524
rect 7832 18522 7856 18524
rect 7912 18522 7918 18524
rect 7672 18470 7674 18522
rect 7854 18470 7856 18522
rect 7610 18468 7616 18470
rect 7672 18468 7696 18470
rect 7752 18468 7776 18470
rect 7832 18468 7856 18470
rect 7912 18468 7918 18470
rect 7610 18459 7918 18468
rect 7472 18420 7524 18426
rect 7472 18362 7524 18368
rect 7610 17436 7918 17445
rect 7610 17434 7616 17436
rect 7672 17434 7696 17436
rect 7752 17434 7776 17436
rect 7832 17434 7856 17436
rect 7912 17434 7918 17436
rect 7672 17382 7674 17434
rect 7854 17382 7856 17434
rect 7610 17380 7616 17382
rect 7672 17380 7696 17382
rect 7752 17380 7776 17382
rect 7832 17380 7856 17382
rect 7912 17380 7918 17382
rect 7610 17371 7918 17380
rect 7472 17264 7524 17270
rect 7472 17206 7524 17212
rect 7380 16584 7432 16590
rect 7380 16526 7432 16532
rect 7380 13184 7432 13190
rect 7380 13126 7432 13132
rect 7288 5160 7340 5166
rect 7288 5102 7340 5108
rect 6950 4924 7258 4933
rect 6950 4922 6956 4924
rect 7012 4922 7036 4924
rect 7092 4922 7116 4924
rect 7172 4922 7196 4924
rect 7252 4922 7258 4924
rect 7012 4870 7014 4922
rect 7194 4870 7196 4922
rect 6950 4868 6956 4870
rect 7012 4868 7036 4870
rect 7092 4868 7116 4870
rect 7172 4868 7196 4870
rect 7252 4868 7258 4870
rect 6950 4859 7258 4868
rect 6840 4678 7052 4706
rect 7024 4622 7052 4678
rect 7012 4616 7064 4622
rect 7012 4558 7064 4564
rect 7300 4486 7328 5102
rect 7392 4826 7420 13126
rect 7380 4820 7432 4826
rect 7380 4762 7432 4768
rect 7484 4690 7512 17206
rect 7610 16348 7918 16357
rect 7610 16346 7616 16348
rect 7672 16346 7696 16348
rect 7752 16346 7776 16348
rect 7832 16346 7856 16348
rect 7912 16346 7918 16348
rect 7672 16294 7674 16346
rect 7854 16294 7856 16346
rect 7610 16292 7616 16294
rect 7672 16292 7696 16294
rect 7752 16292 7776 16294
rect 7832 16292 7856 16294
rect 7912 16292 7918 16294
rect 7610 16283 7918 16292
rect 7610 15260 7918 15269
rect 7610 15258 7616 15260
rect 7672 15258 7696 15260
rect 7752 15258 7776 15260
rect 7832 15258 7856 15260
rect 7912 15258 7918 15260
rect 7672 15206 7674 15258
rect 7854 15206 7856 15258
rect 7610 15204 7616 15206
rect 7672 15204 7696 15206
rect 7752 15204 7776 15206
rect 7832 15204 7856 15206
rect 7912 15204 7918 15206
rect 7610 15195 7918 15204
rect 7610 14172 7918 14181
rect 7610 14170 7616 14172
rect 7672 14170 7696 14172
rect 7752 14170 7776 14172
rect 7832 14170 7856 14172
rect 7912 14170 7918 14172
rect 7672 14118 7674 14170
rect 7854 14118 7856 14170
rect 7610 14116 7616 14118
rect 7672 14116 7696 14118
rect 7752 14116 7776 14118
rect 7832 14116 7856 14118
rect 7912 14116 7918 14118
rect 7610 14107 7918 14116
rect 7610 13084 7918 13093
rect 7610 13082 7616 13084
rect 7672 13082 7696 13084
rect 7752 13082 7776 13084
rect 7832 13082 7856 13084
rect 7912 13082 7918 13084
rect 7672 13030 7674 13082
rect 7854 13030 7856 13082
rect 7610 13028 7616 13030
rect 7672 13028 7696 13030
rect 7752 13028 7776 13030
rect 7832 13028 7856 13030
rect 7912 13028 7918 13030
rect 7610 13019 7918 13028
rect 7610 11996 7918 12005
rect 7610 11994 7616 11996
rect 7672 11994 7696 11996
rect 7752 11994 7776 11996
rect 7832 11994 7856 11996
rect 7912 11994 7918 11996
rect 7672 11942 7674 11994
rect 7854 11942 7856 11994
rect 7610 11940 7616 11942
rect 7672 11940 7696 11942
rect 7752 11940 7776 11942
rect 7832 11940 7856 11942
rect 7912 11940 7918 11942
rect 7610 11931 7918 11940
rect 7610 10908 7918 10917
rect 7610 10906 7616 10908
rect 7672 10906 7696 10908
rect 7752 10906 7776 10908
rect 7832 10906 7856 10908
rect 7912 10906 7918 10908
rect 7672 10854 7674 10906
rect 7854 10854 7856 10906
rect 7610 10852 7616 10854
rect 7672 10852 7696 10854
rect 7752 10852 7776 10854
rect 7832 10852 7856 10854
rect 7912 10852 7918 10854
rect 7610 10843 7918 10852
rect 7610 9820 7918 9829
rect 7610 9818 7616 9820
rect 7672 9818 7696 9820
rect 7752 9818 7776 9820
rect 7832 9818 7856 9820
rect 7912 9818 7918 9820
rect 7672 9766 7674 9818
rect 7854 9766 7856 9818
rect 7610 9764 7616 9766
rect 7672 9764 7696 9766
rect 7752 9764 7776 9766
rect 7832 9764 7856 9766
rect 7912 9764 7918 9766
rect 7610 9755 7918 9764
rect 7610 8732 7918 8741
rect 7610 8730 7616 8732
rect 7672 8730 7696 8732
rect 7752 8730 7776 8732
rect 7832 8730 7856 8732
rect 7912 8730 7918 8732
rect 7672 8678 7674 8730
rect 7854 8678 7856 8730
rect 7610 8676 7616 8678
rect 7672 8676 7696 8678
rect 7752 8676 7776 8678
rect 7832 8676 7856 8678
rect 7912 8676 7918 8678
rect 7610 8667 7918 8676
rect 7610 7644 7918 7653
rect 7610 7642 7616 7644
rect 7672 7642 7696 7644
rect 7752 7642 7776 7644
rect 7832 7642 7856 7644
rect 7912 7642 7918 7644
rect 7672 7590 7674 7642
rect 7854 7590 7856 7642
rect 7610 7588 7616 7590
rect 7672 7588 7696 7590
rect 7752 7588 7776 7590
rect 7832 7588 7856 7590
rect 7912 7588 7918 7590
rect 7610 7579 7918 7588
rect 7610 6556 7918 6565
rect 7610 6554 7616 6556
rect 7672 6554 7696 6556
rect 7752 6554 7776 6556
rect 7832 6554 7856 6556
rect 7912 6554 7918 6556
rect 7672 6502 7674 6554
rect 7854 6502 7856 6554
rect 7610 6500 7616 6502
rect 7672 6500 7696 6502
rect 7752 6500 7776 6502
rect 7832 6500 7856 6502
rect 7912 6500 7918 6502
rect 7610 6491 7918 6500
rect 7610 5468 7918 5477
rect 7610 5466 7616 5468
rect 7672 5466 7696 5468
rect 7752 5466 7776 5468
rect 7832 5466 7856 5468
rect 7912 5466 7918 5468
rect 7672 5414 7674 5466
rect 7854 5414 7856 5466
rect 7610 5412 7616 5414
rect 7672 5412 7696 5414
rect 7752 5412 7776 5414
rect 7832 5412 7856 5414
rect 7912 5412 7918 5414
rect 7610 5403 7918 5412
rect 7472 4684 7524 4690
rect 7472 4626 7524 4632
rect 7288 4480 7340 4486
rect 7288 4422 7340 4428
rect 7610 4380 7918 4389
rect 7610 4378 7616 4380
rect 7672 4378 7696 4380
rect 7752 4378 7776 4380
rect 7832 4378 7856 4380
rect 7912 4378 7918 4380
rect 7672 4326 7674 4378
rect 7854 4326 7856 4378
rect 7610 4324 7616 4326
rect 7672 4324 7696 4326
rect 7752 4324 7776 4326
rect 7832 4324 7856 4326
rect 7912 4324 7918 4326
rect 7610 4315 7918 4324
rect 6460 4140 6512 4146
rect 6460 4082 6512 4088
rect 6950 3836 7258 3845
rect 6950 3834 6956 3836
rect 7012 3834 7036 3836
rect 7092 3834 7116 3836
rect 7172 3834 7196 3836
rect 7252 3834 7258 3836
rect 7012 3782 7014 3834
rect 7194 3782 7196 3834
rect 6950 3780 6956 3782
rect 7012 3780 7036 3782
rect 7092 3780 7116 3782
rect 7172 3780 7196 3782
rect 7252 3780 7258 3782
rect 6950 3771 7258 3780
rect 4804 3528 4856 3534
rect 4804 3470 4856 3476
rect 8036 3466 8064 19246
rect 8128 18578 8156 19654
rect 8220 19310 8248 34711
rect 8312 31210 8340 34870
rect 8404 33454 8432 35822
rect 8392 33448 8444 33454
rect 8392 33390 8444 33396
rect 8300 31204 8352 31210
rect 8300 31146 8352 31152
rect 8668 29504 8720 29510
rect 8668 29446 8720 29452
rect 8392 25968 8444 25974
rect 8392 25910 8444 25916
rect 8300 24404 8352 24410
rect 8300 24346 8352 24352
rect 8312 23866 8340 24346
rect 8300 23860 8352 23866
rect 8300 23802 8352 23808
rect 8312 23662 8340 23802
rect 8300 23656 8352 23662
rect 8300 23598 8352 23604
rect 8404 22506 8432 25910
rect 8484 23520 8536 23526
rect 8484 23462 8536 23468
rect 8392 22500 8444 22506
rect 8392 22442 8444 22448
rect 8208 19304 8260 19310
rect 8208 19246 8260 19252
rect 8128 18550 8248 18578
rect 8116 18420 8168 18426
rect 8116 18362 8168 18368
rect 8128 5030 8156 18362
rect 8220 10538 8248 18550
rect 8208 10532 8260 10538
rect 8208 10474 8260 10480
rect 8208 9104 8260 9110
rect 8208 9046 8260 9052
rect 8220 5234 8248 9046
rect 8392 5296 8444 5302
rect 8392 5238 8444 5244
rect 8208 5228 8260 5234
rect 8208 5170 8260 5176
rect 8116 5024 8168 5030
rect 8116 4966 8168 4972
rect 8404 4758 8432 5238
rect 8496 5234 8524 23462
rect 8680 22982 8708 29446
rect 8668 22976 8720 22982
rect 8668 22918 8720 22924
rect 8680 22710 8708 22918
rect 8668 22704 8720 22710
rect 8668 22646 8720 22652
rect 8484 5228 8536 5234
rect 8484 5170 8536 5176
rect 8392 4752 8444 4758
rect 8392 4694 8444 4700
rect 8208 4616 8260 4622
rect 8208 4558 8260 4564
rect 8024 3460 8076 3466
rect 8024 3402 8076 3408
rect 8220 3398 8248 4558
rect 8208 3392 8260 3398
rect 8208 3334 8260 3340
rect 2610 3292 2918 3301
rect 2610 3290 2616 3292
rect 2672 3290 2696 3292
rect 2752 3290 2776 3292
rect 2832 3290 2856 3292
rect 2912 3290 2918 3292
rect 2672 3238 2674 3290
rect 2854 3238 2856 3290
rect 2610 3236 2616 3238
rect 2672 3236 2696 3238
rect 2752 3236 2776 3238
rect 2832 3236 2856 3238
rect 2912 3236 2918 3238
rect 2610 3227 2918 3236
rect 7610 3292 7918 3301
rect 7610 3290 7616 3292
rect 7672 3290 7696 3292
rect 7752 3290 7776 3292
rect 7832 3290 7856 3292
rect 7912 3290 7918 3292
rect 7672 3238 7674 3290
rect 7854 3238 7856 3290
rect 7610 3236 7616 3238
rect 7672 3236 7696 3238
rect 7752 3236 7776 3238
rect 7832 3236 7856 3238
rect 7912 3236 7918 3238
rect 7610 3227 7918 3236
rect 8496 3194 8524 5170
rect 8772 5098 8800 41414
rect 8864 30190 8892 60454
rect 8956 50318 8984 61134
rect 9036 60716 9088 60722
rect 9036 60658 9088 60664
rect 9048 56982 9076 60658
rect 9036 56976 9088 56982
rect 9036 56918 9088 56924
rect 8944 50312 8996 50318
rect 8944 50254 8996 50260
rect 8956 49774 8984 50254
rect 8944 49768 8996 49774
rect 8944 49710 8996 49716
rect 8944 48680 8996 48686
rect 8944 48622 8996 48628
rect 8956 45490 8984 48622
rect 8944 45484 8996 45490
rect 8944 45426 8996 45432
rect 9048 45422 9076 56918
rect 9232 50454 9260 61134
rect 9404 55820 9456 55826
rect 9404 55762 9456 55768
rect 9312 54596 9364 54602
rect 9312 54538 9364 54544
rect 9324 53650 9352 54538
rect 9312 53644 9364 53650
rect 9312 53586 9364 53592
rect 9220 50448 9272 50454
rect 9220 50390 9272 50396
rect 9416 45554 9444 55762
rect 9496 55752 9548 55758
rect 9496 55694 9548 55700
rect 9232 45526 9444 45554
rect 9036 45416 9088 45422
rect 9036 45358 9088 45364
rect 9048 44198 9076 45358
rect 9232 44402 9260 45526
rect 9220 44396 9272 44402
rect 9220 44338 9272 44344
rect 9036 44192 9088 44198
rect 9036 44134 9088 44140
rect 9128 41812 9180 41818
rect 9128 41754 9180 41760
rect 8944 41744 8996 41750
rect 8944 41686 8996 41692
rect 8956 41546 8984 41686
rect 8944 41540 8996 41546
rect 8944 41482 8996 41488
rect 8852 30184 8904 30190
rect 8852 30126 8904 30132
rect 8864 29322 8892 30126
rect 8956 29510 8984 41482
rect 9036 31816 9088 31822
rect 9036 31758 9088 31764
rect 8944 29504 8996 29510
rect 8944 29446 8996 29452
rect 8864 29294 8984 29322
rect 8852 29164 8904 29170
rect 8852 29106 8904 29112
rect 8760 5092 8812 5098
rect 8760 5034 8812 5040
rect 8864 4078 8892 29106
rect 8956 23254 8984 29294
rect 9048 25906 9076 31758
rect 9140 30326 9168 41754
rect 9128 30320 9180 30326
rect 9128 30262 9180 30268
rect 9232 29850 9260 44338
rect 9508 44266 9536 55694
rect 9496 44260 9548 44266
rect 9496 44202 9548 44208
rect 9312 44192 9364 44198
rect 9312 44134 9364 44140
rect 9324 31890 9352 44134
rect 9404 43104 9456 43110
rect 9404 43046 9456 43052
rect 9312 31884 9364 31890
rect 9312 31826 9364 31832
rect 9220 29844 9272 29850
rect 9220 29786 9272 29792
rect 9128 28960 9180 28966
rect 9128 28902 9180 28908
rect 9036 25900 9088 25906
rect 9036 25842 9088 25848
rect 8944 23248 8996 23254
rect 8944 23190 8996 23196
rect 8944 22976 8996 22982
rect 8944 22918 8996 22924
rect 8956 7546 8984 22918
rect 9048 22166 9076 25842
rect 9036 22160 9088 22166
rect 9036 22102 9088 22108
rect 9140 14618 9168 28902
rect 9312 20868 9364 20874
rect 9312 20810 9364 20816
rect 9220 16108 9272 16114
rect 9220 16050 9272 16056
rect 9128 14612 9180 14618
rect 9128 14554 9180 14560
rect 8944 7540 8996 7546
rect 8944 7482 8996 7488
rect 9232 4146 9260 16050
rect 9324 10470 9352 20810
rect 9416 16046 9444 43046
rect 9508 41818 9536 44202
rect 9600 43314 9628 62630
rect 10324 61124 10376 61130
rect 10324 61066 10376 61072
rect 10140 56908 10192 56914
rect 10140 56850 10192 56856
rect 9956 55752 10008 55758
rect 9956 55694 10008 55700
rect 9680 47728 9732 47734
rect 9680 47670 9732 47676
rect 9692 43314 9720 47670
rect 9968 44334 9996 55694
rect 9956 44328 10008 44334
rect 9956 44270 10008 44276
rect 9968 44198 9996 44270
rect 9956 44192 10008 44198
rect 9956 44134 10008 44140
rect 9588 43308 9640 43314
rect 9588 43250 9640 43256
rect 9680 43308 9732 43314
rect 9680 43250 9732 43256
rect 10048 43308 10100 43314
rect 10048 43250 10100 43256
rect 9496 41812 9548 41818
rect 9496 41754 9548 41760
rect 9864 39092 9916 39098
rect 9864 39034 9916 39040
rect 9588 36168 9640 36174
rect 9588 36110 9640 36116
rect 9494 31240 9550 31249
rect 9494 31175 9550 31184
rect 9508 19378 9536 31175
rect 9600 26450 9628 36110
rect 9772 35760 9824 35766
rect 9772 35702 9824 35708
rect 9784 35290 9812 35702
rect 9772 35284 9824 35290
rect 9772 35226 9824 35232
rect 9876 35086 9904 39034
rect 9772 35080 9824 35086
rect 9772 35022 9824 35028
rect 9864 35080 9916 35086
rect 9864 35022 9916 35028
rect 9784 32570 9812 35022
rect 9772 32564 9824 32570
rect 9772 32506 9824 32512
rect 9876 30734 9904 35022
rect 9864 30728 9916 30734
rect 9864 30670 9916 30676
rect 10060 28966 10088 43250
rect 9680 28960 9732 28966
rect 9680 28902 9732 28908
rect 10048 28960 10100 28966
rect 10048 28902 10100 28908
rect 9588 26444 9640 26450
rect 9588 26386 9640 26392
rect 9692 26314 9720 28902
rect 9680 26308 9732 26314
rect 9680 26250 9732 26256
rect 9496 19372 9548 19378
rect 9496 19314 9548 19320
rect 9404 16040 9456 16046
rect 9404 15982 9456 15988
rect 9312 10464 9364 10470
rect 9312 10406 9364 10412
rect 9220 4140 9272 4146
rect 9220 4082 9272 4088
rect 8852 4072 8904 4078
rect 8852 4014 8904 4020
rect 8484 3188 8536 3194
rect 8484 3130 8536 3136
rect 6950 2748 7258 2757
rect 6950 2746 6956 2748
rect 7012 2746 7036 2748
rect 7092 2746 7116 2748
rect 7172 2746 7196 2748
rect 7252 2746 7258 2748
rect 7012 2694 7014 2746
rect 7194 2694 7196 2746
rect 6950 2692 6956 2694
rect 7012 2692 7036 2694
rect 7092 2692 7116 2694
rect 7172 2692 7196 2694
rect 7252 2692 7258 2694
rect 6950 2683 7258 2692
rect 2504 2508 2556 2514
rect 2504 2450 2556 2456
rect 2320 2304 2372 2310
rect 2320 2246 2372 2252
rect 2516 1170 2544 2450
rect 10152 2446 10180 56850
rect 10336 46442 10364 61066
rect 10324 46436 10376 46442
rect 10324 46378 10376 46384
rect 10428 45014 10456 66574
rect 10520 48278 10548 67050
rect 10876 62892 10928 62898
rect 10876 62834 10928 62840
rect 10692 60784 10744 60790
rect 10692 60726 10744 60732
rect 10704 56914 10732 60726
rect 10692 56908 10744 56914
rect 10692 56850 10744 56856
rect 10784 56840 10836 56846
rect 10782 56808 10784 56817
rect 10836 56808 10838 56817
rect 10782 56743 10838 56752
rect 10692 55956 10744 55962
rect 10692 55898 10744 55904
rect 10704 50930 10732 55898
rect 10888 55214 10916 62834
rect 10968 57928 11020 57934
rect 10968 57870 11020 57876
rect 10980 55894 11008 57870
rect 10968 55888 11020 55894
rect 10968 55830 11020 55836
rect 10888 55186 11008 55214
rect 10876 52080 10928 52086
rect 10876 52022 10928 52028
rect 10784 51876 10836 51882
rect 10784 51818 10836 51824
rect 10692 50924 10744 50930
rect 10692 50866 10744 50872
rect 10796 50810 10824 51818
rect 10888 50930 10916 52022
rect 10876 50924 10928 50930
rect 10876 50866 10928 50872
rect 10796 50782 10916 50810
rect 10600 50448 10652 50454
rect 10600 50390 10652 50396
rect 10508 48272 10560 48278
rect 10508 48214 10560 48220
rect 10416 45008 10468 45014
rect 10416 44950 10468 44956
rect 10232 44260 10284 44266
rect 10232 44202 10284 44208
rect 10244 38758 10272 44202
rect 10508 43240 10560 43246
rect 10508 43182 10560 43188
rect 10416 41064 10468 41070
rect 10416 41006 10468 41012
rect 10428 39914 10456 41006
rect 10416 39908 10468 39914
rect 10416 39850 10468 39856
rect 10232 38752 10284 38758
rect 10232 38694 10284 38700
rect 10324 38208 10376 38214
rect 10324 38150 10376 38156
rect 10232 35828 10284 35834
rect 10232 35770 10284 35776
rect 10244 35086 10272 35770
rect 10232 35080 10284 35086
rect 10232 35022 10284 35028
rect 10244 33114 10272 35022
rect 10232 33108 10284 33114
rect 10232 33050 10284 33056
rect 10232 31884 10284 31890
rect 10232 31826 10284 31832
rect 10244 31278 10272 31826
rect 10232 31272 10284 31278
rect 10232 31214 10284 31220
rect 10336 23186 10364 38150
rect 10428 24682 10456 39850
rect 10520 35290 10548 43182
rect 10612 40934 10640 50390
rect 10692 48612 10744 48618
rect 10692 48554 10744 48560
rect 10600 40928 10652 40934
rect 10600 40870 10652 40876
rect 10612 40118 10640 40870
rect 10600 40112 10652 40118
rect 10600 40054 10652 40060
rect 10508 35284 10560 35290
rect 10508 35226 10560 35232
rect 10600 29096 10652 29102
rect 10600 29038 10652 29044
rect 10508 24812 10560 24818
rect 10508 24754 10560 24760
rect 10416 24676 10468 24682
rect 10416 24618 10468 24624
rect 10520 24410 10548 24754
rect 10508 24404 10560 24410
rect 10508 24346 10560 24352
rect 10324 23180 10376 23186
rect 10324 23122 10376 23128
rect 10612 21010 10640 29038
rect 10704 28490 10732 48554
rect 10784 46368 10836 46374
rect 10784 46310 10836 46316
rect 10796 28558 10824 46310
rect 10888 43450 10916 50782
rect 10876 43444 10928 43450
rect 10876 43386 10928 43392
rect 10980 40662 11008 55186
rect 11244 52012 11296 52018
rect 11244 51954 11296 51960
rect 11152 49768 11204 49774
rect 11152 49710 11204 49716
rect 10968 40656 11020 40662
rect 10968 40598 11020 40604
rect 10876 40112 10928 40118
rect 10876 40054 10928 40060
rect 10784 28552 10836 28558
rect 10784 28494 10836 28500
rect 10692 28484 10744 28490
rect 10692 28426 10744 28432
rect 10704 25294 10732 28426
rect 10692 25288 10744 25294
rect 10692 25230 10744 25236
rect 10600 21004 10652 21010
rect 10600 20946 10652 20952
rect 10888 3602 10916 40054
rect 10980 36242 11008 40598
rect 11060 37936 11112 37942
rect 11060 37878 11112 37884
rect 10968 36236 11020 36242
rect 10968 36178 11020 36184
rect 11072 35154 11100 37878
rect 11060 35148 11112 35154
rect 11060 35090 11112 35096
rect 11060 25832 11112 25838
rect 11060 25774 11112 25780
rect 10968 24268 11020 24274
rect 10968 24210 11020 24216
rect 10980 18834 11008 24210
rect 11072 22710 11100 25774
rect 11060 22704 11112 22710
rect 11060 22646 11112 22652
rect 10968 18828 11020 18834
rect 10968 18770 11020 18776
rect 10968 10736 11020 10742
rect 10968 10678 11020 10684
rect 10980 3670 11008 10678
rect 10968 3664 11020 3670
rect 10968 3606 11020 3612
rect 10876 3596 10928 3602
rect 10876 3538 10928 3544
rect 11164 3534 11192 49710
rect 11256 43246 11284 51954
rect 11440 50862 11468 68750
rect 11520 68740 11572 68746
rect 11520 68682 11572 68688
rect 11428 50856 11480 50862
rect 11428 50798 11480 50804
rect 11440 48754 11468 50798
rect 11428 48748 11480 48754
rect 11428 48690 11480 48696
rect 11440 48550 11468 48690
rect 11532 48686 11560 68682
rect 12610 68572 12918 68581
rect 12610 68570 12616 68572
rect 12672 68570 12696 68572
rect 12752 68570 12776 68572
rect 12832 68570 12856 68572
rect 12912 68570 12918 68572
rect 12672 68518 12674 68570
rect 12854 68518 12856 68570
rect 12610 68516 12616 68518
rect 12672 68516 12696 68518
rect 12752 68516 12776 68518
rect 12832 68516 12856 68518
rect 12912 68516 12918 68518
rect 12610 68507 12918 68516
rect 11950 68028 12258 68037
rect 11950 68026 11956 68028
rect 12012 68026 12036 68028
rect 12092 68026 12116 68028
rect 12172 68026 12196 68028
rect 12252 68026 12258 68028
rect 12012 67974 12014 68026
rect 12194 67974 12196 68026
rect 11950 67972 11956 67974
rect 12012 67972 12036 67974
rect 12092 67972 12116 67974
rect 12172 67972 12196 67974
rect 12252 67972 12258 67974
rect 11950 67963 12258 67972
rect 13084 67720 13136 67726
rect 13084 67662 13136 67668
rect 12992 67652 13044 67658
rect 12992 67594 13044 67600
rect 12610 67484 12918 67493
rect 12610 67482 12616 67484
rect 12672 67482 12696 67484
rect 12752 67482 12776 67484
rect 12832 67482 12856 67484
rect 12912 67482 12918 67484
rect 12672 67430 12674 67482
rect 12854 67430 12856 67482
rect 12610 67428 12616 67430
rect 12672 67428 12696 67430
rect 12752 67428 12776 67430
rect 12832 67428 12856 67430
rect 12912 67428 12918 67430
rect 12610 67419 12918 67428
rect 11950 66940 12258 66949
rect 11950 66938 11956 66940
rect 12012 66938 12036 66940
rect 12092 66938 12116 66940
rect 12172 66938 12196 66940
rect 12252 66938 12258 66940
rect 12012 66886 12014 66938
rect 12194 66886 12196 66938
rect 11950 66884 11956 66886
rect 12012 66884 12036 66886
rect 12092 66884 12116 66886
rect 12172 66884 12196 66886
rect 12252 66884 12258 66886
rect 11950 66875 12258 66884
rect 12610 66396 12918 66405
rect 12610 66394 12616 66396
rect 12672 66394 12696 66396
rect 12752 66394 12776 66396
rect 12832 66394 12856 66396
rect 12912 66394 12918 66396
rect 12672 66342 12674 66394
rect 12854 66342 12856 66394
rect 12610 66340 12616 66342
rect 12672 66340 12696 66342
rect 12752 66340 12776 66342
rect 12832 66340 12856 66342
rect 12912 66340 12918 66342
rect 12610 66331 12918 66340
rect 11950 65852 12258 65861
rect 11950 65850 11956 65852
rect 12012 65850 12036 65852
rect 12092 65850 12116 65852
rect 12172 65850 12196 65852
rect 12252 65850 12258 65852
rect 12012 65798 12014 65850
rect 12194 65798 12196 65850
rect 11950 65796 11956 65798
rect 12012 65796 12036 65798
rect 12092 65796 12116 65798
rect 12172 65796 12196 65798
rect 12252 65796 12258 65798
rect 11950 65787 12258 65796
rect 11888 65544 11940 65550
rect 11888 65486 11940 65492
rect 11900 65210 11928 65486
rect 12348 65476 12400 65482
rect 12348 65418 12400 65424
rect 11888 65204 11940 65210
rect 11888 65146 11940 65152
rect 11950 64764 12258 64773
rect 11950 64762 11956 64764
rect 12012 64762 12036 64764
rect 12092 64762 12116 64764
rect 12172 64762 12196 64764
rect 12252 64762 12258 64764
rect 12012 64710 12014 64762
rect 12194 64710 12196 64762
rect 11950 64708 11956 64710
rect 12012 64708 12036 64710
rect 12092 64708 12116 64710
rect 12172 64708 12196 64710
rect 12252 64708 12258 64710
rect 11950 64699 12258 64708
rect 11950 63676 12258 63685
rect 11950 63674 11956 63676
rect 12012 63674 12036 63676
rect 12092 63674 12116 63676
rect 12172 63674 12196 63676
rect 12252 63674 12258 63676
rect 12012 63622 12014 63674
rect 12194 63622 12196 63674
rect 11950 63620 11956 63622
rect 12012 63620 12036 63622
rect 12092 63620 12116 63622
rect 12172 63620 12196 63622
rect 12252 63620 12258 63622
rect 11950 63611 12258 63620
rect 11950 62588 12258 62597
rect 11950 62586 11956 62588
rect 12012 62586 12036 62588
rect 12092 62586 12116 62588
rect 12172 62586 12196 62588
rect 12252 62586 12258 62588
rect 12012 62534 12014 62586
rect 12194 62534 12196 62586
rect 11950 62532 11956 62534
rect 12012 62532 12036 62534
rect 12092 62532 12116 62534
rect 12172 62532 12196 62534
rect 12252 62532 12258 62534
rect 11950 62523 12258 62532
rect 11796 61736 11848 61742
rect 11796 61678 11848 61684
rect 11704 55752 11756 55758
rect 11704 55694 11756 55700
rect 11612 50992 11664 50998
rect 11612 50934 11664 50940
rect 11624 50250 11652 50934
rect 11612 50244 11664 50250
rect 11612 50186 11664 50192
rect 11520 48680 11572 48686
rect 11520 48622 11572 48628
rect 11428 48544 11480 48550
rect 11428 48486 11480 48492
rect 11336 48272 11388 48278
rect 11336 48214 11388 48220
rect 11244 43240 11296 43246
rect 11244 43182 11296 43188
rect 11348 30122 11376 48214
rect 11428 43240 11480 43246
rect 11428 43182 11480 43188
rect 11440 32502 11468 43182
rect 11520 33040 11572 33046
rect 11520 32982 11572 32988
rect 11428 32496 11480 32502
rect 11428 32438 11480 32444
rect 11336 30116 11388 30122
rect 11336 30058 11388 30064
rect 11348 29102 11376 30058
rect 11336 29096 11388 29102
rect 11336 29038 11388 29044
rect 11532 29034 11560 32982
rect 11624 32978 11652 50186
rect 11716 36378 11744 55694
rect 11808 41478 11836 61678
rect 11950 61500 12258 61509
rect 11950 61498 11956 61500
rect 12012 61498 12036 61500
rect 12092 61498 12116 61500
rect 12172 61498 12196 61500
rect 12252 61498 12258 61500
rect 12012 61446 12014 61498
rect 12194 61446 12196 61498
rect 11950 61444 11956 61446
rect 12012 61444 12036 61446
rect 12092 61444 12116 61446
rect 12172 61444 12196 61446
rect 12252 61444 12258 61446
rect 11950 61435 12258 61444
rect 11950 60412 12258 60421
rect 11950 60410 11956 60412
rect 12012 60410 12036 60412
rect 12092 60410 12116 60412
rect 12172 60410 12196 60412
rect 12252 60410 12258 60412
rect 12012 60358 12014 60410
rect 12194 60358 12196 60410
rect 11950 60356 11956 60358
rect 12012 60356 12036 60358
rect 12092 60356 12116 60358
rect 12172 60356 12196 60358
rect 12252 60356 12258 60358
rect 11950 60347 12258 60356
rect 11950 59324 12258 59333
rect 11950 59322 11956 59324
rect 12012 59322 12036 59324
rect 12092 59322 12116 59324
rect 12172 59322 12196 59324
rect 12252 59322 12258 59324
rect 12012 59270 12014 59322
rect 12194 59270 12196 59322
rect 11950 59268 11956 59270
rect 12012 59268 12036 59270
rect 12092 59268 12116 59270
rect 12172 59268 12196 59270
rect 12252 59268 12258 59270
rect 11950 59259 12258 59268
rect 11950 58236 12258 58245
rect 11950 58234 11956 58236
rect 12012 58234 12036 58236
rect 12092 58234 12116 58236
rect 12172 58234 12196 58236
rect 12252 58234 12258 58236
rect 12012 58182 12014 58234
rect 12194 58182 12196 58234
rect 11950 58180 11956 58182
rect 12012 58180 12036 58182
rect 12092 58180 12116 58182
rect 12172 58180 12196 58182
rect 12252 58180 12258 58182
rect 11950 58171 12258 58180
rect 11950 57148 12258 57157
rect 11950 57146 11956 57148
rect 12012 57146 12036 57148
rect 12092 57146 12116 57148
rect 12172 57146 12196 57148
rect 12252 57146 12258 57148
rect 12012 57094 12014 57146
rect 12194 57094 12196 57146
rect 11950 57092 11956 57094
rect 12012 57092 12036 57094
rect 12092 57092 12116 57094
rect 12172 57092 12196 57094
rect 12252 57092 12258 57094
rect 11950 57083 12258 57092
rect 11950 56060 12258 56069
rect 11950 56058 11956 56060
rect 12012 56058 12036 56060
rect 12092 56058 12116 56060
rect 12172 56058 12196 56060
rect 12252 56058 12258 56060
rect 12012 56006 12014 56058
rect 12194 56006 12196 56058
rect 11950 56004 11956 56006
rect 12012 56004 12036 56006
rect 12092 56004 12116 56006
rect 12172 56004 12196 56006
rect 12252 56004 12258 56006
rect 11950 55995 12258 56004
rect 11950 54972 12258 54981
rect 11950 54970 11956 54972
rect 12012 54970 12036 54972
rect 12092 54970 12116 54972
rect 12172 54970 12196 54972
rect 12252 54970 12258 54972
rect 12012 54918 12014 54970
rect 12194 54918 12196 54970
rect 11950 54916 11956 54918
rect 12012 54916 12036 54918
rect 12092 54916 12116 54918
rect 12172 54916 12196 54918
rect 12252 54916 12258 54918
rect 11950 54907 12258 54916
rect 11950 53884 12258 53893
rect 11950 53882 11956 53884
rect 12012 53882 12036 53884
rect 12092 53882 12116 53884
rect 12172 53882 12196 53884
rect 12252 53882 12258 53884
rect 12012 53830 12014 53882
rect 12194 53830 12196 53882
rect 11950 53828 11956 53830
rect 12012 53828 12036 53830
rect 12092 53828 12116 53830
rect 12172 53828 12196 53830
rect 12252 53828 12258 53830
rect 11950 53819 12258 53828
rect 11950 52796 12258 52805
rect 11950 52794 11956 52796
rect 12012 52794 12036 52796
rect 12092 52794 12116 52796
rect 12172 52794 12196 52796
rect 12252 52794 12258 52796
rect 12012 52742 12014 52794
rect 12194 52742 12196 52794
rect 11950 52740 11956 52742
rect 12012 52740 12036 52742
rect 12092 52740 12116 52742
rect 12172 52740 12196 52742
rect 12252 52740 12258 52742
rect 11950 52731 12258 52740
rect 11950 51708 12258 51717
rect 11950 51706 11956 51708
rect 12012 51706 12036 51708
rect 12092 51706 12116 51708
rect 12172 51706 12196 51708
rect 12252 51706 12258 51708
rect 12012 51654 12014 51706
rect 12194 51654 12196 51706
rect 11950 51652 11956 51654
rect 12012 51652 12036 51654
rect 12092 51652 12116 51654
rect 12172 51652 12196 51654
rect 12252 51652 12258 51654
rect 11950 51643 12258 51652
rect 11950 50620 12258 50629
rect 11950 50618 11956 50620
rect 12012 50618 12036 50620
rect 12092 50618 12116 50620
rect 12172 50618 12196 50620
rect 12252 50618 12258 50620
rect 12012 50566 12014 50618
rect 12194 50566 12196 50618
rect 11950 50564 11956 50566
rect 12012 50564 12036 50566
rect 12092 50564 12116 50566
rect 12172 50564 12196 50566
rect 12252 50564 12258 50566
rect 11950 50555 12258 50564
rect 11950 49532 12258 49541
rect 11950 49530 11956 49532
rect 12012 49530 12036 49532
rect 12092 49530 12116 49532
rect 12172 49530 12196 49532
rect 12252 49530 12258 49532
rect 12012 49478 12014 49530
rect 12194 49478 12196 49530
rect 11950 49476 11956 49478
rect 12012 49476 12036 49478
rect 12092 49476 12116 49478
rect 12172 49476 12196 49478
rect 12252 49476 12258 49478
rect 11950 49467 12258 49476
rect 11950 48444 12258 48453
rect 11950 48442 11956 48444
rect 12012 48442 12036 48444
rect 12092 48442 12116 48444
rect 12172 48442 12196 48444
rect 12252 48442 12258 48444
rect 12012 48390 12014 48442
rect 12194 48390 12196 48442
rect 11950 48388 11956 48390
rect 12012 48388 12036 48390
rect 12092 48388 12116 48390
rect 12172 48388 12196 48390
rect 12252 48388 12258 48390
rect 11950 48379 12258 48388
rect 11950 47356 12258 47365
rect 11950 47354 11956 47356
rect 12012 47354 12036 47356
rect 12092 47354 12116 47356
rect 12172 47354 12196 47356
rect 12252 47354 12258 47356
rect 12012 47302 12014 47354
rect 12194 47302 12196 47354
rect 11950 47300 11956 47302
rect 12012 47300 12036 47302
rect 12092 47300 12116 47302
rect 12172 47300 12196 47302
rect 12252 47300 12258 47302
rect 11950 47291 12258 47300
rect 11950 46268 12258 46277
rect 11950 46266 11956 46268
rect 12012 46266 12036 46268
rect 12092 46266 12116 46268
rect 12172 46266 12196 46268
rect 12252 46266 12258 46268
rect 12012 46214 12014 46266
rect 12194 46214 12196 46266
rect 11950 46212 11956 46214
rect 12012 46212 12036 46214
rect 12092 46212 12116 46214
rect 12172 46212 12196 46214
rect 12252 46212 12258 46214
rect 11950 46203 12258 46212
rect 11950 45180 12258 45189
rect 11950 45178 11956 45180
rect 12012 45178 12036 45180
rect 12092 45178 12116 45180
rect 12172 45178 12196 45180
rect 12252 45178 12258 45180
rect 12012 45126 12014 45178
rect 12194 45126 12196 45178
rect 11950 45124 11956 45126
rect 12012 45124 12036 45126
rect 12092 45124 12116 45126
rect 12172 45124 12196 45126
rect 12252 45124 12258 45126
rect 11950 45115 12258 45124
rect 12360 44946 12388 65418
rect 12610 65308 12918 65317
rect 12610 65306 12616 65308
rect 12672 65306 12696 65308
rect 12752 65306 12776 65308
rect 12832 65306 12856 65308
rect 12912 65306 12918 65308
rect 12672 65254 12674 65306
rect 12854 65254 12856 65306
rect 12610 65252 12616 65254
rect 12672 65252 12696 65254
rect 12752 65252 12776 65254
rect 12832 65252 12856 65254
rect 12912 65252 12918 65254
rect 12610 65243 12918 65252
rect 12610 64220 12918 64229
rect 12610 64218 12616 64220
rect 12672 64218 12696 64220
rect 12752 64218 12776 64220
rect 12832 64218 12856 64220
rect 12912 64218 12918 64220
rect 12672 64166 12674 64218
rect 12854 64166 12856 64218
rect 12610 64164 12616 64166
rect 12672 64164 12696 64166
rect 12752 64164 12776 64166
rect 12832 64164 12856 64166
rect 12912 64164 12918 64166
rect 12610 64155 12918 64164
rect 12610 63132 12918 63141
rect 12610 63130 12616 63132
rect 12672 63130 12696 63132
rect 12752 63130 12776 63132
rect 12832 63130 12856 63132
rect 12912 63130 12918 63132
rect 12672 63078 12674 63130
rect 12854 63078 12856 63130
rect 12610 63076 12616 63078
rect 12672 63076 12696 63078
rect 12752 63076 12776 63078
rect 12832 63076 12856 63078
rect 12912 63076 12918 63078
rect 12610 63067 12918 63076
rect 13004 62914 13032 67594
rect 13096 65686 13124 67662
rect 13188 67250 13216 68750
rect 13268 68740 13320 68746
rect 13268 68682 13320 68688
rect 13176 67244 13228 67250
rect 13176 67186 13228 67192
rect 13188 66094 13216 67186
rect 13176 66088 13228 66094
rect 13176 66030 13228 66036
rect 13084 65680 13136 65686
rect 13084 65622 13136 65628
rect 13188 64874 13216 66030
rect 12912 62886 13032 62914
rect 13096 64846 13216 64874
rect 12912 62490 12940 62886
rect 12900 62484 12952 62490
rect 12900 62426 12952 62432
rect 12912 62286 12940 62426
rect 12532 62280 12584 62286
rect 12532 62222 12584 62228
rect 12900 62280 12952 62286
rect 12900 62222 12952 62228
rect 12544 59498 12572 62222
rect 12610 62044 12918 62053
rect 12610 62042 12616 62044
rect 12672 62042 12696 62044
rect 12752 62042 12776 62044
rect 12832 62042 12856 62044
rect 12912 62042 12918 62044
rect 12672 61990 12674 62042
rect 12854 61990 12856 62042
rect 12610 61988 12616 61990
rect 12672 61988 12696 61990
rect 12752 61988 12776 61990
rect 12832 61988 12856 61990
rect 12912 61988 12918 61990
rect 12610 61979 12918 61988
rect 12610 60956 12918 60965
rect 12610 60954 12616 60956
rect 12672 60954 12696 60956
rect 12752 60954 12776 60956
rect 12832 60954 12856 60956
rect 12912 60954 12918 60956
rect 12672 60902 12674 60954
rect 12854 60902 12856 60954
rect 12610 60900 12616 60902
rect 12672 60900 12696 60902
rect 12752 60900 12776 60902
rect 12832 60900 12856 60902
rect 12912 60900 12918 60902
rect 12610 60891 12918 60900
rect 12610 59868 12918 59877
rect 12610 59866 12616 59868
rect 12672 59866 12696 59868
rect 12752 59866 12776 59868
rect 12832 59866 12856 59868
rect 12912 59866 12918 59868
rect 12672 59814 12674 59866
rect 12854 59814 12856 59866
rect 12610 59812 12616 59814
rect 12672 59812 12696 59814
rect 12752 59812 12776 59814
rect 12832 59812 12856 59814
rect 12912 59812 12918 59814
rect 12610 59803 12918 59812
rect 12532 59492 12584 59498
rect 12532 59434 12584 59440
rect 12610 58780 12918 58789
rect 12610 58778 12616 58780
rect 12672 58778 12696 58780
rect 12752 58778 12776 58780
rect 12832 58778 12856 58780
rect 12912 58778 12918 58780
rect 12672 58726 12674 58778
rect 12854 58726 12856 58778
rect 12610 58724 12616 58726
rect 12672 58724 12696 58726
rect 12752 58724 12776 58726
rect 12832 58724 12856 58726
rect 12912 58724 12918 58726
rect 12610 58715 12918 58724
rect 12440 57792 12492 57798
rect 12440 57734 12492 57740
rect 12452 50726 12480 57734
rect 12610 57692 12918 57701
rect 12610 57690 12616 57692
rect 12672 57690 12696 57692
rect 12752 57690 12776 57692
rect 12832 57690 12856 57692
rect 12912 57690 12918 57692
rect 12672 57638 12674 57690
rect 12854 57638 12856 57690
rect 12610 57636 12616 57638
rect 12672 57636 12696 57638
rect 12752 57636 12776 57638
rect 12832 57636 12856 57638
rect 12912 57636 12918 57638
rect 12610 57627 12918 57636
rect 12610 56604 12918 56613
rect 12610 56602 12616 56604
rect 12672 56602 12696 56604
rect 12752 56602 12776 56604
rect 12832 56602 12856 56604
rect 12912 56602 12918 56604
rect 12672 56550 12674 56602
rect 12854 56550 12856 56602
rect 12610 56548 12616 56550
rect 12672 56548 12696 56550
rect 12752 56548 12776 56550
rect 12832 56548 12856 56550
rect 12912 56548 12918 56550
rect 12610 56539 12918 56548
rect 12610 55516 12918 55525
rect 12610 55514 12616 55516
rect 12672 55514 12696 55516
rect 12752 55514 12776 55516
rect 12832 55514 12856 55516
rect 12912 55514 12918 55516
rect 12672 55462 12674 55514
rect 12854 55462 12856 55514
rect 12610 55460 12616 55462
rect 12672 55460 12696 55462
rect 12752 55460 12776 55462
rect 12832 55460 12856 55462
rect 12912 55460 12918 55462
rect 12610 55451 12918 55460
rect 12610 54428 12918 54437
rect 12610 54426 12616 54428
rect 12672 54426 12696 54428
rect 12752 54426 12776 54428
rect 12832 54426 12856 54428
rect 12912 54426 12918 54428
rect 12672 54374 12674 54426
rect 12854 54374 12856 54426
rect 12610 54372 12616 54374
rect 12672 54372 12696 54374
rect 12752 54372 12776 54374
rect 12832 54372 12856 54374
rect 12912 54372 12918 54374
rect 12610 54363 12918 54372
rect 12610 53340 12918 53349
rect 12610 53338 12616 53340
rect 12672 53338 12696 53340
rect 12752 53338 12776 53340
rect 12832 53338 12856 53340
rect 12912 53338 12918 53340
rect 12672 53286 12674 53338
rect 12854 53286 12856 53338
rect 12610 53284 12616 53286
rect 12672 53284 12696 53286
rect 12752 53284 12776 53286
rect 12832 53284 12856 53286
rect 12912 53284 12918 53286
rect 12610 53275 12918 53284
rect 12610 52252 12918 52261
rect 12610 52250 12616 52252
rect 12672 52250 12696 52252
rect 12752 52250 12776 52252
rect 12832 52250 12856 52252
rect 12912 52250 12918 52252
rect 12672 52198 12674 52250
rect 12854 52198 12856 52250
rect 12610 52196 12616 52198
rect 12672 52196 12696 52198
rect 12752 52196 12776 52198
rect 12832 52196 12856 52198
rect 12912 52196 12918 52198
rect 12610 52187 12918 52196
rect 12610 51164 12918 51173
rect 12610 51162 12616 51164
rect 12672 51162 12696 51164
rect 12752 51162 12776 51164
rect 12832 51162 12856 51164
rect 12912 51162 12918 51164
rect 12672 51110 12674 51162
rect 12854 51110 12856 51162
rect 12610 51108 12616 51110
rect 12672 51108 12696 51110
rect 12752 51108 12776 51110
rect 12832 51108 12856 51110
rect 12912 51108 12918 51110
rect 12610 51099 12918 51108
rect 12992 50924 13044 50930
rect 12992 50866 13044 50872
rect 12440 50720 12492 50726
rect 12440 50662 12492 50668
rect 12808 50720 12860 50726
rect 12808 50662 12860 50668
rect 12348 44940 12400 44946
rect 12348 44882 12400 44888
rect 12452 44470 12480 50662
rect 12820 50318 12848 50662
rect 12808 50312 12860 50318
rect 12808 50254 12860 50260
rect 12610 50076 12918 50085
rect 12610 50074 12616 50076
rect 12672 50074 12696 50076
rect 12752 50074 12776 50076
rect 12832 50074 12856 50076
rect 12912 50074 12918 50076
rect 12672 50022 12674 50074
rect 12854 50022 12856 50074
rect 12610 50020 12616 50022
rect 12672 50020 12696 50022
rect 12752 50020 12776 50022
rect 12832 50020 12856 50022
rect 12912 50020 12918 50022
rect 12610 50011 12918 50020
rect 12610 48988 12918 48997
rect 12610 48986 12616 48988
rect 12672 48986 12696 48988
rect 12752 48986 12776 48988
rect 12832 48986 12856 48988
rect 12912 48986 12918 48988
rect 12672 48934 12674 48986
rect 12854 48934 12856 48986
rect 12610 48932 12616 48934
rect 12672 48932 12696 48934
rect 12752 48932 12776 48934
rect 12832 48932 12856 48934
rect 12912 48932 12918 48934
rect 12610 48923 12918 48932
rect 12610 47900 12918 47909
rect 12610 47898 12616 47900
rect 12672 47898 12696 47900
rect 12752 47898 12776 47900
rect 12832 47898 12856 47900
rect 12912 47898 12918 47900
rect 12672 47846 12674 47898
rect 12854 47846 12856 47898
rect 12610 47844 12616 47846
rect 12672 47844 12696 47846
rect 12752 47844 12776 47846
rect 12832 47844 12856 47846
rect 12912 47844 12918 47846
rect 12610 47835 12918 47844
rect 12610 46812 12918 46821
rect 12610 46810 12616 46812
rect 12672 46810 12696 46812
rect 12752 46810 12776 46812
rect 12832 46810 12856 46812
rect 12912 46810 12918 46812
rect 12672 46758 12674 46810
rect 12854 46758 12856 46810
rect 12610 46756 12616 46758
rect 12672 46756 12696 46758
rect 12752 46756 12776 46758
rect 12832 46756 12856 46758
rect 12912 46756 12918 46758
rect 12610 46747 12918 46756
rect 12610 45724 12918 45733
rect 12610 45722 12616 45724
rect 12672 45722 12696 45724
rect 12752 45722 12776 45724
rect 12832 45722 12856 45724
rect 12912 45722 12918 45724
rect 12672 45670 12674 45722
rect 12854 45670 12856 45722
rect 12610 45668 12616 45670
rect 12672 45668 12696 45670
rect 12752 45668 12776 45670
rect 12832 45668 12856 45670
rect 12912 45668 12918 45670
rect 12610 45659 12918 45668
rect 12610 44636 12918 44645
rect 12610 44634 12616 44636
rect 12672 44634 12696 44636
rect 12752 44634 12776 44636
rect 12832 44634 12856 44636
rect 12912 44634 12918 44636
rect 12672 44582 12674 44634
rect 12854 44582 12856 44634
rect 12610 44580 12616 44582
rect 12672 44580 12696 44582
rect 12752 44580 12776 44582
rect 12832 44580 12856 44582
rect 12912 44580 12918 44582
rect 12610 44571 12918 44580
rect 12440 44464 12492 44470
rect 12440 44406 12492 44412
rect 11950 44092 12258 44101
rect 11950 44090 11956 44092
rect 12012 44090 12036 44092
rect 12092 44090 12116 44092
rect 12172 44090 12196 44092
rect 12252 44090 12258 44092
rect 12012 44038 12014 44090
rect 12194 44038 12196 44090
rect 11950 44036 11956 44038
rect 12012 44036 12036 44038
rect 12092 44036 12116 44038
rect 12172 44036 12196 44038
rect 12252 44036 12258 44038
rect 11950 44027 12258 44036
rect 12610 43548 12918 43557
rect 12610 43546 12616 43548
rect 12672 43546 12696 43548
rect 12752 43546 12776 43548
rect 12832 43546 12856 43548
rect 12912 43546 12918 43548
rect 12672 43494 12674 43546
rect 12854 43494 12856 43546
rect 12610 43492 12616 43494
rect 12672 43492 12696 43494
rect 12752 43492 12776 43494
rect 12832 43492 12856 43494
rect 12912 43492 12918 43494
rect 12610 43483 12918 43492
rect 12348 43172 12400 43178
rect 12348 43114 12400 43120
rect 11950 43004 12258 43013
rect 11950 43002 11956 43004
rect 12012 43002 12036 43004
rect 12092 43002 12116 43004
rect 12172 43002 12196 43004
rect 12252 43002 12258 43004
rect 12012 42950 12014 43002
rect 12194 42950 12196 43002
rect 11950 42948 11956 42950
rect 12012 42948 12036 42950
rect 12092 42948 12116 42950
rect 12172 42948 12196 42950
rect 12252 42948 12258 42950
rect 11950 42939 12258 42948
rect 11950 41916 12258 41925
rect 11950 41914 11956 41916
rect 12012 41914 12036 41916
rect 12092 41914 12116 41916
rect 12172 41914 12196 41916
rect 12252 41914 12258 41916
rect 12012 41862 12014 41914
rect 12194 41862 12196 41914
rect 11950 41860 11956 41862
rect 12012 41860 12036 41862
rect 12092 41860 12116 41862
rect 12172 41860 12196 41862
rect 12252 41860 12258 41862
rect 11950 41851 12258 41860
rect 11796 41472 11848 41478
rect 11796 41414 11848 41420
rect 11950 40828 12258 40837
rect 11950 40826 11956 40828
rect 12012 40826 12036 40828
rect 12092 40826 12116 40828
rect 12172 40826 12196 40828
rect 12252 40826 12258 40828
rect 12012 40774 12014 40826
rect 12194 40774 12196 40826
rect 11950 40772 11956 40774
rect 12012 40772 12036 40774
rect 12092 40772 12116 40774
rect 12172 40772 12196 40774
rect 12252 40772 12258 40774
rect 11950 40763 12258 40772
rect 11950 39740 12258 39749
rect 11950 39738 11956 39740
rect 12012 39738 12036 39740
rect 12092 39738 12116 39740
rect 12172 39738 12196 39740
rect 12252 39738 12258 39740
rect 12012 39686 12014 39738
rect 12194 39686 12196 39738
rect 11950 39684 11956 39686
rect 12012 39684 12036 39686
rect 12092 39684 12116 39686
rect 12172 39684 12196 39686
rect 12252 39684 12258 39686
rect 11950 39675 12258 39684
rect 11950 38652 12258 38661
rect 11950 38650 11956 38652
rect 12012 38650 12036 38652
rect 12092 38650 12116 38652
rect 12172 38650 12196 38652
rect 12252 38650 12258 38652
rect 12012 38598 12014 38650
rect 12194 38598 12196 38650
rect 11950 38596 11956 38598
rect 12012 38596 12036 38598
rect 12092 38596 12116 38598
rect 12172 38596 12196 38598
rect 12252 38596 12258 38598
rect 11950 38587 12258 38596
rect 11950 37564 12258 37573
rect 11950 37562 11956 37564
rect 12012 37562 12036 37564
rect 12092 37562 12116 37564
rect 12172 37562 12196 37564
rect 12252 37562 12258 37564
rect 12012 37510 12014 37562
rect 12194 37510 12196 37562
rect 11950 37508 11956 37510
rect 12012 37508 12036 37510
rect 12092 37508 12116 37510
rect 12172 37508 12196 37510
rect 12252 37508 12258 37510
rect 11950 37499 12258 37508
rect 11950 36476 12258 36485
rect 11950 36474 11956 36476
rect 12012 36474 12036 36476
rect 12092 36474 12116 36476
rect 12172 36474 12196 36476
rect 12252 36474 12258 36476
rect 12012 36422 12014 36474
rect 12194 36422 12196 36474
rect 11950 36420 11956 36422
rect 12012 36420 12036 36422
rect 12092 36420 12116 36422
rect 12172 36420 12196 36422
rect 12252 36420 12258 36422
rect 11950 36411 12258 36420
rect 11704 36372 11756 36378
rect 11704 36314 11756 36320
rect 11950 35388 12258 35397
rect 11950 35386 11956 35388
rect 12012 35386 12036 35388
rect 12092 35386 12116 35388
rect 12172 35386 12196 35388
rect 12252 35386 12258 35388
rect 12012 35334 12014 35386
rect 12194 35334 12196 35386
rect 11950 35332 11956 35334
rect 12012 35332 12036 35334
rect 12092 35332 12116 35334
rect 12172 35332 12196 35334
rect 12252 35332 12258 35334
rect 11950 35323 12258 35332
rect 11950 34300 12258 34309
rect 11950 34298 11956 34300
rect 12012 34298 12036 34300
rect 12092 34298 12116 34300
rect 12172 34298 12196 34300
rect 12252 34298 12258 34300
rect 12012 34246 12014 34298
rect 12194 34246 12196 34298
rect 11950 34244 11956 34246
rect 12012 34244 12036 34246
rect 12092 34244 12116 34246
rect 12172 34244 12196 34246
rect 12252 34244 12258 34246
rect 11950 34235 12258 34244
rect 11704 33924 11756 33930
rect 11704 33866 11756 33872
rect 11612 32972 11664 32978
rect 11612 32914 11664 32920
rect 11520 29028 11572 29034
rect 11520 28970 11572 28976
rect 11716 28014 11744 33866
rect 11950 33212 12258 33221
rect 11950 33210 11956 33212
rect 12012 33210 12036 33212
rect 12092 33210 12116 33212
rect 12172 33210 12196 33212
rect 12252 33210 12258 33212
rect 12012 33158 12014 33210
rect 12194 33158 12196 33210
rect 11950 33156 11956 33158
rect 12012 33156 12036 33158
rect 12092 33156 12116 33158
rect 12172 33156 12196 33158
rect 12252 33156 12258 33158
rect 11950 33147 12258 33156
rect 11950 32124 12258 32133
rect 11950 32122 11956 32124
rect 12012 32122 12036 32124
rect 12092 32122 12116 32124
rect 12172 32122 12196 32124
rect 12252 32122 12258 32124
rect 12012 32070 12014 32122
rect 12194 32070 12196 32122
rect 11950 32068 11956 32070
rect 12012 32068 12036 32070
rect 12092 32068 12116 32070
rect 12172 32068 12196 32070
rect 12252 32068 12258 32070
rect 11950 32059 12258 32068
rect 11950 31036 12258 31045
rect 11950 31034 11956 31036
rect 12012 31034 12036 31036
rect 12092 31034 12116 31036
rect 12172 31034 12196 31036
rect 12252 31034 12258 31036
rect 12012 30982 12014 31034
rect 12194 30982 12196 31034
rect 11950 30980 11956 30982
rect 12012 30980 12036 30982
rect 12092 30980 12116 30982
rect 12172 30980 12196 30982
rect 12252 30980 12258 30982
rect 11950 30971 12258 30980
rect 11950 29948 12258 29957
rect 11950 29946 11956 29948
rect 12012 29946 12036 29948
rect 12092 29946 12116 29948
rect 12172 29946 12196 29948
rect 12252 29946 12258 29948
rect 12012 29894 12014 29946
rect 12194 29894 12196 29946
rect 11950 29892 11956 29894
rect 12012 29892 12036 29894
rect 12092 29892 12116 29894
rect 12172 29892 12196 29894
rect 12252 29892 12258 29894
rect 11950 29883 12258 29892
rect 12256 29300 12308 29306
rect 12256 29242 12308 29248
rect 12268 29170 12296 29242
rect 11980 29164 12032 29170
rect 11980 29106 12032 29112
rect 12256 29164 12308 29170
rect 12256 29106 12308 29112
rect 11992 29034 12020 29106
rect 11796 29028 11848 29034
rect 11796 28970 11848 28976
rect 11980 29028 12032 29034
rect 11980 28970 12032 28976
rect 11704 28008 11756 28014
rect 11704 27950 11756 27956
rect 11716 23254 11744 27950
rect 11704 23248 11756 23254
rect 11704 23190 11756 23196
rect 11612 22772 11664 22778
rect 11612 22714 11664 22720
rect 11624 22166 11652 22714
rect 11612 22160 11664 22166
rect 11612 22102 11664 22108
rect 11704 21412 11756 21418
rect 11704 21354 11756 21360
rect 11152 3528 11204 3534
rect 11152 3470 11204 3476
rect 11716 2514 11744 21354
rect 11808 15910 11836 28970
rect 11950 28860 12258 28869
rect 11950 28858 11956 28860
rect 12012 28858 12036 28860
rect 12092 28858 12116 28860
rect 12172 28858 12196 28860
rect 12252 28858 12258 28860
rect 12012 28806 12014 28858
rect 12194 28806 12196 28858
rect 11950 28804 11956 28806
rect 12012 28804 12036 28806
rect 12092 28804 12116 28806
rect 12172 28804 12196 28806
rect 12252 28804 12258 28806
rect 11950 28795 12258 28804
rect 11950 27772 12258 27781
rect 11950 27770 11956 27772
rect 12012 27770 12036 27772
rect 12092 27770 12116 27772
rect 12172 27770 12196 27772
rect 12252 27770 12258 27772
rect 12012 27718 12014 27770
rect 12194 27718 12196 27770
rect 11950 27716 11956 27718
rect 12012 27716 12036 27718
rect 12092 27716 12116 27718
rect 12172 27716 12196 27718
rect 12252 27716 12258 27718
rect 11950 27707 12258 27716
rect 11950 26684 12258 26693
rect 11950 26682 11956 26684
rect 12012 26682 12036 26684
rect 12092 26682 12116 26684
rect 12172 26682 12196 26684
rect 12252 26682 12258 26684
rect 12012 26630 12014 26682
rect 12194 26630 12196 26682
rect 11950 26628 11956 26630
rect 12012 26628 12036 26630
rect 12092 26628 12116 26630
rect 12172 26628 12196 26630
rect 12252 26628 12258 26630
rect 11950 26619 12258 26628
rect 11950 25596 12258 25605
rect 11950 25594 11956 25596
rect 12012 25594 12036 25596
rect 12092 25594 12116 25596
rect 12172 25594 12196 25596
rect 12252 25594 12258 25596
rect 12012 25542 12014 25594
rect 12194 25542 12196 25594
rect 11950 25540 11956 25542
rect 12012 25540 12036 25542
rect 12092 25540 12116 25542
rect 12172 25540 12196 25542
rect 12252 25540 12258 25542
rect 11950 25531 12258 25540
rect 11950 24508 12258 24517
rect 11950 24506 11956 24508
rect 12012 24506 12036 24508
rect 12092 24506 12116 24508
rect 12172 24506 12196 24508
rect 12252 24506 12258 24508
rect 12012 24454 12014 24506
rect 12194 24454 12196 24506
rect 11950 24452 11956 24454
rect 12012 24452 12036 24454
rect 12092 24452 12116 24454
rect 12172 24452 12196 24454
rect 12252 24452 12258 24454
rect 11950 24443 12258 24452
rect 12360 24206 12388 43114
rect 13004 42702 13032 50866
rect 13096 49706 13124 64846
rect 13280 62150 13308 68682
rect 13636 67856 13688 67862
rect 13636 67798 13688 67804
rect 13452 67720 13504 67726
rect 13452 67662 13504 67668
rect 13544 67720 13596 67726
rect 13544 67662 13596 67668
rect 13464 64530 13492 67662
rect 13452 64524 13504 64530
rect 13452 64466 13504 64472
rect 13556 64462 13584 67662
rect 13544 64456 13596 64462
rect 13544 64398 13596 64404
rect 13360 62756 13412 62762
rect 13360 62698 13412 62704
rect 13372 62286 13400 62698
rect 13360 62280 13412 62286
rect 13360 62222 13412 62228
rect 13268 62144 13320 62150
rect 13268 62086 13320 62092
rect 13452 55208 13504 55214
rect 13452 55150 13504 55156
rect 13176 54052 13228 54058
rect 13176 53994 13228 54000
rect 13084 49700 13136 49706
rect 13084 49642 13136 49648
rect 12992 42696 13044 42702
rect 12992 42638 13044 42644
rect 12610 42460 12918 42469
rect 12610 42458 12616 42460
rect 12672 42458 12696 42460
rect 12752 42458 12776 42460
rect 12832 42458 12856 42460
rect 12912 42458 12918 42460
rect 12672 42406 12674 42458
rect 12854 42406 12856 42458
rect 12610 42404 12616 42406
rect 12672 42404 12696 42406
rect 12752 42404 12776 42406
rect 12832 42404 12856 42406
rect 12912 42404 12918 42406
rect 12610 42395 12918 42404
rect 12610 41372 12918 41381
rect 12610 41370 12616 41372
rect 12672 41370 12696 41372
rect 12752 41370 12776 41372
rect 12832 41370 12856 41372
rect 12912 41370 12918 41372
rect 12672 41318 12674 41370
rect 12854 41318 12856 41370
rect 12610 41316 12616 41318
rect 12672 41316 12696 41318
rect 12752 41316 12776 41318
rect 12832 41316 12856 41318
rect 12912 41316 12918 41318
rect 12610 41307 12918 41316
rect 12610 40284 12918 40293
rect 12610 40282 12616 40284
rect 12672 40282 12696 40284
rect 12752 40282 12776 40284
rect 12832 40282 12856 40284
rect 12912 40282 12918 40284
rect 12672 40230 12674 40282
rect 12854 40230 12856 40282
rect 12610 40228 12616 40230
rect 12672 40228 12696 40230
rect 12752 40228 12776 40230
rect 12832 40228 12856 40230
rect 12912 40228 12918 40230
rect 12610 40219 12918 40228
rect 12610 39196 12918 39205
rect 12610 39194 12616 39196
rect 12672 39194 12696 39196
rect 12752 39194 12776 39196
rect 12832 39194 12856 39196
rect 12912 39194 12918 39196
rect 12672 39142 12674 39194
rect 12854 39142 12856 39194
rect 12610 39140 12616 39142
rect 12672 39140 12696 39142
rect 12752 39140 12776 39142
rect 12832 39140 12856 39142
rect 12912 39140 12918 39142
rect 12610 39131 12918 39140
rect 12610 38108 12918 38117
rect 12610 38106 12616 38108
rect 12672 38106 12696 38108
rect 12752 38106 12776 38108
rect 12832 38106 12856 38108
rect 12912 38106 12918 38108
rect 12672 38054 12674 38106
rect 12854 38054 12856 38106
rect 12610 38052 12616 38054
rect 12672 38052 12696 38054
rect 12752 38052 12776 38054
rect 12832 38052 12856 38054
rect 12912 38052 12918 38054
rect 12610 38043 12918 38052
rect 12610 37020 12918 37029
rect 12610 37018 12616 37020
rect 12672 37018 12696 37020
rect 12752 37018 12776 37020
rect 12832 37018 12856 37020
rect 12912 37018 12918 37020
rect 12672 36966 12674 37018
rect 12854 36966 12856 37018
rect 12610 36964 12616 36966
rect 12672 36964 12696 36966
rect 12752 36964 12776 36966
rect 12832 36964 12856 36966
rect 12912 36964 12918 36966
rect 12610 36955 12918 36964
rect 12610 35932 12918 35941
rect 12610 35930 12616 35932
rect 12672 35930 12696 35932
rect 12752 35930 12776 35932
rect 12832 35930 12856 35932
rect 12912 35930 12918 35932
rect 12672 35878 12674 35930
rect 12854 35878 12856 35930
rect 12610 35876 12616 35878
rect 12672 35876 12696 35878
rect 12752 35876 12776 35878
rect 12832 35876 12856 35878
rect 12912 35876 12918 35878
rect 12610 35867 12918 35876
rect 12440 35148 12492 35154
rect 12440 35090 12492 35096
rect 12348 24200 12400 24206
rect 12348 24142 12400 24148
rect 11950 23420 12258 23429
rect 11950 23418 11956 23420
rect 12012 23418 12036 23420
rect 12092 23418 12116 23420
rect 12172 23418 12196 23420
rect 12252 23418 12258 23420
rect 12012 23366 12014 23418
rect 12194 23366 12196 23418
rect 11950 23364 11956 23366
rect 12012 23364 12036 23366
rect 12092 23364 12116 23366
rect 12172 23364 12196 23366
rect 12252 23364 12258 23366
rect 11950 23355 12258 23364
rect 12256 23248 12308 23254
rect 12256 23190 12308 23196
rect 11980 22772 12032 22778
rect 11980 22714 12032 22720
rect 11992 22506 12020 22714
rect 12268 22710 12296 23190
rect 12256 22704 12308 22710
rect 12256 22646 12308 22652
rect 11980 22500 12032 22506
rect 11980 22442 12032 22448
rect 11950 22332 12258 22341
rect 11950 22330 11956 22332
rect 12012 22330 12036 22332
rect 12092 22330 12116 22332
rect 12172 22330 12196 22332
rect 12252 22330 12258 22332
rect 12012 22278 12014 22330
rect 12194 22278 12196 22330
rect 11950 22276 11956 22278
rect 12012 22276 12036 22278
rect 12092 22276 12116 22278
rect 12172 22276 12196 22278
rect 12252 22276 12258 22278
rect 11950 22267 12258 22276
rect 11950 21244 12258 21253
rect 11950 21242 11956 21244
rect 12012 21242 12036 21244
rect 12092 21242 12116 21244
rect 12172 21242 12196 21244
rect 12252 21242 12258 21244
rect 12012 21190 12014 21242
rect 12194 21190 12196 21242
rect 11950 21188 11956 21190
rect 12012 21188 12036 21190
rect 12092 21188 12116 21190
rect 12172 21188 12196 21190
rect 12252 21188 12258 21190
rect 11950 21179 12258 21188
rect 11950 20156 12258 20165
rect 11950 20154 11956 20156
rect 12012 20154 12036 20156
rect 12092 20154 12116 20156
rect 12172 20154 12196 20156
rect 12252 20154 12258 20156
rect 12012 20102 12014 20154
rect 12194 20102 12196 20154
rect 11950 20100 11956 20102
rect 12012 20100 12036 20102
rect 12092 20100 12116 20102
rect 12172 20100 12196 20102
rect 12252 20100 12258 20102
rect 11950 20091 12258 20100
rect 11950 19068 12258 19077
rect 11950 19066 11956 19068
rect 12012 19066 12036 19068
rect 12092 19066 12116 19068
rect 12172 19066 12196 19068
rect 12252 19066 12258 19068
rect 12012 19014 12014 19066
rect 12194 19014 12196 19066
rect 11950 19012 11956 19014
rect 12012 19012 12036 19014
rect 12092 19012 12116 19014
rect 12172 19012 12196 19014
rect 12252 19012 12258 19014
rect 11950 19003 12258 19012
rect 11950 17980 12258 17989
rect 11950 17978 11956 17980
rect 12012 17978 12036 17980
rect 12092 17978 12116 17980
rect 12172 17978 12196 17980
rect 12252 17978 12258 17980
rect 12012 17926 12014 17978
rect 12194 17926 12196 17978
rect 11950 17924 11956 17926
rect 12012 17924 12036 17926
rect 12092 17924 12116 17926
rect 12172 17924 12196 17926
rect 12252 17924 12258 17926
rect 11950 17915 12258 17924
rect 11950 16892 12258 16901
rect 11950 16890 11956 16892
rect 12012 16890 12036 16892
rect 12092 16890 12116 16892
rect 12172 16890 12196 16892
rect 12252 16890 12258 16892
rect 12012 16838 12014 16890
rect 12194 16838 12196 16890
rect 11950 16836 11956 16838
rect 12012 16836 12036 16838
rect 12092 16836 12116 16838
rect 12172 16836 12196 16838
rect 12252 16836 12258 16838
rect 11950 16827 12258 16836
rect 11796 15904 11848 15910
rect 11796 15846 11848 15852
rect 11950 15804 12258 15813
rect 11950 15802 11956 15804
rect 12012 15802 12036 15804
rect 12092 15802 12116 15804
rect 12172 15802 12196 15804
rect 12252 15802 12258 15804
rect 12012 15750 12014 15802
rect 12194 15750 12196 15802
rect 11950 15748 11956 15750
rect 12012 15748 12036 15750
rect 12092 15748 12116 15750
rect 12172 15748 12196 15750
rect 12252 15748 12258 15750
rect 11950 15739 12258 15748
rect 11950 14716 12258 14725
rect 11950 14714 11956 14716
rect 12012 14714 12036 14716
rect 12092 14714 12116 14716
rect 12172 14714 12196 14716
rect 12252 14714 12258 14716
rect 12012 14662 12014 14714
rect 12194 14662 12196 14714
rect 11950 14660 11956 14662
rect 12012 14660 12036 14662
rect 12092 14660 12116 14662
rect 12172 14660 12196 14662
rect 12252 14660 12258 14662
rect 11950 14651 12258 14660
rect 11950 13628 12258 13637
rect 11950 13626 11956 13628
rect 12012 13626 12036 13628
rect 12092 13626 12116 13628
rect 12172 13626 12196 13628
rect 12252 13626 12258 13628
rect 12012 13574 12014 13626
rect 12194 13574 12196 13626
rect 11950 13572 11956 13574
rect 12012 13572 12036 13574
rect 12092 13572 12116 13574
rect 12172 13572 12196 13574
rect 12252 13572 12258 13574
rect 11950 13563 12258 13572
rect 11950 12540 12258 12549
rect 11950 12538 11956 12540
rect 12012 12538 12036 12540
rect 12092 12538 12116 12540
rect 12172 12538 12196 12540
rect 12252 12538 12258 12540
rect 12012 12486 12014 12538
rect 12194 12486 12196 12538
rect 11950 12484 11956 12486
rect 12012 12484 12036 12486
rect 12092 12484 12116 12486
rect 12172 12484 12196 12486
rect 12252 12484 12258 12486
rect 11950 12475 12258 12484
rect 11950 11452 12258 11461
rect 11950 11450 11956 11452
rect 12012 11450 12036 11452
rect 12092 11450 12116 11452
rect 12172 11450 12196 11452
rect 12252 11450 12258 11452
rect 12012 11398 12014 11450
rect 12194 11398 12196 11450
rect 11950 11396 11956 11398
rect 12012 11396 12036 11398
rect 12092 11396 12116 11398
rect 12172 11396 12196 11398
rect 12252 11396 12258 11398
rect 11950 11387 12258 11396
rect 12360 10606 12388 24142
rect 12452 21418 12480 35090
rect 12610 34844 12918 34853
rect 12610 34842 12616 34844
rect 12672 34842 12696 34844
rect 12752 34842 12776 34844
rect 12832 34842 12856 34844
rect 12912 34842 12918 34844
rect 12672 34790 12674 34842
rect 12854 34790 12856 34842
rect 12610 34788 12616 34790
rect 12672 34788 12696 34790
rect 12752 34788 12776 34790
rect 12832 34788 12856 34790
rect 12912 34788 12918 34790
rect 12610 34779 12918 34788
rect 13004 34610 13032 42638
rect 13084 35080 13136 35086
rect 13084 35022 13136 35028
rect 12992 34604 13044 34610
rect 12992 34546 13044 34552
rect 12610 33756 12918 33765
rect 12610 33754 12616 33756
rect 12672 33754 12696 33756
rect 12752 33754 12776 33756
rect 12832 33754 12856 33756
rect 12912 33754 12918 33756
rect 12672 33702 12674 33754
rect 12854 33702 12856 33754
rect 12610 33700 12616 33702
rect 12672 33700 12696 33702
rect 12752 33700 12776 33702
rect 12832 33700 12856 33702
rect 12912 33700 12918 33702
rect 12610 33691 12918 33700
rect 12992 33380 13044 33386
rect 12992 33322 13044 33328
rect 12610 32668 12918 32677
rect 12610 32666 12616 32668
rect 12672 32666 12696 32668
rect 12752 32666 12776 32668
rect 12832 32666 12856 32668
rect 12912 32666 12918 32668
rect 12672 32614 12674 32666
rect 12854 32614 12856 32666
rect 12610 32612 12616 32614
rect 12672 32612 12696 32614
rect 12752 32612 12776 32614
rect 12832 32612 12856 32614
rect 12912 32612 12918 32614
rect 12610 32603 12918 32612
rect 13004 31754 13032 33322
rect 13096 33114 13124 35022
rect 13084 33108 13136 33114
rect 13084 33050 13136 33056
rect 13004 31726 13124 31754
rect 12610 31580 12918 31589
rect 12610 31578 12616 31580
rect 12672 31578 12696 31580
rect 12752 31578 12776 31580
rect 12832 31578 12856 31580
rect 12912 31578 12918 31580
rect 12672 31526 12674 31578
rect 12854 31526 12856 31578
rect 12610 31524 12616 31526
rect 12672 31524 12696 31526
rect 12752 31524 12776 31526
rect 12832 31524 12856 31526
rect 12912 31524 12918 31526
rect 12610 31515 12918 31524
rect 12610 30492 12918 30501
rect 12610 30490 12616 30492
rect 12672 30490 12696 30492
rect 12752 30490 12776 30492
rect 12832 30490 12856 30492
rect 12912 30490 12918 30492
rect 12672 30438 12674 30490
rect 12854 30438 12856 30490
rect 12610 30436 12616 30438
rect 12672 30436 12696 30438
rect 12752 30436 12776 30438
rect 12832 30436 12856 30438
rect 12912 30436 12918 30438
rect 12610 30427 12918 30436
rect 12610 29404 12918 29413
rect 12610 29402 12616 29404
rect 12672 29402 12696 29404
rect 12752 29402 12776 29404
rect 12832 29402 12856 29404
rect 12912 29402 12918 29404
rect 12672 29350 12674 29402
rect 12854 29350 12856 29402
rect 12610 29348 12616 29350
rect 12672 29348 12696 29350
rect 12752 29348 12776 29350
rect 12832 29348 12856 29350
rect 12912 29348 12918 29350
rect 12610 29339 12918 29348
rect 12532 29232 12584 29238
rect 12532 29174 12584 29180
rect 12544 29034 12572 29174
rect 12532 29028 12584 29034
rect 12532 28970 12584 28976
rect 12610 28316 12918 28325
rect 12610 28314 12616 28316
rect 12672 28314 12696 28316
rect 12752 28314 12776 28316
rect 12832 28314 12856 28316
rect 12912 28314 12918 28316
rect 12672 28262 12674 28314
rect 12854 28262 12856 28314
rect 12610 28260 12616 28262
rect 12672 28260 12696 28262
rect 12752 28260 12776 28262
rect 12832 28260 12856 28262
rect 12912 28260 12918 28262
rect 12610 28251 12918 28260
rect 12610 27228 12918 27237
rect 12610 27226 12616 27228
rect 12672 27226 12696 27228
rect 12752 27226 12776 27228
rect 12832 27226 12856 27228
rect 12912 27226 12918 27228
rect 12672 27174 12674 27226
rect 12854 27174 12856 27226
rect 12610 27172 12616 27174
rect 12672 27172 12696 27174
rect 12752 27172 12776 27174
rect 12832 27172 12856 27174
rect 12912 27172 12918 27174
rect 12610 27163 12918 27172
rect 12610 26140 12918 26149
rect 12610 26138 12616 26140
rect 12672 26138 12696 26140
rect 12752 26138 12776 26140
rect 12832 26138 12856 26140
rect 12912 26138 12918 26140
rect 12672 26086 12674 26138
rect 12854 26086 12856 26138
rect 12610 26084 12616 26086
rect 12672 26084 12696 26086
rect 12752 26084 12776 26086
rect 12832 26084 12856 26086
rect 12912 26084 12918 26086
rect 12610 26075 12918 26084
rect 12610 25052 12918 25061
rect 12610 25050 12616 25052
rect 12672 25050 12696 25052
rect 12752 25050 12776 25052
rect 12832 25050 12856 25052
rect 12912 25050 12918 25052
rect 12672 24998 12674 25050
rect 12854 24998 12856 25050
rect 12610 24996 12616 24998
rect 12672 24996 12696 24998
rect 12752 24996 12776 24998
rect 12832 24996 12856 24998
rect 12912 24996 12918 24998
rect 12610 24987 12918 24996
rect 12610 23964 12918 23973
rect 12610 23962 12616 23964
rect 12672 23962 12696 23964
rect 12752 23962 12776 23964
rect 12832 23962 12856 23964
rect 12912 23962 12918 23964
rect 12672 23910 12674 23962
rect 12854 23910 12856 23962
rect 12610 23908 12616 23910
rect 12672 23908 12696 23910
rect 12752 23908 12776 23910
rect 12832 23908 12856 23910
rect 12912 23908 12918 23910
rect 12610 23899 12918 23908
rect 12610 22876 12918 22885
rect 12610 22874 12616 22876
rect 12672 22874 12696 22876
rect 12752 22874 12776 22876
rect 12832 22874 12856 22876
rect 12912 22874 12918 22876
rect 12672 22822 12674 22874
rect 12854 22822 12856 22874
rect 12610 22820 12616 22822
rect 12672 22820 12696 22822
rect 12752 22820 12776 22822
rect 12832 22820 12856 22822
rect 12912 22820 12918 22822
rect 12610 22811 12918 22820
rect 12610 21788 12918 21797
rect 12610 21786 12616 21788
rect 12672 21786 12696 21788
rect 12752 21786 12776 21788
rect 12832 21786 12856 21788
rect 12912 21786 12918 21788
rect 12672 21734 12674 21786
rect 12854 21734 12856 21786
rect 12610 21732 12616 21734
rect 12672 21732 12696 21734
rect 12752 21732 12776 21734
rect 12832 21732 12856 21734
rect 12912 21732 12918 21734
rect 12610 21723 12918 21732
rect 12440 21412 12492 21418
rect 12440 21354 12492 21360
rect 12992 21140 13044 21146
rect 12992 21082 13044 21088
rect 12610 20700 12918 20709
rect 12610 20698 12616 20700
rect 12672 20698 12696 20700
rect 12752 20698 12776 20700
rect 12832 20698 12856 20700
rect 12912 20698 12918 20700
rect 12672 20646 12674 20698
rect 12854 20646 12856 20698
rect 12610 20644 12616 20646
rect 12672 20644 12696 20646
rect 12752 20644 12776 20646
rect 12832 20644 12856 20646
rect 12912 20644 12918 20646
rect 12610 20635 12918 20644
rect 12610 19612 12918 19621
rect 12610 19610 12616 19612
rect 12672 19610 12696 19612
rect 12752 19610 12776 19612
rect 12832 19610 12856 19612
rect 12912 19610 12918 19612
rect 12672 19558 12674 19610
rect 12854 19558 12856 19610
rect 12610 19556 12616 19558
rect 12672 19556 12696 19558
rect 12752 19556 12776 19558
rect 12832 19556 12856 19558
rect 12912 19556 12918 19558
rect 12610 19547 12918 19556
rect 12610 18524 12918 18533
rect 12610 18522 12616 18524
rect 12672 18522 12696 18524
rect 12752 18522 12776 18524
rect 12832 18522 12856 18524
rect 12912 18522 12918 18524
rect 12672 18470 12674 18522
rect 12854 18470 12856 18522
rect 12610 18468 12616 18470
rect 12672 18468 12696 18470
rect 12752 18468 12776 18470
rect 12832 18468 12856 18470
rect 12912 18468 12918 18470
rect 12610 18459 12918 18468
rect 12610 17436 12918 17445
rect 12610 17434 12616 17436
rect 12672 17434 12696 17436
rect 12752 17434 12776 17436
rect 12832 17434 12856 17436
rect 12912 17434 12918 17436
rect 12672 17382 12674 17434
rect 12854 17382 12856 17434
rect 12610 17380 12616 17382
rect 12672 17380 12696 17382
rect 12752 17380 12776 17382
rect 12832 17380 12856 17382
rect 12912 17380 12918 17382
rect 12610 17371 12918 17380
rect 12610 16348 12918 16357
rect 12610 16346 12616 16348
rect 12672 16346 12696 16348
rect 12752 16346 12776 16348
rect 12832 16346 12856 16348
rect 12912 16346 12918 16348
rect 12672 16294 12674 16346
rect 12854 16294 12856 16346
rect 12610 16292 12616 16294
rect 12672 16292 12696 16294
rect 12752 16292 12776 16294
rect 12832 16292 12856 16294
rect 12912 16292 12918 16294
rect 12610 16283 12918 16292
rect 13004 15706 13032 21082
rect 12992 15700 13044 15706
rect 12992 15642 13044 15648
rect 13096 15434 13124 31726
rect 13188 30598 13216 53994
rect 13464 51066 13492 55150
rect 13452 51060 13504 51066
rect 13452 51002 13504 51008
rect 13268 50720 13320 50726
rect 13268 50662 13320 50668
rect 13280 40730 13308 50662
rect 13360 49700 13412 49706
rect 13360 49642 13412 49648
rect 13372 48822 13400 49642
rect 13360 48816 13412 48822
rect 13360 48758 13412 48764
rect 13544 48340 13596 48346
rect 13544 48282 13596 48288
rect 13556 41414 13584 48282
rect 13464 41386 13584 41414
rect 13268 40724 13320 40730
rect 13268 40666 13320 40672
rect 13464 39846 13492 41386
rect 13544 40384 13596 40390
rect 13544 40326 13596 40332
rect 13452 39840 13504 39846
rect 13452 39782 13504 39788
rect 13268 39432 13320 39438
rect 13268 39374 13320 39380
rect 13280 33930 13308 39374
rect 13556 35086 13584 40326
rect 13544 35080 13596 35086
rect 13544 35022 13596 35028
rect 13544 34604 13596 34610
rect 13544 34546 13596 34552
rect 13268 33924 13320 33930
rect 13268 33866 13320 33872
rect 13556 33522 13584 34546
rect 13544 33516 13596 33522
rect 13544 33458 13596 33464
rect 13556 33402 13584 33458
rect 13464 33374 13584 33402
rect 13176 30592 13228 30598
rect 13176 30534 13228 30540
rect 13176 19916 13228 19922
rect 13176 19858 13228 19864
rect 13188 15502 13216 19858
rect 13464 15706 13492 33374
rect 13544 33040 13596 33046
rect 13544 32982 13596 32988
rect 13452 15700 13504 15706
rect 13452 15642 13504 15648
rect 13176 15496 13228 15502
rect 13176 15438 13228 15444
rect 13084 15428 13136 15434
rect 13084 15370 13136 15376
rect 13268 15428 13320 15434
rect 13268 15370 13320 15376
rect 12610 15260 12918 15269
rect 12610 15258 12616 15260
rect 12672 15258 12696 15260
rect 12752 15258 12776 15260
rect 12832 15258 12856 15260
rect 12912 15258 12918 15260
rect 12672 15206 12674 15258
rect 12854 15206 12856 15258
rect 12610 15204 12616 15206
rect 12672 15204 12696 15206
rect 12752 15204 12776 15206
rect 12832 15204 12856 15206
rect 12912 15204 12918 15206
rect 12610 15195 12918 15204
rect 12610 14172 12918 14181
rect 12610 14170 12616 14172
rect 12672 14170 12696 14172
rect 12752 14170 12776 14172
rect 12832 14170 12856 14172
rect 12912 14170 12918 14172
rect 12672 14118 12674 14170
rect 12854 14118 12856 14170
rect 12610 14116 12616 14118
rect 12672 14116 12696 14118
rect 12752 14116 12776 14118
rect 12832 14116 12856 14118
rect 12912 14116 12918 14118
rect 12610 14107 12918 14116
rect 12610 13084 12918 13093
rect 12610 13082 12616 13084
rect 12672 13082 12696 13084
rect 12752 13082 12776 13084
rect 12832 13082 12856 13084
rect 12912 13082 12918 13084
rect 12672 13030 12674 13082
rect 12854 13030 12856 13082
rect 12610 13028 12616 13030
rect 12672 13028 12696 13030
rect 12752 13028 12776 13030
rect 12832 13028 12856 13030
rect 12912 13028 12918 13030
rect 12610 13019 12918 13028
rect 12610 11996 12918 12005
rect 12610 11994 12616 11996
rect 12672 11994 12696 11996
rect 12752 11994 12776 11996
rect 12832 11994 12856 11996
rect 12912 11994 12918 11996
rect 12672 11942 12674 11994
rect 12854 11942 12856 11994
rect 12610 11940 12616 11942
rect 12672 11940 12696 11942
rect 12752 11940 12776 11942
rect 12832 11940 12856 11942
rect 12912 11940 12918 11942
rect 12610 11931 12918 11940
rect 13280 11286 13308 15370
rect 13556 13870 13584 32982
rect 13544 13864 13596 13870
rect 13544 13806 13596 13812
rect 13268 11280 13320 11286
rect 13268 11222 13320 11228
rect 12610 10908 12918 10917
rect 12610 10906 12616 10908
rect 12672 10906 12696 10908
rect 12752 10906 12776 10908
rect 12832 10906 12856 10908
rect 12912 10906 12918 10908
rect 12672 10854 12674 10906
rect 12854 10854 12856 10906
rect 12610 10852 12616 10854
rect 12672 10852 12696 10854
rect 12752 10852 12776 10854
rect 12832 10852 12856 10854
rect 12912 10852 12918 10854
rect 12610 10843 12918 10852
rect 12348 10600 12400 10606
rect 12348 10542 12400 10548
rect 11950 10364 12258 10373
rect 11950 10362 11956 10364
rect 12012 10362 12036 10364
rect 12092 10362 12116 10364
rect 12172 10362 12196 10364
rect 12252 10362 12258 10364
rect 12012 10310 12014 10362
rect 12194 10310 12196 10362
rect 11950 10308 11956 10310
rect 12012 10308 12036 10310
rect 12092 10308 12116 10310
rect 12172 10308 12196 10310
rect 12252 10308 12258 10310
rect 11950 10299 12258 10308
rect 12610 9820 12918 9829
rect 12610 9818 12616 9820
rect 12672 9818 12696 9820
rect 12752 9818 12776 9820
rect 12832 9818 12856 9820
rect 12912 9818 12918 9820
rect 12672 9766 12674 9818
rect 12854 9766 12856 9818
rect 12610 9764 12616 9766
rect 12672 9764 12696 9766
rect 12752 9764 12776 9766
rect 12832 9764 12856 9766
rect 12912 9764 12918 9766
rect 12610 9755 12918 9764
rect 12992 9648 13044 9654
rect 12992 9590 13044 9596
rect 11950 9276 12258 9285
rect 11950 9274 11956 9276
rect 12012 9274 12036 9276
rect 12092 9274 12116 9276
rect 12172 9274 12196 9276
rect 12252 9274 12258 9276
rect 12012 9222 12014 9274
rect 12194 9222 12196 9274
rect 11950 9220 11956 9222
rect 12012 9220 12036 9222
rect 12092 9220 12116 9222
rect 12172 9220 12196 9222
rect 12252 9220 12258 9222
rect 11950 9211 12258 9220
rect 12610 8732 12918 8741
rect 12610 8730 12616 8732
rect 12672 8730 12696 8732
rect 12752 8730 12776 8732
rect 12832 8730 12856 8732
rect 12912 8730 12918 8732
rect 12672 8678 12674 8730
rect 12854 8678 12856 8730
rect 12610 8676 12616 8678
rect 12672 8676 12696 8678
rect 12752 8676 12776 8678
rect 12832 8676 12856 8678
rect 12912 8676 12918 8678
rect 12610 8667 12918 8676
rect 11950 8188 12258 8197
rect 11950 8186 11956 8188
rect 12012 8186 12036 8188
rect 12092 8186 12116 8188
rect 12172 8186 12196 8188
rect 12252 8186 12258 8188
rect 12012 8134 12014 8186
rect 12194 8134 12196 8186
rect 11950 8132 11956 8134
rect 12012 8132 12036 8134
rect 12092 8132 12116 8134
rect 12172 8132 12196 8134
rect 12252 8132 12258 8134
rect 11950 8123 12258 8132
rect 12610 7644 12918 7653
rect 12610 7642 12616 7644
rect 12672 7642 12696 7644
rect 12752 7642 12776 7644
rect 12832 7642 12856 7644
rect 12912 7642 12918 7644
rect 12672 7590 12674 7642
rect 12854 7590 12856 7642
rect 12610 7588 12616 7590
rect 12672 7588 12696 7590
rect 12752 7588 12776 7590
rect 12832 7588 12856 7590
rect 12912 7588 12918 7590
rect 12610 7579 12918 7588
rect 11950 7100 12258 7109
rect 11950 7098 11956 7100
rect 12012 7098 12036 7100
rect 12092 7098 12116 7100
rect 12172 7098 12196 7100
rect 12252 7098 12258 7100
rect 12012 7046 12014 7098
rect 12194 7046 12196 7098
rect 11950 7044 11956 7046
rect 12012 7044 12036 7046
rect 12092 7044 12116 7046
rect 12172 7044 12196 7046
rect 12252 7044 12258 7046
rect 11950 7035 12258 7044
rect 12610 6556 12918 6565
rect 12610 6554 12616 6556
rect 12672 6554 12696 6556
rect 12752 6554 12776 6556
rect 12832 6554 12856 6556
rect 12912 6554 12918 6556
rect 12672 6502 12674 6554
rect 12854 6502 12856 6554
rect 12610 6500 12616 6502
rect 12672 6500 12696 6502
rect 12752 6500 12776 6502
rect 12832 6500 12856 6502
rect 12912 6500 12918 6502
rect 12610 6491 12918 6500
rect 11950 6012 12258 6021
rect 11950 6010 11956 6012
rect 12012 6010 12036 6012
rect 12092 6010 12116 6012
rect 12172 6010 12196 6012
rect 12252 6010 12258 6012
rect 12012 5958 12014 6010
rect 12194 5958 12196 6010
rect 11950 5956 11956 5958
rect 12012 5956 12036 5958
rect 12092 5956 12116 5958
rect 12172 5956 12196 5958
rect 12252 5956 12258 5958
rect 11950 5947 12258 5956
rect 12610 5468 12918 5477
rect 12610 5466 12616 5468
rect 12672 5466 12696 5468
rect 12752 5466 12776 5468
rect 12832 5466 12856 5468
rect 12912 5466 12918 5468
rect 12672 5414 12674 5466
rect 12854 5414 12856 5466
rect 12610 5412 12616 5414
rect 12672 5412 12696 5414
rect 12752 5412 12776 5414
rect 12832 5412 12856 5414
rect 12912 5412 12918 5414
rect 12610 5403 12918 5412
rect 13004 5370 13032 9590
rect 13648 9586 13676 67798
rect 14556 65748 14608 65754
rect 14556 65690 14608 65696
rect 14004 64660 14056 64666
rect 14004 64602 14056 64608
rect 13912 62144 13964 62150
rect 13912 62086 13964 62092
rect 13820 61804 13872 61810
rect 13820 61746 13872 61752
rect 13728 61736 13780 61742
rect 13728 61678 13780 61684
rect 13740 55350 13768 61678
rect 13832 56166 13860 61746
rect 13924 61402 13952 62086
rect 13912 61396 13964 61402
rect 13912 61338 13964 61344
rect 14016 60734 14044 64602
rect 13924 60706 14044 60734
rect 13820 56160 13872 56166
rect 13820 56102 13872 56108
rect 13728 55344 13780 55350
rect 13728 55286 13780 55292
rect 13924 54210 13952 60706
rect 14372 58540 14424 58546
rect 14372 58482 14424 58488
rect 14004 58472 14056 58478
rect 14004 58414 14056 58420
rect 13832 54182 13952 54210
rect 13728 48612 13780 48618
rect 13728 48554 13780 48560
rect 13740 35086 13768 48554
rect 13832 35086 13860 54182
rect 13912 52488 13964 52494
rect 13912 52430 13964 52436
rect 13924 49842 13952 52430
rect 13912 49836 13964 49842
rect 13912 49778 13964 49784
rect 13728 35080 13780 35086
rect 13728 35022 13780 35028
rect 13820 35080 13872 35086
rect 13820 35022 13872 35028
rect 13728 34468 13780 34474
rect 13728 34410 13780 34416
rect 13740 33522 13768 34410
rect 13728 33516 13780 33522
rect 13728 33458 13780 33464
rect 13740 33046 13768 33458
rect 13728 33040 13780 33046
rect 13728 32982 13780 32988
rect 13820 32972 13872 32978
rect 13820 32914 13872 32920
rect 13832 9586 13860 32914
rect 13924 26994 13952 49778
rect 14016 42362 14044 58414
rect 14188 58404 14240 58410
rect 14188 58346 14240 58352
rect 14200 50454 14228 58346
rect 14384 54602 14412 58482
rect 14464 55344 14516 55350
rect 14464 55286 14516 55292
rect 14372 54596 14424 54602
rect 14372 54538 14424 54544
rect 14188 50448 14240 50454
rect 14188 50390 14240 50396
rect 14188 49836 14240 49842
rect 14188 49778 14240 49784
rect 14096 48136 14148 48142
rect 14096 48078 14148 48084
rect 14004 42356 14056 42362
rect 14004 42298 14056 42304
rect 14004 35148 14056 35154
rect 14004 35090 14056 35096
rect 14016 33318 14044 35090
rect 14004 33312 14056 33318
rect 14004 33254 14056 33260
rect 13912 26988 13964 26994
rect 13912 26930 13964 26936
rect 13636 9580 13688 9586
rect 13636 9522 13688 9528
rect 13820 9580 13872 9586
rect 13820 9522 13872 9528
rect 13648 7818 13676 9522
rect 13636 7812 13688 7818
rect 13636 7754 13688 7760
rect 12532 5364 12584 5370
rect 12532 5306 12584 5312
rect 12992 5364 13044 5370
rect 12992 5306 13044 5312
rect 11950 4924 12258 4933
rect 11950 4922 11956 4924
rect 12012 4922 12036 4924
rect 12092 4922 12116 4924
rect 12172 4922 12196 4924
rect 12252 4922 12258 4924
rect 12012 4870 12014 4922
rect 12194 4870 12196 4922
rect 11950 4868 11956 4870
rect 12012 4868 12036 4870
rect 12092 4868 12116 4870
rect 12172 4868 12196 4870
rect 12252 4868 12258 4870
rect 11950 4859 12258 4868
rect 11950 3836 12258 3845
rect 11950 3834 11956 3836
rect 12012 3834 12036 3836
rect 12092 3834 12116 3836
rect 12172 3834 12196 3836
rect 12252 3834 12258 3836
rect 12012 3782 12014 3834
rect 12194 3782 12196 3834
rect 11950 3780 11956 3782
rect 12012 3780 12036 3782
rect 12092 3780 12116 3782
rect 12172 3780 12196 3782
rect 12252 3780 12258 3782
rect 11950 3771 12258 3780
rect 12544 3534 12572 5306
rect 14108 4690 14136 48078
rect 14200 43450 14228 49778
rect 14476 47802 14504 55286
rect 14464 47796 14516 47802
rect 14464 47738 14516 47744
rect 14464 46572 14516 46578
rect 14464 46514 14516 46520
rect 14280 44192 14332 44198
rect 14280 44134 14332 44140
rect 14188 43444 14240 43450
rect 14188 43386 14240 43392
rect 14188 35692 14240 35698
rect 14188 35634 14240 35640
rect 14200 33522 14228 35634
rect 14188 33516 14240 33522
rect 14188 33458 14240 33464
rect 14292 33454 14320 44134
rect 14280 33448 14332 33454
rect 14280 33390 14332 33396
rect 14188 33108 14240 33114
rect 14188 33050 14240 33056
rect 14200 9654 14228 33050
rect 14280 22500 14332 22506
rect 14280 22442 14332 22448
rect 14188 9648 14240 9654
rect 14188 9590 14240 9596
rect 14096 4684 14148 4690
rect 14096 4626 14148 4632
rect 14292 4622 14320 22442
rect 14372 22432 14424 22438
rect 14372 22374 14424 22380
rect 14280 4616 14332 4622
rect 14280 4558 14332 4564
rect 12610 4380 12918 4389
rect 12610 4378 12616 4380
rect 12672 4378 12696 4380
rect 12752 4378 12776 4380
rect 12832 4378 12856 4380
rect 12912 4378 12918 4380
rect 12672 4326 12674 4378
rect 12854 4326 12856 4378
rect 12610 4324 12616 4326
rect 12672 4324 12696 4326
rect 12752 4324 12776 4326
rect 12832 4324 12856 4326
rect 12912 4324 12918 4326
rect 12610 4315 12918 4324
rect 12532 3528 12584 3534
rect 12532 3470 12584 3476
rect 12610 3292 12918 3301
rect 12610 3290 12616 3292
rect 12672 3290 12696 3292
rect 12752 3290 12776 3292
rect 12832 3290 12856 3292
rect 12912 3290 12918 3292
rect 12672 3238 12674 3290
rect 12854 3238 12856 3290
rect 12610 3236 12616 3238
rect 12672 3236 12696 3238
rect 12752 3236 12776 3238
rect 12832 3236 12856 3238
rect 12912 3236 12918 3238
rect 12610 3227 12918 3236
rect 11950 2748 12258 2757
rect 11950 2746 11956 2748
rect 12012 2746 12036 2748
rect 12092 2746 12116 2748
rect 12172 2746 12196 2748
rect 12252 2746 12258 2748
rect 12012 2694 12014 2746
rect 12194 2694 12196 2746
rect 11950 2692 11956 2694
rect 12012 2692 12036 2694
rect 12092 2692 12116 2694
rect 12172 2692 12196 2694
rect 12252 2692 12258 2694
rect 11950 2683 12258 2692
rect 14384 2582 14412 22374
rect 14476 3534 14504 46514
rect 14568 39642 14596 65690
rect 15108 64048 15160 64054
rect 15108 63990 15160 63996
rect 14648 62960 14700 62966
rect 14648 62902 14700 62908
rect 14660 55214 14688 62902
rect 15120 62354 15148 63990
rect 15108 62348 15160 62354
rect 15108 62290 15160 62296
rect 14648 55208 14700 55214
rect 14648 55150 14700 55156
rect 14924 53712 14976 53718
rect 14924 53654 14976 53660
rect 14936 53514 14964 53654
rect 14924 53508 14976 53514
rect 14924 53450 14976 53456
rect 14740 48000 14792 48006
rect 14740 47942 14792 47948
rect 14556 39636 14608 39642
rect 14556 39578 14608 39584
rect 14752 34202 14780 47942
rect 15016 39840 15068 39846
rect 15016 39782 15068 39788
rect 14924 39568 14976 39574
rect 14924 39510 14976 39516
rect 14832 38276 14884 38282
rect 14832 38218 14884 38224
rect 14844 35154 14872 38218
rect 14832 35148 14884 35154
rect 14832 35090 14884 35096
rect 14740 34196 14792 34202
rect 14740 34138 14792 34144
rect 14648 33312 14700 33318
rect 14648 33254 14700 33260
rect 14660 22642 14688 33254
rect 14752 31754 14780 34138
rect 14936 33998 14964 39510
rect 15028 35698 15056 39782
rect 15016 35692 15068 35698
rect 15016 35634 15068 35640
rect 14924 33992 14976 33998
rect 14924 33934 14976 33940
rect 14936 33658 14964 33934
rect 14832 33652 14884 33658
rect 14832 33594 14884 33600
rect 14924 33652 14976 33658
rect 14924 33594 14976 33600
rect 14844 33522 14872 33594
rect 14832 33516 14884 33522
rect 14832 33458 14884 33464
rect 14844 33318 14872 33458
rect 15016 33448 15068 33454
rect 15016 33390 15068 33396
rect 14832 33312 14884 33318
rect 14832 33254 14884 33260
rect 14752 31726 14872 31754
rect 14648 22636 14700 22642
rect 14648 22578 14700 22584
rect 14844 22030 14872 31726
rect 15028 30054 15056 33390
rect 15016 30048 15068 30054
rect 15016 29990 15068 29996
rect 15016 23180 15068 23186
rect 15016 23122 15068 23128
rect 14922 22808 14978 22817
rect 14922 22743 14978 22752
rect 14936 22710 14964 22743
rect 15028 22710 15056 23122
rect 14924 22704 14976 22710
rect 14924 22646 14976 22652
rect 15016 22704 15068 22710
rect 15016 22646 15068 22652
rect 14832 22024 14884 22030
rect 14832 21966 14884 21972
rect 14556 17536 14608 17542
rect 14556 17478 14608 17484
rect 14568 15094 14596 17478
rect 14556 15088 14608 15094
rect 14556 15030 14608 15036
rect 14568 12434 14596 15030
rect 14568 12406 14688 12434
rect 14660 8022 14688 12406
rect 15120 11150 15148 62290
rect 15476 54732 15528 54738
rect 15476 54674 15528 54680
rect 15292 54188 15344 54194
rect 15292 54130 15344 54136
rect 15304 53446 15332 54130
rect 15384 53712 15436 53718
rect 15384 53654 15436 53660
rect 15396 53582 15424 53654
rect 15384 53576 15436 53582
rect 15384 53518 15436 53524
rect 15292 53440 15344 53446
rect 15292 53382 15344 53388
rect 15292 53100 15344 53106
rect 15292 53042 15344 53048
rect 15200 52964 15252 52970
rect 15200 52906 15252 52912
rect 15212 35193 15240 52906
rect 15304 37942 15332 53042
rect 15396 52018 15424 53518
rect 15488 53514 15516 54674
rect 15476 53508 15528 53514
rect 15476 53450 15528 53456
rect 15580 53106 15608 68750
rect 20168 68672 20220 68678
rect 20168 68614 20220 68620
rect 17610 68572 17918 68581
rect 17610 68570 17616 68572
rect 17672 68570 17696 68572
rect 17752 68570 17776 68572
rect 17832 68570 17856 68572
rect 17912 68570 17918 68572
rect 17672 68518 17674 68570
rect 17854 68518 17856 68570
rect 17610 68516 17616 68518
rect 17672 68516 17696 68518
rect 17752 68516 17776 68518
rect 17832 68516 17856 68518
rect 17912 68516 17918 68518
rect 17610 68507 17918 68516
rect 19800 68332 19852 68338
rect 19800 68274 19852 68280
rect 16950 68028 17258 68037
rect 16950 68026 16956 68028
rect 17012 68026 17036 68028
rect 17092 68026 17116 68028
rect 17172 68026 17196 68028
rect 17252 68026 17258 68028
rect 17012 67974 17014 68026
rect 17194 67974 17196 68026
rect 16950 67972 16956 67974
rect 17012 67972 17036 67974
rect 17092 67972 17116 67974
rect 17172 67972 17196 67974
rect 17252 67972 17258 67974
rect 16950 67963 17258 67972
rect 17610 67484 17918 67493
rect 17610 67482 17616 67484
rect 17672 67482 17696 67484
rect 17752 67482 17776 67484
rect 17832 67482 17856 67484
rect 17912 67482 17918 67484
rect 17672 67430 17674 67482
rect 17854 67430 17856 67482
rect 17610 67428 17616 67430
rect 17672 67428 17696 67430
rect 17752 67428 17776 67430
rect 17832 67428 17856 67430
rect 17912 67428 17918 67430
rect 17610 67419 17918 67428
rect 18144 67312 18196 67318
rect 18144 67254 18196 67260
rect 16950 66940 17258 66949
rect 16950 66938 16956 66940
rect 17012 66938 17036 66940
rect 17092 66938 17116 66940
rect 17172 66938 17196 66940
rect 17252 66938 17258 66940
rect 17012 66886 17014 66938
rect 17194 66886 17196 66938
rect 16950 66884 16956 66886
rect 17012 66884 17036 66886
rect 17092 66884 17116 66886
rect 17172 66884 17196 66886
rect 17252 66884 17258 66886
rect 16950 66875 17258 66884
rect 17610 66396 17918 66405
rect 17610 66394 17616 66396
rect 17672 66394 17696 66396
rect 17752 66394 17776 66396
rect 17832 66394 17856 66396
rect 17912 66394 17918 66396
rect 17672 66342 17674 66394
rect 17854 66342 17856 66394
rect 17610 66340 17616 66342
rect 17672 66340 17696 66342
rect 17752 66340 17776 66342
rect 17832 66340 17856 66342
rect 17912 66340 17918 66342
rect 17610 66331 17918 66340
rect 16950 65852 17258 65861
rect 16950 65850 16956 65852
rect 17012 65850 17036 65852
rect 17092 65850 17116 65852
rect 17172 65850 17196 65852
rect 17252 65850 17258 65852
rect 17012 65798 17014 65850
rect 17194 65798 17196 65850
rect 16950 65796 16956 65798
rect 17012 65796 17036 65798
rect 17092 65796 17116 65798
rect 17172 65796 17196 65798
rect 17252 65796 17258 65798
rect 16950 65787 17258 65796
rect 17610 65308 17918 65317
rect 17610 65306 17616 65308
rect 17672 65306 17696 65308
rect 17752 65306 17776 65308
rect 17832 65306 17856 65308
rect 17912 65306 17918 65308
rect 17672 65254 17674 65306
rect 17854 65254 17856 65306
rect 17610 65252 17616 65254
rect 17672 65252 17696 65254
rect 17752 65252 17776 65254
rect 17832 65252 17856 65254
rect 17912 65252 17918 65254
rect 17610 65243 17918 65252
rect 16396 65204 16448 65210
rect 16396 65146 16448 65152
rect 16408 63578 16436 65146
rect 16950 64764 17258 64773
rect 16950 64762 16956 64764
rect 17012 64762 17036 64764
rect 17092 64762 17116 64764
rect 17172 64762 17196 64764
rect 17252 64762 17258 64764
rect 17012 64710 17014 64762
rect 17194 64710 17196 64762
rect 16950 64708 16956 64710
rect 17012 64708 17036 64710
rect 17092 64708 17116 64710
rect 17172 64708 17196 64710
rect 17252 64708 17258 64710
rect 16950 64699 17258 64708
rect 17316 64388 17368 64394
rect 17316 64330 17368 64336
rect 16950 63676 17258 63685
rect 16950 63674 16956 63676
rect 17012 63674 17036 63676
rect 17092 63674 17116 63676
rect 17172 63674 17196 63676
rect 17252 63674 17258 63676
rect 17012 63622 17014 63674
rect 17194 63622 17196 63674
rect 16950 63620 16956 63622
rect 17012 63620 17036 63622
rect 17092 63620 17116 63622
rect 17172 63620 17196 63622
rect 17252 63620 17258 63622
rect 16950 63611 17258 63620
rect 16396 63572 16448 63578
rect 16396 63514 16448 63520
rect 16304 63028 16356 63034
rect 16304 62970 16356 62976
rect 16120 57316 16172 57322
rect 16120 57258 16172 57264
rect 15936 55888 15988 55894
rect 15936 55830 15988 55836
rect 15948 54058 15976 55830
rect 15936 54052 15988 54058
rect 15936 53994 15988 54000
rect 15844 53508 15896 53514
rect 15844 53450 15896 53456
rect 15568 53100 15620 53106
rect 15568 53042 15620 53048
rect 15384 52012 15436 52018
rect 15384 51954 15436 51960
rect 15568 41608 15620 41614
rect 15568 41550 15620 41556
rect 15292 37936 15344 37942
rect 15292 37878 15344 37884
rect 15292 36576 15344 36582
rect 15292 36518 15344 36524
rect 15198 35184 15254 35193
rect 15198 35119 15254 35128
rect 15212 26314 15240 35119
rect 15200 26308 15252 26314
rect 15200 26250 15252 26256
rect 15304 22098 15332 36518
rect 15580 34610 15608 41550
rect 15568 34604 15620 34610
rect 15568 34546 15620 34552
rect 15752 34604 15804 34610
rect 15752 34546 15804 34552
rect 15660 33992 15712 33998
rect 15660 33934 15712 33940
rect 15672 31754 15700 33934
rect 15764 33386 15792 34546
rect 15752 33380 15804 33386
rect 15752 33322 15804 33328
rect 15580 31726 15700 31754
rect 15292 22092 15344 22098
rect 15580 22094 15608 31726
rect 15856 29594 15884 53450
rect 15936 53032 15988 53038
rect 15936 52974 15988 52980
rect 15948 33046 15976 52974
rect 16132 33862 16160 57258
rect 16316 56846 16344 62970
rect 16304 56840 16356 56846
rect 16304 56782 16356 56788
rect 16316 55622 16344 56782
rect 16304 55616 16356 55622
rect 16304 55558 16356 55564
rect 16212 53100 16264 53106
rect 16212 53042 16264 53048
rect 16120 33856 16172 33862
rect 16120 33798 16172 33804
rect 15936 33040 15988 33046
rect 15936 32982 15988 32988
rect 16028 32564 16080 32570
rect 16028 32506 16080 32512
rect 15936 31136 15988 31142
rect 15936 31078 15988 31084
rect 15672 29566 15884 29594
rect 15672 25702 15700 29566
rect 15844 29504 15896 29510
rect 15844 29446 15896 29452
rect 15660 25696 15712 25702
rect 15660 25638 15712 25644
rect 15856 22094 15884 29446
rect 15948 28558 15976 31078
rect 15936 28552 15988 28558
rect 15936 28494 15988 28500
rect 15948 25430 15976 28494
rect 15936 25424 15988 25430
rect 15936 25366 15988 25372
rect 15580 22066 15792 22094
rect 15856 22066 15976 22094
rect 15292 22034 15344 22040
rect 15764 19854 15792 22066
rect 15948 21078 15976 22066
rect 15936 21072 15988 21078
rect 15936 21014 15988 21020
rect 15752 19848 15804 19854
rect 15752 19790 15804 19796
rect 15108 11144 15160 11150
rect 15108 11086 15160 11092
rect 15660 9512 15712 9518
rect 15660 9454 15712 9460
rect 14648 8016 14700 8022
rect 14648 7958 14700 7964
rect 15672 7886 15700 9454
rect 15660 7880 15712 7886
rect 15660 7822 15712 7828
rect 15764 7410 15792 19790
rect 16040 9518 16068 32506
rect 16132 30938 16160 33798
rect 16120 30932 16172 30938
rect 16120 30874 16172 30880
rect 16224 30818 16252 53042
rect 16316 39506 16344 55558
rect 16408 51074 16436 63514
rect 16580 62824 16632 62830
rect 16580 62766 16632 62772
rect 16488 55616 16540 55622
rect 16488 55558 16540 55564
rect 16500 55321 16528 55558
rect 16486 55312 16542 55321
rect 16486 55247 16542 55256
rect 16408 51046 16528 51074
rect 16500 41614 16528 51046
rect 16592 48890 16620 62766
rect 16950 62588 17258 62597
rect 16950 62586 16956 62588
rect 17012 62586 17036 62588
rect 17092 62586 17116 62588
rect 17172 62586 17196 62588
rect 17252 62586 17258 62588
rect 17012 62534 17014 62586
rect 17194 62534 17196 62586
rect 16950 62532 16956 62534
rect 17012 62532 17036 62534
rect 17092 62532 17116 62534
rect 17172 62532 17196 62534
rect 17252 62532 17258 62534
rect 16950 62523 17258 62532
rect 16950 61500 17258 61509
rect 16950 61498 16956 61500
rect 17012 61498 17036 61500
rect 17092 61498 17116 61500
rect 17172 61498 17196 61500
rect 17252 61498 17258 61500
rect 17012 61446 17014 61498
rect 17194 61446 17196 61498
rect 16950 61444 16956 61446
rect 17012 61444 17036 61446
rect 17092 61444 17116 61446
rect 17172 61444 17196 61446
rect 17252 61444 17258 61446
rect 16950 61435 17258 61444
rect 16950 60412 17258 60421
rect 16950 60410 16956 60412
rect 17012 60410 17036 60412
rect 17092 60410 17116 60412
rect 17172 60410 17196 60412
rect 17252 60410 17258 60412
rect 17012 60358 17014 60410
rect 17194 60358 17196 60410
rect 16950 60356 16956 60358
rect 17012 60356 17036 60358
rect 17092 60356 17116 60358
rect 17172 60356 17196 60358
rect 17252 60356 17258 60358
rect 16950 60347 17258 60356
rect 16950 59324 17258 59333
rect 16950 59322 16956 59324
rect 17012 59322 17036 59324
rect 17092 59322 17116 59324
rect 17172 59322 17196 59324
rect 17252 59322 17258 59324
rect 17012 59270 17014 59322
rect 17194 59270 17196 59322
rect 16950 59268 16956 59270
rect 17012 59268 17036 59270
rect 17092 59268 17116 59270
rect 17172 59268 17196 59270
rect 17252 59268 17258 59270
rect 16950 59259 17258 59268
rect 16950 58236 17258 58245
rect 16950 58234 16956 58236
rect 17012 58234 17036 58236
rect 17092 58234 17116 58236
rect 17172 58234 17196 58236
rect 17252 58234 17258 58236
rect 17012 58182 17014 58234
rect 17194 58182 17196 58234
rect 16950 58180 16956 58182
rect 17012 58180 17036 58182
rect 17092 58180 17116 58182
rect 17172 58180 17196 58182
rect 17252 58180 17258 58182
rect 16950 58171 17258 58180
rect 16856 57452 16908 57458
rect 16856 57394 16908 57400
rect 16672 57384 16724 57390
rect 16672 57326 16724 57332
rect 16580 48884 16632 48890
rect 16580 48826 16632 48832
rect 16580 43240 16632 43246
rect 16580 43182 16632 43188
rect 16488 41608 16540 41614
rect 16488 41550 16540 41556
rect 16592 41414 16620 43182
rect 16500 41386 16620 41414
rect 16500 40186 16528 41386
rect 16580 41268 16632 41274
rect 16580 41210 16632 41216
rect 16488 40180 16540 40186
rect 16488 40122 16540 40128
rect 16304 39500 16356 39506
rect 16304 39442 16356 39448
rect 16316 39098 16344 39442
rect 16304 39092 16356 39098
rect 16304 39034 16356 39040
rect 16592 35986 16620 41210
rect 16500 35958 16620 35986
rect 16500 35630 16528 35958
rect 16684 35850 16712 57326
rect 16868 52154 16896 57394
rect 16950 57148 17258 57157
rect 16950 57146 16956 57148
rect 17012 57146 17036 57148
rect 17092 57146 17116 57148
rect 17172 57146 17196 57148
rect 17252 57146 17258 57148
rect 17012 57094 17014 57146
rect 17194 57094 17196 57146
rect 16950 57092 16956 57094
rect 17012 57092 17036 57094
rect 17092 57092 17116 57094
rect 17172 57092 17196 57094
rect 17252 57092 17258 57094
rect 16950 57083 17258 57092
rect 16950 56060 17258 56069
rect 16950 56058 16956 56060
rect 17012 56058 17036 56060
rect 17092 56058 17116 56060
rect 17172 56058 17196 56060
rect 17252 56058 17258 56060
rect 17012 56006 17014 56058
rect 17194 56006 17196 56058
rect 16950 56004 16956 56006
rect 17012 56004 17036 56006
rect 17092 56004 17116 56006
rect 17172 56004 17196 56006
rect 17252 56004 17258 56006
rect 16950 55995 17258 56004
rect 16950 54972 17258 54981
rect 16950 54970 16956 54972
rect 17012 54970 17036 54972
rect 17092 54970 17116 54972
rect 17172 54970 17196 54972
rect 17252 54970 17258 54972
rect 17012 54918 17014 54970
rect 17194 54918 17196 54970
rect 16950 54916 16956 54918
rect 17012 54916 17036 54918
rect 17092 54916 17116 54918
rect 17172 54916 17196 54918
rect 17252 54916 17258 54918
rect 16950 54907 17258 54916
rect 16950 53884 17258 53893
rect 16950 53882 16956 53884
rect 17012 53882 17036 53884
rect 17092 53882 17116 53884
rect 17172 53882 17196 53884
rect 17252 53882 17258 53884
rect 17012 53830 17014 53882
rect 17194 53830 17196 53882
rect 16950 53828 16956 53830
rect 17012 53828 17036 53830
rect 17092 53828 17116 53830
rect 17172 53828 17196 53830
rect 17252 53828 17258 53830
rect 16950 53819 17258 53828
rect 16950 52796 17258 52805
rect 16950 52794 16956 52796
rect 17012 52794 17036 52796
rect 17092 52794 17116 52796
rect 17172 52794 17196 52796
rect 17252 52794 17258 52796
rect 17012 52742 17014 52794
rect 17194 52742 17196 52794
rect 16950 52740 16956 52742
rect 17012 52740 17036 52742
rect 17092 52740 17116 52742
rect 17172 52740 17196 52742
rect 17252 52740 17258 52742
rect 16950 52731 17258 52740
rect 16856 52148 16908 52154
rect 16856 52090 16908 52096
rect 16764 48544 16816 48550
rect 16764 48486 16816 48492
rect 16776 43246 16804 48486
rect 16764 43240 16816 43246
rect 16764 43182 16816 43188
rect 16764 43104 16816 43110
rect 16764 43046 16816 43052
rect 16776 40526 16804 43046
rect 16764 40520 16816 40526
rect 16764 40462 16816 40468
rect 16764 40180 16816 40186
rect 16764 40122 16816 40128
rect 16776 37126 16804 40122
rect 16868 37874 16896 52090
rect 16950 51708 17258 51717
rect 16950 51706 16956 51708
rect 17012 51706 17036 51708
rect 17092 51706 17116 51708
rect 17172 51706 17196 51708
rect 17252 51706 17258 51708
rect 17012 51654 17014 51706
rect 17194 51654 17196 51706
rect 16950 51652 16956 51654
rect 17012 51652 17036 51654
rect 17092 51652 17116 51654
rect 17172 51652 17196 51654
rect 17252 51652 17258 51654
rect 16950 51643 17258 51652
rect 16950 50620 17258 50629
rect 16950 50618 16956 50620
rect 17012 50618 17036 50620
rect 17092 50618 17116 50620
rect 17172 50618 17196 50620
rect 17252 50618 17258 50620
rect 17012 50566 17014 50618
rect 17194 50566 17196 50618
rect 16950 50564 16956 50566
rect 17012 50564 17036 50566
rect 17092 50564 17116 50566
rect 17172 50564 17196 50566
rect 17252 50564 17258 50566
rect 16950 50555 17258 50564
rect 16950 49532 17258 49541
rect 16950 49530 16956 49532
rect 17012 49530 17036 49532
rect 17092 49530 17116 49532
rect 17172 49530 17196 49532
rect 17252 49530 17258 49532
rect 17012 49478 17014 49530
rect 17194 49478 17196 49530
rect 16950 49476 16956 49478
rect 17012 49476 17036 49478
rect 17092 49476 17116 49478
rect 17172 49476 17196 49478
rect 17252 49476 17258 49478
rect 16950 49467 17258 49476
rect 17328 48754 17356 64330
rect 17610 64220 17918 64229
rect 17610 64218 17616 64220
rect 17672 64218 17696 64220
rect 17752 64218 17776 64220
rect 17832 64218 17856 64220
rect 17912 64218 17918 64220
rect 17672 64166 17674 64218
rect 17854 64166 17856 64218
rect 17610 64164 17616 64166
rect 17672 64164 17696 64166
rect 17752 64164 17776 64166
rect 17832 64164 17856 64166
rect 17912 64164 17918 64166
rect 17610 64155 17918 64164
rect 17960 63232 18012 63238
rect 17960 63174 18012 63180
rect 17610 63132 17918 63141
rect 17610 63130 17616 63132
rect 17672 63130 17696 63132
rect 17752 63130 17776 63132
rect 17832 63130 17856 63132
rect 17912 63130 17918 63132
rect 17672 63078 17674 63130
rect 17854 63078 17856 63130
rect 17610 63076 17616 63078
rect 17672 63076 17696 63078
rect 17752 63076 17776 63078
rect 17832 63076 17856 63078
rect 17912 63076 17918 63078
rect 17610 63067 17918 63076
rect 17972 62694 18000 63174
rect 17960 62688 18012 62694
rect 17960 62630 18012 62636
rect 17972 62150 18000 62630
rect 18156 62422 18184 67254
rect 18604 67244 18656 67250
rect 18604 67186 18656 67192
rect 18236 67176 18288 67182
rect 18236 67118 18288 67124
rect 18144 62416 18196 62422
rect 18144 62358 18196 62364
rect 18248 62354 18276 67118
rect 18328 67108 18380 67114
rect 18328 67050 18380 67056
rect 18236 62348 18288 62354
rect 18236 62290 18288 62296
rect 17960 62144 18012 62150
rect 17960 62086 18012 62092
rect 17610 62044 17918 62053
rect 17610 62042 17616 62044
rect 17672 62042 17696 62044
rect 17752 62042 17776 62044
rect 17832 62042 17856 62044
rect 17912 62042 17918 62044
rect 17672 61990 17674 62042
rect 17854 61990 17856 62042
rect 17610 61988 17616 61990
rect 17672 61988 17696 61990
rect 17752 61988 17776 61990
rect 17832 61988 17856 61990
rect 17912 61988 17918 61990
rect 17610 61979 17918 61988
rect 17972 61606 18000 62086
rect 17960 61600 18012 61606
rect 17960 61542 18012 61548
rect 17960 61260 18012 61266
rect 17960 61202 18012 61208
rect 17610 60956 17918 60965
rect 17610 60954 17616 60956
rect 17672 60954 17696 60956
rect 17752 60954 17776 60956
rect 17832 60954 17856 60956
rect 17912 60954 17918 60956
rect 17672 60902 17674 60954
rect 17854 60902 17856 60954
rect 17610 60900 17616 60902
rect 17672 60900 17696 60902
rect 17752 60900 17776 60902
rect 17832 60900 17856 60902
rect 17912 60900 17918 60902
rect 17610 60891 17918 60900
rect 17610 59868 17918 59877
rect 17610 59866 17616 59868
rect 17672 59866 17696 59868
rect 17752 59866 17776 59868
rect 17832 59866 17856 59868
rect 17912 59866 17918 59868
rect 17672 59814 17674 59866
rect 17854 59814 17856 59866
rect 17610 59812 17616 59814
rect 17672 59812 17696 59814
rect 17752 59812 17776 59814
rect 17832 59812 17856 59814
rect 17912 59812 17918 59814
rect 17610 59803 17918 59812
rect 17610 58780 17918 58789
rect 17610 58778 17616 58780
rect 17672 58778 17696 58780
rect 17752 58778 17776 58780
rect 17832 58778 17856 58780
rect 17912 58778 17918 58780
rect 17672 58726 17674 58778
rect 17854 58726 17856 58778
rect 17610 58724 17616 58726
rect 17672 58724 17696 58726
rect 17752 58724 17776 58726
rect 17832 58724 17856 58726
rect 17912 58724 17918 58726
rect 17610 58715 17918 58724
rect 17610 57692 17918 57701
rect 17610 57690 17616 57692
rect 17672 57690 17696 57692
rect 17752 57690 17776 57692
rect 17832 57690 17856 57692
rect 17912 57690 17918 57692
rect 17672 57638 17674 57690
rect 17854 57638 17856 57690
rect 17610 57636 17616 57638
rect 17672 57636 17696 57638
rect 17752 57636 17776 57638
rect 17832 57636 17856 57638
rect 17912 57636 17918 57638
rect 17610 57627 17918 57636
rect 17610 56604 17918 56613
rect 17610 56602 17616 56604
rect 17672 56602 17696 56604
rect 17752 56602 17776 56604
rect 17832 56602 17856 56604
rect 17912 56602 17918 56604
rect 17672 56550 17674 56602
rect 17854 56550 17856 56602
rect 17610 56548 17616 56550
rect 17672 56548 17696 56550
rect 17752 56548 17776 56550
rect 17832 56548 17856 56550
rect 17912 56548 17918 56550
rect 17610 56539 17918 56548
rect 17972 55758 18000 61202
rect 17960 55752 18012 55758
rect 17960 55694 18012 55700
rect 17610 55516 17918 55525
rect 17610 55514 17616 55516
rect 17672 55514 17696 55516
rect 17752 55514 17776 55516
rect 17832 55514 17856 55516
rect 17912 55514 17918 55516
rect 17672 55462 17674 55514
rect 17854 55462 17856 55514
rect 17610 55460 17616 55462
rect 17672 55460 17696 55462
rect 17752 55460 17776 55462
rect 17832 55460 17856 55462
rect 17912 55460 17918 55462
rect 17610 55451 17918 55460
rect 17610 54428 17918 54437
rect 17610 54426 17616 54428
rect 17672 54426 17696 54428
rect 17752 54426 17776 54428
rect 17832 54426 17856 54428
rect 17912 54426 17918 54428
rect 17672 54374 17674 54426
rect 17854 54374 17856 54426
rect 17610 54372 17616 54374
rect 17672 54372 17696 54374
rect 17752 54372 17776 54374
rect 17832 54372 17856 54374
rect 17912 54372 17918 54374
rect 17610 54363 17918 54372
rect 17610 53340 17918 53349
rect 17610 53338 17616 53340
rect 17672 53338 17696 53340
rect 17752 53338 17776 53340
rect 17832 53338 17856 53340
rect 17912 53338 17918 53340
rect 17672 53286 17674 53338
rect 17854 53286 17856 53338
rect 17610 53284 17616 53286
rect 17672 53284 17696 53286
rect 17752 53284 17776 53286
rect 17832 53284 17856 53286
rect 17912 53284 17918 53286
rect 17610 53275 17918 53284
rect 17610 52252 17918 52261
rect 17610 52250 17616 52252
rect 17672 52250 17696 52252
rect 17752 52250 17776 52252
rect 17832 52250 17856 52252
rect 17912 52250 17918 52252
rect 17672 52198 17674 52250
rect 17854 52198 17856 52250
rect 17610 52196 17616 52198
rect 17672 52196 17696 52198
rect 17752 52196 17776 52198
rect 17832 52196 17856 52198
rect 17912 52196 17918 52198
rect 17610 52187 17918 52196
rect 18144 51944 18196 51950
rect 18144 51886 18196 51892
rect 17610 51164 17918 51173
rect 17610 51162 17616 51164
rect 17672 51162 17696 51164
rect 17752 51162 17776 51164
rect 17832 51162 17856 51164
rect 17912 51162 17918 51164
rect 17672 51110 17674 51162
rect 17854 51110 17856 51162
rect 17610 51108 17616 51110
rect 17672 51108 17696 51110
rect 17752 51108 17776 51110
rect 17832 51108 17856 51110
rect 17912 51108 17918 51110
rect 17610 51099 17918 51108
rect 17500 50856 17552 50862
rect 17500 50798 17552 50804
rect 17316 48748 17368 48754
rect 17316 48690 17368 48696
rect 16948 48680 17000 48686
rect 16948 48622 17000 48628
rect 16960 48550 16988 48622
rect 16948 48544 17000 48550
rect 16948 48486 17000 48492
rect 16950 48444 17258 48453
rect 16950 48442 16956 48444
rect 17012 48442 17036 48444
rect 17092 48442 17116 48444
rect 17172 48442 17196 48444
rect 17252 48442 17258 48444
rect 17012 48390 17014 48442
rect 17194 48390 17196 48442
rect 16950 48388 16956 48390
rect 17012 48388 17036 48390
rect 17092 48388 17116 48390
rect 17172 48388 17196 48390
rect 17252 48388 17258 48390
rect 16950 48379 17258 48388
rect 16950 47356 17258 47365
rect 16950 47354 16956 47356
rect 17012 47354 17036 47356
rect 17092 47354 17116 47356
rect 17172 47354 17196 47356
rect 17252 47354 17258 47356
rect 17012 47302 17014 47354
rect 17194 47302 17196 47354
rect 16950 47300 16956 47302
rect 17012 47300 17036 47302
rect 17092 47300 17116 47302
rect 17172 47300 17196 47302
rect 17252 47300 17258 47302
rect 16950 47291 17258 47300
rect 16950 46268 17258 46277
rect 16950 46266 16956 46268
rect 17012 46266 17036 46268
rect 17092 46266 17116 46268
rect 17172 46266 17196 46268
rect 17252 46266 17258 46268
rect 17012 46214 17014 46266
rect 17194 46214 17196 46266
rect 16950 46212 16956 46214
rect 17012 46212 17036 46214
rect 17092 46212 17116 46214
rect 17172 46212 17196 46214
rect 17252 46212 17258 46214
rect 16950 46203 17258 46212
rect 16950 45180 17258 45189
rect 16950 45178 16956 45180
rect 17012 45178 17036 45180
rect 17092 45178 17116 45180
rect 17172 45178 17196 45180
rect 17252 45178 17258 45180
rect 17012 45126 17014 45178
rect 17194 45126 17196 45178
rect 16950 45124 16956 45126
rect 17012 45124 17036 45126
rect 17092 45124 17116 45126
rect 17172 45124 17196 45126
rect 17252 45124 17258 45126
rect 16950 45115 17258 45124
rect 16950 44092 17258 44101
rect 16950 44090 16956 44092
rect 17012 44090 17036 44092
rect 17092 44090 17116 44092
rect 17172 44090 17196 44092
rect 17252 44090 17258 44092
rect 17012 44038 17014 44090
rect 17194 44038 17196 44090
rect 16950 44036 16956 44038
rect 17012 44036 17036 44038
rect 17092 44036 17116 44038
rect 17172 44036 17196 44038
rect 17252 44036 17258 44038
rect 16950 44027 17258 44036
rect 16950 43004 17258 43013
rect 16950 43002 16956 43004
rect 17012 43002 17036 43004
rect 17092 43002 17116 43004
rect 17172 43002 17196 43004
rect 17252 43002 17258 43004
rect 17012 42950 17014 43002
rect 17194 42950 17196 43002
rect 16950 42948 16956 42950
rect 17012 42948 17036 42950
rect 17092 42948 17116 42950
rect 17172 42948 17196 42950
rect 17252 42948 17258 42950
rect 16950 42939 17258 42948
rect 16950 41916 17258 41925
rect 16950 41914 16956 41916
rect 17012 41914 17036 41916
rect 17092 41914 17116 41916
rect 17172 41914 17196 41916
rect 17252 41914 17258 41916
rect 17012 41862 17014 41914
rect 17194 41862 17196 41914
rect 16950 41860 16956 41862
rect 17012 41860 17036 41862
rect 17092 41860 17116 41862
rect 17172 41860 17196 41862
rect 17252 41860 17258 41862
rect 16950 41851 17258 41860
rect 17328 41274 17356 48690
rect 17408 48680 17460 48686
rect 17408 48622 17460 48628
rect 17316 41268 17368 41274
rect 17316 41210 17368 41216
rect 17316 41132 17368 41138
rect 17316 41074 17368 41080
rect 16950 40828 17258 40837
rect 16950 40826 16956 40828
rect 17012 40826 17036 40828
rect 17092 40826 17116 40828
rect 17172 40826 17196 40828
rect 17252 40826 17258 40828
rect 17012 40774 17014 40826
rect 17194 40774 17196 40826
rect 16950 40772 16956 40774
rect 17012 40772 17036 40774
rect 17092 40772 17116 40774
rect 17172 40772 17196 40774
rect 17252 40772 17258 40774
rect 16950 40763 17258 40772
rect 17328 40118 17356 41074
rect 17316 40112 17368 40118
rect 17316 40054 17368 40060
rect 16950 39740 17258 39749
rect 16950 39738 16956 39740
rect 17012 39738 17036 39740
rect 17092 39738 17116 39740
rect 17172 39738 17196 39740
rect 17252 39738 17258 39740
rect 17012 39686 17014 39738
rect 17194 39686 17196 39738
rect 16950 39684 16956 39686
rect 17012 39684 17036 39686
rect 17092 39684 17116 39686
rect 17172 39684 17196 39686
rect 17252 39684 17258 39686
rect 16950 39675 17258 39684
rect 16950 38652 17258 38661
rect 16950 38650 16956 38652
rect 17012 38650 17036 38652
rect 17092 38650 17116 38652
rect 17172 38650 17196 38652
rect 17252 38650 17258 38652
rect 17012 38598 17014 38650
rect 17194 38598 17196 38650
rect 16950 38596 16956 38598
rect 17012 38596 17036 38598
rect 17092 38596 17116 38598
rect 17172 38596 17196 38598
rect 17252 38596 17258 38598
rect 16950 38587 17258 38596
rect 17420 38162 17448 48622
rect 17328 38134 17448 38162
rect 16856 37868 16908 37874
rect 16856 37810 16908 37816
rect 16950 37564 17258 37573
rect 16950 37562 16956 37564
rect 17012 37562 17036 37564
rect 17092 37562 17116 37564
rect 17172 37562 17196 37564
rect 17252 37562 17258 37564
rect 17012 37510 17014 37562
rect 17194 37510 17196 37562
rect 16950 37508 16956 37510
rect 17012 37508 17036 37510
rect 17092 37508 17116 37510
rect 17172 37508 17196 37510
rect 17252 37508 17258 37510
rect 16950 37499 17258 37508
rect 16764 37120 16816 37126
rect 16764 37062 16816 37068
rect 16592 35822 16712 35850
rect 16488 35624 16540 35630
rect 16488 35566 16540 35572
rect 16396 35556 16448 35562
rect 16396 35498 16448 35504
rect 16408 35154 16436 35498
rect 16396 35148 16448 35154
rect 16396 35090 16448 35096
rect 16396 31952 16448 31958
rect 16592 31906 16620 35822
rect 16672 35760 16724 35766
rect 16672 35702 16724 35708
rect 16684 35154 16712 35702
rect 16672 35148 16724 35154
rect 16672 35090 16724 35096
rect 16672 34536 16724 34542
rect 16672 34478 16724 34484
rect 16396 31894 16448 31900
rect 16408 31226 16436 31894
rect 16500 31878 16620 31906
rect 16500 31362 16528 31878
rect 16684 31482 16712 34478
rect 16776 31958 16804 37062
rect 16950 36476 17258 36485
rect 16950 36474 16956 36476
rect 17012 36474 17036 36476
rect 17092 36474 17116 36476
rect 17172 36474 17196 36476
rect 17252 36474 17258 36476
rect 17012 36422 17014 36474
rect 17194 36422 17196 36474
rect 16950 36420 16956 36422
rect 17012 36420 17036 36422
rect 17092 36420 17116 36422
rect 17172 36420 17196 36422
rect 17252 36420 17258 36422
rect 16950 36411 17258 36420
rect 17328 36258 17356 38134
rect 17408 37324 17460 37330
rect 17408 37266 17460 37272
rect 17236 36230 17356 36258
rect 17236 35698 17264 36230
rect 17224 35692 17276 35698
rect 17224 35634 17276 35640
rect 16856 35624 16908 35630
rect 16856 35566 16908 35572
rect 16868 34678 16896 35566
rect 16950 35388 17258 35397
rect 16950 35386 16956 35388
rect 17012 35386 17036 35388
rect 17092 35386 17116 35388
rect 17172 35386 17196 35388
rect 17252 35386 17258 35388
rect 17012 35334 17014 35386
rect 17194 35334 17196 35386
rect 16950 35332 16956 35334
rect 17012 35332 17036 35334
rect 17092 35332 17116 35334
rect 17172 35332 17196 35334
rect 17252 35332 17258 35334
rect 16950 35323 17258 35332
rect 16856 34672 16908 34678
rect 16856 34614 16908 34620
rect 16950 34300 17258 34309
rect 16950 34298 16956 34300
rect 17012 34298 17036 34300
rect 17092 34298 17116 34300
rect 17172 34298 17196 34300
rect 17252 34298 17258 34300
rect 17012 34246 17014 34298
rect 17194 34246 17196 34298
rect 16950 34244 16956 34246
rect 17012 34244 17036 34246
rect 17092 34244 17116 34246
rect 17172 34244 17196 34246
rect 17252 34244 17258 34246
rect 16950 34235 17258 34244
rect 17316 33924 17368 33930
rect 17316 33866 17368 33872
rect 17328 33590 17356 33866
rect 17316 33584 17368 33590
rect 17316 33526 17368 33532
rect 17420 33538 17448 37266
rect 17512 33658 17540 50798
rect 17610 50076 17918 50085
rect 17610 50074 17616 50076
rect 17672 50074 17696 50076
rect 17752 50074 17776 50076
rect 17832 50074 17856 50076
rect 17912 50074 17918 50076
rect 17672 50022 17674 50074
rect 17854 50022 17856 50074
rect 17610 50020 17616 50022
rect 17672 50020 17696 50022
rect 17752 50020 17776 50022
rect 17832 50020 17856 50022
rect 17912 50020 17918 50022
rect 17610 50011 17918 50020
rect 17610 48988 17918 48997
rect 17610 48986 17616 48988
rect 17672 48986 17696 48988
rect 17752 48986 17776 48988
rect 17832 48986 17856 48988
rect 17912 48986 17918 48988
rect 17672 48934 17674 48986
rect 17854 48934 17856 48986
rect 17610 48932 17616 48934
rect 17672 48932 17696 48934
rect 17752 48932 17776 48934
rect 17832 48932 17856 48934
rect 17912 48932 17918 48934
rect 17610 48923 17918 48932
rect 17610 47900 17918 47909
rect 17610 47898 17616 47900
rect 17672 47898 17696 47900
rect 17752 47898 17776 47900
rect 17832 47898 17856 47900
rect 17912 47898 17918 47900
rect 17672 47846 17674 47898
rect 17854 47846 17856 47898
rect 17610 47844 17616 47846
rect 17672 47844 17696 47846
rect 17752 47844 17776 47846
rect 17832 47844 17856 47846
rect 17912 47844 17918 47846
rect 17610 47835 17918 47844
rect 17610 46812 17918 46821
rect 17610 46810 17616 46812
rect 17672 46810 17696 46812
rect 17752 46810 17776 46812
rect 17832 46810 17856 46812
rect 17912 46810 17918 46812
rect 17672 46758 17674 46810
rect 17854 46758 17856 46810
rect 17610 46756 17616 46758
rect 17672 46756 17696 46758
rect 17752 46756 17776 46758
rect 17832 46756 17856 46758
rect 17912 46756 17918 46758
rect 17610 46747 17918 46756
rect 18156 45898 18184 51886
rect 18144 45892 18196 45898
rect 18144 45834 18196 45840
rect 17610 45724 17918 45733
rect 17610 45722 17616 45724
rect 17672 45722 17696 45724
rect 17752 45722 17776 45724
rect 17832 45722 17856 45724
rect 17912 45722 17918 45724
rect 17672 45670 17674 45722
rect 17854 45670 17856 45722
rect 17610 45668 17616 45670
rect 17672 45668 17696 45670
rect 17752 45668 17776 45670
rect 17832 45668 17856 45670
rect 17912 45668 17918 45670
rect 17610 45659 17918 45668
rect 17610 44636 17918 44645
rect 17610 44634 17616 44636
rect 17672 44634 17696 44636
rect 17752 44634 17776 44636
rect 17832 44634 17856 44636
rect 17912 44634 17918 44636
rect 17672 44582 17674 44634
rect 17854 44582 17856 44634
rect 17610 44580 17616 44582
rect 17672 44580 17696 44582
rect 17752 44580 17776 44582
rect 17832 44580 17856 44582
rect 17912 44580 17918 44582
rect 17610 44571 17918 44580
rect 17610 43548 17918 43557
rect 17610 43546 17616 43548
rect 17672 43546 17696 43548
rect 17752 43546 17776 43548
rect 17832 43546 17856 43548
rect 17912 43546 17918 43548
rect 17672 43494 17674 43546
rect 17854 43494 17856 43546
rect 17610 43492 17616 43494
rect 17672 43492 17696 43494
rect 17752 43492 17776 43494
rect 17832 43492 17856 43494
rect 17912 43492 17918 43494
rect 17610 43483 17918 43492
rect 17610 42460 17918 42469
rect 17610 42458 17616 42460
rect 17672 42458 17696 42460
rect 17752 42458 17776 42460
rect 17832 42458 17856 42460
rect 17912 42458 17918 42460
rect 17672 42406 17674 42458
rect 17854 42406 17856 42458
rect 17610 42404 17616 42406
rect 17672 42404 17696 42406
rect 17752 42404 17776 42406
rect 17832 42404 17856 42406
rect 17912 42404 17918 42406
rect 17610 42395 17918 42404
rect 17610 41372 17918 41381
rect 17610 41370 17616 41372
rect 17672 41370 17696 41372
rect 17752 41370 17776 41372
rect 17832 41370 17856 41372
rect 17912 41370 17918 41372
rect 17672 41318 17674 41370
rect 17854 41318 17856 41370
rect 17610 41316 17616 41318
rect 17672 41316 17696 41318
rect 17752 41316 17776 41318
rect 17832 41316 17856 41318
rect 17912 41316 17918 41318
rect 17610 41307 17918 41316
rect 17610 40284 17918 40293
rect 17610 40282 17616 40284
rect 17672 40282 17696 40284
rect 17752 40282 17776 40284
rect 17832 40282 17856 40284
rect 17912 40282 17918 40284
rect 17672 40230 17674 40282
rect 17854 40230 17856 40282
rect 17610 40228 17616 40230
rect 17672 40228 17696 40230
rect 17752 40228 17776 40230
rect 17832 40228 17856 40230
rect 17912 40228 17918 40230
rect 17610 40219 17918 40228
rect 17610 39196 17918 39205
rect 17610 39194 17616 39196
rect 17672 39194 17696 39196
rect 17752 39194 17776 39196
rect 17832 39194 17856 39196
rect 17912 39194 17918 39196
rect 17672 39142 17674 39194
rect 17854 39142 17856 39194
rect 17610 39140 17616 39142
rect 17672 39140 17696 39142
rect 17752 39140 17776 39142
rect 17832 39140 17856 39142
rect 17912 39140 17918 39142
rect 17610 39131 17918 39140
rect 17610 38108 17918 38117
rect 17610 38106 17616 38108
rect 17672 38106 17696 38108
rect 17752 38106 17776 38108
rect 17832 38106 17856 38108
rect 17912 38106 17918 38108
rect 17672 38054 17674 38106
rect 17854 38054 17856 38106
rect 17610 38052 17616 38054
rect 17672 38052 17696 38054
rect 17752 38052 17776 38054
rect 17832 38052 17856 38054
rect 17912 38052 17918 38054
rect 17610 38043 17918 38052
rect 18052 37732 18104 37738
rect 18052 37674 18104 37680
rect 17960 37120 18012 37126
rect 17960 37062 18012 37068
rect 17610 37020 17918 37029
rect 17610 37018 17616 37020
rect 17672 37018 17696 37020
rect 17752 37018 17776 37020
rect 17832 37018 17856 37020
rect 17912 37018 17918 37020
rect 17672 36966 17674 37018
rect 17854 36966 17856 37018
rect 17610 36964 17616 36966
rect 17672 36964 17696 36966
rect 17752 36964 17776 36966
rect 17832 36964 17856 36966
rect 17912 36964 17918 36966
rect 17610 36955 17918 36964
rect 17610 35932 17918 35941
rect 17610 35930 17616 35932
rect 17672 35930 17696 35932
rect 17752 35930 17776 35932
rect 17832 35930 17856 35932
rect 17912 35930 17918 35932
rect 17672 35878 17674 35930
rect 17854 35878 17856 35930
rect 17610 35876 17616 35878
rect 17672 35876 17696 35878
rect 17752 35876 17776 35878
rect 17832 35876 17856 35878
rect 17912 35876 17918 35878
rect 17610 35867 17918 35876
rect 17592 35692 17644 35698
rect 17592 35634 17644 35640
rect 17604 35018 17632 35634
rect 17684 35624 17736 35630
rect 17684 35566 17736 35572
rect 17696 35086 17724 35566
rect 17684 35080 17736 35086
rect 17684 35022 17736 35028
rect 17592 35012 17644 35018
rect 17592 34954 17644 34960
rect 17610 34844 17918 34853
rect 17610 34842 17616 34844
rect 17672 34842 17696 34844
rect 17752 34842 17776 34844
rect 17832 34842 17856 34844
rect 17912 34842 17918 34844
rect 17672 34790 17674 34842
rect 17854 34790 17856 34842
rect 17610 34788 17616 34790
rect 17672 34788 17696 34790
rect 17752 34788 17776 34790
rect 17832 34788 17856 34790
rect 17912 34788 17918 34790
rect 17610 34779 17918 34788
rect 17610 33756 17918 33765
rect 17610 33754 17616 33756
rect 17672 33754 17696 33756
rect 17752 33754 17776 33756
rect 17832 33754 17856 33756
rect 17912 33754 17918 33756
rect 17672 33702 17674 33754
rect 17854 33702 17856 33754
rect 17610 33700 17616 33702
rect 17672 33700 17696 33702
rect 17752 33700 17776 33702
rect 17832 33700 17856 33702
rect 17912 33700 17918 33702
rect 17610 33691 17918 33700
rect 17500 33652 17552 33658
rect 17500 33594 17552 33600
rect 17420 33522 17908 33538
rect 17420 33516 17920 33522
rect 17420 33510 17868 33516
rect 16950 33212 17258 33221
rect 16950 33210 16956 33212
rect 17012 33210 17036 33212
rect 17092 33210 17116 33212
rect 17172 33210 17196 33212
rect 17252 33210 17258 33212
rect 17012 33158 17014 33210
rect 17194 33158 17196 33210
rect 16950 33156 16956 33158
rect 17012 33156 17036 33158
rect 17092 33156 17116 33158
rect 17172 33156 17196 33158
rect 17252 33156 17258 33158
rect 16950 33147 17258 33156
rect 17408 32904 17460 32910
rect 17408 32846 17460 32852
rect 16856 32836 16908 32842
rect 16856 32778 16908 32784
rect 16764 31952 16816 31958
rect 16764 31894 16816 31900
rect 16868 31754 16896 32778
rect 16948 32496 17000 32502
rect 17132 32496 17184 32502
rect 17000 32444 17132 32450
rect 16948 32438 17184 32444
rect 16960 32422 17172 32438
rect 16950 32124 17258 32133
rect 16950 32122 16956 32124
rect 17012 32122 17036 32124
rect 17092 32122 17116 32124
rect 17172 32122 17196 32124
rect 17252 32122 17258 32124
rect 17012 32070 17014 32122
rect 17194 32070 17196 32122
rect 16950 32068 16956 32070
rect 17012 32068 17036 32070
rect 17092 32068 17116 32070
rect 17172 32068 17196 32070
rect 17252 32068 17258 32070
rect 16950 32059 17258 32068
rect 17316 31952 17368 31958
rect 17316 31894 17368 31900
rect 16776 31726 16896 31754
rect 16672 31476 16724 31482
rect 16672 31418 16724 31424
rect 16500 31334 16712 31362
rect 16408 31198 16620 31226
rect 16488 30932 16540 30938
rect 16488 30874 16540 30880
rect 16132 30790 16252 30818
rect 16132 22094 16160 30790
rect 16304 29096 16356 29102
rect 16304 29038 16356 29044
rect 16316 25498 16344 29038
rect 16396 26444 16448 26450
rect 16396 26386 16448 26392
rect 16304 25492 16356 25498
rect 16304 25434 16356 25440
rect 16132 22066 16252 22094
rect 16028 9512 16080 9518
rect 16028 9454 16080 9460
rect 16224 8362 16252 22066
rect 16212 8356 16264 8362
rect 16212 8298 16264 8304
rect 16408 7954 16436 26386
rect 16500 12238 16528 30874
rect 16592 27062 16620 31198
rect 16684 30258 16712 31334
rect 16672 30252 16724 30258
rect 16672 30194 16724 30200
rect 16684 29034 16712 30194
rect 16672 29028 16724 29034
rect 16672 28970 16724 28976
rect 16672 28484 16724 28490
rect 16672 28426 16724 28432
rect 16580 27056 16632 27062
rect 16580 26998 16632 27004
rect 16578 26888 16634 26897
rect 16578 26823 16634 26832
rect 16592 15094 16620 26823
rect 16580 15088 16632 15094
rect 16580 15030 16632 15036
rect 16578 13424 16634 13433
rect 16578 13359 16634 13368
rect 16488 12232 16540 12238
rect 16488 12174 16540 12180
rect 16592 11150 16620 13359
rect 16580 11144 16632 11150
rect 16580 11086 16632 11092
rect 16580 9580 16632 9586
rect 16580 9522 16632 9528
rect 16592 8906 16620 9522
rect 16684 9382 16712 28426
rect 16672 9376 16724 9382
rect 16672 9318 16724 9324
rect 16580 8900 16632 8906
rect 16580 8842 16632 8848
rect 16672 8356 16724 8362
rect 16672 8298 16724 8304
rect 16396 7948 16448 7954
rect 16396 7890 16448 7896
rect 15752 7404 15804 7410
rect 15752 7346 15804 7352
rect 16684 6322 16712 8298
rect 16776 6322 16804 31726
rect 16856 31680 16908 31686
rect 16856 31622 16908 31628
rect 16868 28762 16896 31622
rect 16950 31036 17258 31045
rect 16950 31034 16956 31036
rect 17012 31034 17036 31036
rect 17092 31034 17116 31036
rect 17172 31034 17196 31036
rect 17252 31034 17258 31036
rect 17012 30982 17014 31034
rect 17194 30982 17196 31034
rect 16950 30980 16956 30982
rect 17012 30980 17036 30982
rect 17092 30980 17116 30982
rect 17172 30980 17196 30982
rect 17252 30980 17258 30982
rect 16950 30971 17258 30980
rect 16950 29948 17258 29957
rect 16950 29946 16956 29948
rect 17012 29946 17036 29948
rect 17092 29946 17116 29948
rect 17172 29946 17196 29948
rect 17252 29946 17258 29948
rect 17012 29894 17014 29946
rect 17194 29894 17196 29946
rect 16950 29892 16956 29894
rect 17012 29892 17036 29894
rect 17092 29892 17116 29894
rect 17172 29892 17196 29894
rect 17252 29892 17258 29894
rect 16950 29883 17258 29892
rect 16948 29572 17000 29578
rect 16948 29514 17000 29520
rect 16960 29102 16988 29514
rect 16948 29096 17000 29102
rect 16948 29038 17000 29044
rect 16950 28860 17258 28869
rect 16950 28858 16956 28860
rect 17012 28858 17036 28860
rect 17092 28858 17116 28860
rect 17172 28858 17196 28860
rect 17252 28858 17258 28860
rect 17012 28806 17014 28858
rect 17194 28806 17196 28858
rect 16950 28804 16956 28806
rect 17012 28804 17036 28806
rect 17092 28804 17116 28806
rect 17172 28804 17196 28806
rect 17252 28804 17258 28806
rect 16950 28795 17258 28804
rect 16856 28756 16908 28762
rect 16856 28698 16908 28704
rect 16948 28756 17000 28762
rect 16948 28698 17000 28704
rect 16868 25770 16896 28698
rect 16960 28558 16988 28698
rect 16948 28552 17000 28558
rect 16948 28494 17000 28500
rect 16960 28218 16988 28494
rect 16948 28212 17000 28218
rect 16948 28154 17000 28160
rect 16950 27772 17258 27781
rect 16950 27770 16956 27772
rect 17012 27770 17036 27772
rect 17092 27770 17116 27772
rect 17172 27770 17196 27772
rect 17252 27770 17258 27772
rect 17012 27718 17014 27770
rect 17194 27718 17196 27770
rect 16950 27716 16956 27718
rect 17012 27716 17036 27718
rect 17092 27716 17116 27718
rect 17172 27716 17196 27718
rect 17252 27716 17258 27718
rect 16950 27707 17258 27716
rect 17224 27668 17276 27674
rect 17224 27610 17276 27616
rect 17236 26874 17264 27610
rect 17328 27033 17356 31894
rect 17420 31822 17448 32846
rect 17408 31816 17460 31822
rect 17408 31758 17460 31764
rect 17420 31346 17448 31758
rect 17408 31340 17460 31346
rect 17408 31282 17460 31288
rect 17408 29708 17460 29714
rect 17408 29650 17460 29656
rect 17420 29170 17448 29650
rect 17408 29164 17460 29170
rect 17408 29106 17460 29112
rect 17420 28626 17448 29106
rect 17408 28620 17460 28626
rect 17408 28562 17460 28568
rect 17408 28212 17460 28218
rect 17408 28154 17460 28160
rect 17420 27674 17448 28154
rect 17408 27668 17460 27674
rect 17408 27610 17460 27616
rect 17408 27056 17460 27062
rect 17314 27024 17370 27033
rect 17408 26998 17460 27004
rect 17314 26959 17370 26968
rect 17236 26846 17356 26874
rect 16950 26684 17258 26693
rect 16950 26682 16956 26684
rect 17012 26682 17036 26684
rect 17092 26682 17116 26684
rect 17172 26682 17196 26684
rect 17252 26682 17258 26684
rect 17012 26630 17014 26682
rect 17194 26630 17196 26682
rect 16950 26628 16956 26630
rect 17012 26628 17036 26630
rect 17092 26628 17116 26630
rect 17172 26628 17196 26630
rect 17252 26628 17258 26630
rect 16950 26619 17258 26628
rect 17224 26376 17276 26382
rect 17224 26318 17276 26324
rect 17236 25838 17264 26318
rect 17224 25832 17276 25838
rect 17224 25774 17276 25780
rect 16856 25764 16908 25770
rect 16856 25706 16908 25712
rect 16950 25596 17258 25605
rect 16950 25594 16956 25596
rect 17012 25594 17036 25596
rect 17092 25594 17116 25596
rect 17172 25594 17196 25596
rect 17252 25594 17258 25596
rect 17012 25542 17014 25594
rect 17194 25542 17196 25594
rect 16950 25540 16956 25542
rect 17012 25540 17036 25542
rect 17092 25540 17116 25542
rect 17172 25540 17196 25542
rect 17252 25540 17258 25542
rect 16950 25531 17258 25540
rect 16856 25492 16908 25498
rect 16856 25434 16908 25440
rect 16868 9654 16896 25434
rect 17328 25362 17356 26846
rect 17420 25922 17448 26998
rect 17512 26042 17540 33510
rect 17868 33458 17920 33464
rect 17610 32668 17918 32677
rect 17610 32666 17616 32668
rect 17672 32666 17696 32668
rect 17752 32666 17776 32668
rect 17832 32666 17856 32668
rect 17912 32666 17918 32668
rect 17672 32614 17674 32666
rect 17854 32614 17856 32666
rect 17610 32612 17616 32614
rect 17672 32612 17696 32614
rect 17752 32612 17776 32614
rect 17832 32612 17856 32614
rect 17912 32612 17918 32614
rect 17610 32603 17918 32612
rect 17610 31580 17918 31589
rect 17610 31578 17616 31580
rect 17672 31578 17696 31580
rect 17752 31578 17776 31580
rect 17832 31578 17856 31580
rect 17912 31578 17918 31580
rect 17672 31526 17674 31578
rect 17854 31526 17856 31578
rect 17610 31524 17616 31526
rect 17672 31524 17696 31526
rect 17752 31524 17776 31526
rect 17832 31524 17856 31526
rect 17912 31524 17918 31526
rect 17610 31515 17918 31524
rect 17868 30932 17920 30938
rect 17868 30874 17920 30880
rect 17880 30682 17908 30874
rect 17972 30802 18000 37062
rect 18064 32978 18092 37674
rect 18052 32972 18104 32978
rect 18052 32914 18104 32920
rect 18052 32224 18104 32230
rect 18052 32166 18104 32172
rect 17960 30796 18012 30802
rect 17960 30738 18012 30744
rect 17880 30654 18000 30682
rect 17610 30492 17918 30501
rect 17610 30490 17616 30492
rect 17672 30490 17696 30492
rect 17752 30490 17776 30492
rect 17832 30490 17856 30492
rect 17912 30490 17918 30492
rect 17672 30438 17674 30490
rect 17854 30438 17856 30490
rect 17610 30436 17616 30438
rect 17672 30436 17696 30438
rect 17752 30436 17776 30438
rect 17832 30436 17856 30438
rect 17912 30436 17918 30438
rect 17610 30427 17918 30436
rect 17972 30274 18000 30654
rect 17880 30246 18000 30274
rect 17880 29578 17908 30246
rect 17868 29572 17920 29578
rect 17868 29514 17920 29520
rect 17610 29404 17918 29413
rect 17610 29402 17616 29404
rect 17672 29402 17696 29404
rect 17752 29402 17776 29404
rect 17832 29402 17856 29404
rect 17912 29402 17918 29404
rect 17672 29350 17674 29402
rect 17854 29350 17856 29402
rect 17610 29348 17616 29350
rect 17672 29348 17696 29350
rect 17752 29348 17776 29350
rect 17832 29348 17856 29350
rect 17912 29348 17918 29350
rect 17610 29339 17918 29348
rect 17868 29028 17920 29034
rect 17868 28970 17920 28976
rect 17776 28960 17828 28966
rect 17776 28902 17828 28908
rect 17788 28626 17816 28902
rect 17776 28620 17828 28626
rect 17776 28562 17828 28568
rect 17880 28506 17908 28970
rect 17880 28478 18000 28506
rect 17610 28316 17918 28325
rect 17610 28314 17616 28316
rect 17672 28314 17696 28316
rect 17752 28314 17776 28316
rect 17832 28314 17856 28316
rect 17912 28314 17918 28316
rect 17672 28262 17674 28314
rect 17854 28262 17856 28314
rect 17610 28260 17616 28262
rect 17672 28260 17696 28262
rect 17752 28260 17776 28262
rect 17832 28260 17856 28262
rect 17912 28260 17918 28262
rect 17610 28251 17918 28260
rect 17972 28098 18000 28478
rect 17880 28070 18000 28098
rect 17880 27418 17908 28070
rect 17880 27390 18000 27418
rect 17610 27228 17918 27237
rect 17610 27226 17616 27228
rect 17672 27226 17696 27228
rect 17752 27226 17776 27228
rect 17832 27226 17856 27228
rect 17912 27226 17918 27228
rect 17672 27174 17674 27226
rect 17854 27174 17856 27226
rect 17610 27172 17616 27174
rect 17672 27172 17696 27174
rect 17752 27172 17776 27174
rect 17832 27172 17856 27174
rect 17912 27172 17918 27174
rect 17610 27163 17918 27172
rect 17972 27010 18000 27390
rect 17880 26982 18000 27010
rect 17592 26852 17644 26858
rect 17592 26794 17644 26800
rect 17604 26382 17632 26794
rect 17592 26376 17644 26382
rect 17592 26318 17644 26324
rect 17880 26330 17908 26982
rect 17880 26302 18000 26330
rect 17610 26140 17918 26149
rect 17610 26138 17616 26140
rect 17672 26138 17696 26140
rect 17752 26138 17776 26140
rect 17832 26138 17856 26140
rect 17912 26138 17918 26140
rect 17672 26086 17674 26138
rect 17854 26086 17856 26138
rect 17610 26084 17616 26086
rect 17672 26084 17696 26086
rect 17752 26084 17776 26086
rect 17832 26084 17856 26086
rect 17912 26084 17918 26086
rect 17610 26075 17918 26084
rect 17500 26036 17552 26042
rect 17500 25978 17552 25984
rect 17972 25922 18000 26302
rect 18064 25974 18092 32166
rect 17420 25894 17540 25922
rect 17408 25832 17460 25838
rect 17408 25774 17460 25780
rect 17316 25356 17368 25362
rect 17316 25298 17368 25304
rect 17316 25220 17368 25226
rect 17316 25162 17368 25168
rect 16950 24508 17258 24517
rect 16950 24506 16956 24508
rect 17012 24506 17036 24508
rect 17092 24506 17116 24508
rect 17172 24506 17196 24508
rect 17252 24506 17258 24508
rect 17012 24454 17014 24506
rect 17194 24454 17196 24506
rect 16950 24452 16956 24454
rect 17012 24452 17036 24454
rect 17092 24452 17116 24454
rect 17172 24452 17196 24454
rect 17252 24452 17258 24454
rect 16950 24443 17258 24452
rect 16950 23420 17258 23429
rect 16950 23418 16956 23420
rect 17012 23418 17036 23420
rect 17092 23418 17116 23420
rect 17172 23418 17196 23420
rect 17252 23418 17258 23420
rect 17012 23366 17014 23418
rect 17194 23366 17196 23418
rect 16950 23364 16956 23366
rect 17012 23364 17036 23366
rect 17092 23364 17116 23366
rect 17172 23364 17196 23366
rect 17252 23364 17258 23366
rect 16950 23355 17258 23364
rect 17328 23322 17356 25162
rect 17316 23316 17368 23322
rect 17316 23258 17368 23264
rect 17420 22778 17448 25774
rect 17408 22772 17460 22778
rect 17408 22714 17460 22720
rect 17316 22636 17368 22642
rect 17316 22578 17368 22584
rect 17328 22386 17356 22578
rect 17328 22358 17448 22386
rect 16950 22332 17258 22341
rect 16950 22330 16956 22332
rect 17012 22330 17036 22332
rect 17092 22330 17116 22332
rect 17172 22330 17196 22332
rect 17252 22330 17258 22332
rect 17012 22278 17014 22330
rect 17194 22278 17196 22330
rect 16950 22276 16956 22278
rect 17012 22276 17036 22278
rect 17092 22276 17116 22278
rect 17172 22276 17196 22278
rect 17252 22276 17258 22278
rect 16950 22267 17258 22276
rect 17316 22228 17368 22234
rect 17316 22170 17368 22176
rect 17224 22092 17276 22098
rect 17224 22034 17276 22040
rect 17236 21418 17264 22034
rect 17224 21412 17276 21418
rect 17224 21354 17276 21360
rect 16950 21244 17258 21253
rect 16950 21242 16956 21244
rect 17012 21242 17036 21244
rect 17092 21242 17116 21244
rect 17172 21242 17196 21244
rect 17252 21242 17258 21244
rect 17012 21190 17014 21242
rect 17194 21190 17196 21242
rect 16950 21188 16956 21190
rect 17012 21188 17036 21190
rect 17092 21188 17116 21190
rect 17172 21188 17196 21190
rect 17252 21188 17258 21190
rect 16950 21179 17258 21188
rect 16950 20156 17258 20165
rect 16950 20154 16956 20156
rect 17012 20154 17036 20156
rect 17092 20154 17116 20156
rect 17172 20154 17196 20156
rect 17252 20154 17258 20156
rect 17012 20102 17014 20154
rect 17194 20102 17196 20154
rect 16950 20100 16956 20102
rect 17012 20100 17036 20102
rect 17092 20100 17116 20102
rect 17172 20100 17196 20102
rect 17252 20100 17258 20102
rect 16950 20091 17258 20100
rect 16950 19068 17258 19077
rect 16950 19066 16956 19068
rect 17012 19066 17036 19068
rect 17092 19066 17116 19068
rect 17172 19066 17196 19068
rect 17252 19066 17258 19068
rect 17012 19014 17014 19066
rect 17194 19014 17196 19066
rect 16950 19012 16956 19014
rect 17012 19012 17036 19014
rect 17092 19012 17116 19014
rect 17172 19012 17196 19014
rect 17252 19012 17258 19014
rect 16950 19003 17258 19012
rect 16950 17980 17258 17989
rect 16950 17978 16956 17980
rect 17012 17978 17036 17980
rect 17092 17978 17116 17980
rect 17172 17978 17196 17980
rect 17252 17978 17258 17980
rect 17012 17926 17014 17978
rect 17194 17926 17196 17978
rect 16950 17924 16956 17926
rect 17012 17924 17036 17926
rect 17092 17924 17116 17926
rect 17172 17924 17196 17926
rect 17252 17924 17258 17926
rect 16950 17915 17258 17924
rect 16950 16892 17258 16901
rect 16950 16890 16956 16892
rect 17012 16890 17036 16892
rect 17092 16890 17116 16892
rect 17172 16890 17196 16892
rect 17252 16890 17258 16892
rect 17012 16838 17014 16890
rect 17194 16838 17196 16890
rect 16950 16836 16956 16838
rect 17012 16836 17036 16838
rect 17092 16836 17116 16838
rect 17172 16836 17196 16838
rect 17252 16836 17258 16838
rect 16950 16827 17258 16836
rect 16950 15804 17258 15813
rect 16950 15802 16956 15804
rect 17012 15802 17036 15804
rect 17092 15802 17116 15804
rect 17172 15802 17196 15804
rect 17252 15802 17258 15804
rect 17012 15750 17014 15802
rect 17194 15750 17196 15802
rect 16950 15748 16956 15750
rect 17012 15748 17036 15750
rect 17092 15748 17116 15750
rect 17172 15748 17196 15750
rect 17252 15748 17258 15750
rect 16950 15739 17258 15748
rect 17224 15156 17276 15162
rect 17224 15098 17276 15104
rect 17236 14958 17264 15098
rect 17224 14952 17276 14958
rect 17224 14894 17276 14900
rect 16950 14716 17258 14725
rect 16950 14714 16956 14716
rect 17012 14714 17036 14716
rect 17092 14714 17116 14716
rect 17172 14714 17196 14716
rect 17252 14714 17258 14716
rect 17012 14662 17014 14714
rect 17194 14662 17196 14714
rect 16950 14660 16956 14662
rect 17012 14660 17036 14662
rect 17092 14660 17116 14662
rect 17172 14660 17196 14662
rect 17252 14660 17258 14662
rect 16950 14651 17258 14660
rect 16950 13628 17258 13637
rect 16950 13626 16956 13628
rect 17012 13626 17036 13628
rect 17092 13626 17116 13628
rect 17172 13626 17196 13628
rect 17252 13626 17258 13628
rect 17012 13574 17014 13626
rect 17194 13574 17196 13626
rect 16950 13572 16956 13574
rect 17012 13572 17036 13574
rect 17092 13572 17116 13574
rect 17172 13572 17196 13574
rect 17252 13572 17258 13574
rect 16950 13563 17258 13572
rect 16950 12540 17258 12549
rect 16950 12538 16956 12540
rect 17012 12538 17036 12540
rect 17092 12538 17116 12540
rect 17172 12538 17196 12540
rect 17252 12538 17258 12540
rect 17012 12486 17014 12538
rect 17194 12486 17196 12538
rect 16950 12484 16956 12486
rect 17012 12484 17036 12486
rect 17092 12484 17116 12486
rect 17172 12484 17196 12486
rect 17252 12484 17258 12486
rect 16950 12475 17258 12484
rect 16950 11452 17258 11461
rect 16950 11450 16956 11452
rect 17012 11450 17036 11452
rect 17092 11450 17116 11452
rect 17172 11450 17196 11452
rect 17252 11450 17258 11452
rect 17012 11398 17014 11450
rect 17194 11398 17196 11450
rect 16950 11396 16956 11398
rect 17012 11396 17036 11398
rect 17092 11396 17116 11398
rect 17172 11396 17196 11398
rect 17252 11396 17258 11398
rect 16950 11387 17258 11396
rect 16950 10364 17258 10373
rect 16950 10362 16956 10364
rect 17012 10362 17036 10364
rect 17092 10362 17116 10364
rect 17172 10362 17196 10364
rect 17252 10362 17258 10364
rect 17012 10310 17014 10362
rect 17194 10310 17196 10362
rect 16950 10308 16956 10310
rect 17012 10308 17036 10310
rect 17092 10308 17116 10310
rect 17172 10308 17196 10310
rect 17252 10308 17258 10310
rect 16950 10299 17258 10308
rect 16856 9648 16908 9654
rect 16856 9590 16908 9596
rect 16950 9276 17258 9285
rect 16950 9274 16956 9276
rect 17012 9274 17036 9276
rect 17092 9274 17116 9276
rect 17172 9274 17196 9276
rect 17252 9274 17258 9276
rect 17012 9222 17014 9274
rect 17194 9222 17196 9274
rect 16950 9220 16956 9222
rect 17012 9220 17036 9222
rect 17092 9220 17116 9222
rect 17172 9220 17196 9222
rect 17252 9220 17258 9222
rect 16950 9211 17258 9220
rect 16950 8188 17258 8197
rect 16950 8186 16956 8188
rect 17012 8186 17036 8188
rect 17092 8186 17116 8188
rect 17172 8186 17196 8188
rect 17252 8186 17258 8188
rect 17012 8134 17014 8186
rect 17194 8134 17196 8186
rect 16950 8132 16956 8134
rect 17012 8132 17036 8134
rect 17092 8132 17116 8134
rect 17172 8132 17196 8134
rect 17252 8132 17258 8134
rect 16950 8123 17258 8132
rect 16950 7100 17258 7109
rect 16950 7098 16956 7100
rect 17012 7098 17036 7100
rect 17092 7098 17116 7100
rect 17172 7098 17196 7100
rect 17252 7098 17258 7100
rect 17012 7046 17014 7098
rect 17194 7046 17196 7098
rect 16950 7044 16956 7046
rect 17012 7044 17036 7046
rect 17092 7044 17116 7046
rect 17172 7044 17196 7046
rect 17252 7044 17258 7046
rect 16950 7035 17258 7044
rect 16948 6724 17000 6730
rect 16948 6666 17000 6672
rect 16960 6322 16988 6666
rect 16672 6316 16724 6322
rect 16672 6258 16724 6264
rect 16764 6316 16816 6322
rect 16764 6258 16816 6264
rect 16948 6316 17000 6322
rect 16948 6258 17000 6264
rect 16950 6012 17258 6021
rect 16950 6010 16956 6012
rect 17012 6010 17036 6012
rect 17092 6010 17116 6012
rect 17172 6010 17196 6012
rect 17252 6010 17258 6012
rect 17012 5958 17014 6010
rect 17194 5958 17196 6010
rect 16950 5956 16956 5958
rect 17012 5956 17036 5958
rect 17092 5956 17116 5958
rect 17172 5956 17196 5958
rect 17252 5956 17258 5958
rect 16950 5947 17258 5956
rect 16950 4924 17258 4933
rect 16950 4922 16956 4924
rect 17012 4922 17036 4924
rect 17092 4922 17116 4924
rect 17172 4922 17196 4924
rect 17252 4922 17258 4924
rect 17012 4870 17014 4922
rect 17194 4870 17196 4922
rect 16950 4868 16956 4870
rect 17012 4868 17036 4870
rect 17092 4868 17116 4870
rect 17172 4868 17196 4870
rect 17252 4868 17258 4870
rect 16950 4859 17258 4868
rect 16950 3836 17258 3845
rect 16950 3834 16956 3836
rect 17012 3834 17036 3836
rect 17092 3834 17116 3836
rect 17172 3834 17196 3836
rect 17252 3834 17258 3836
rect 17012 3782 17014 3834
rect 17194 3782 17196 3834
rect 16950 3780 16956 3782
rect 17012 3780 17036 3782
rect 17092 3780 17116 3782
rect 17172 3780 17196 3782
rect 17252 3780 17258 3782
rect 16950 3771 17258 3780
rect 14464 3528 14516 3534
rect 14464 3470 14516 3476
rect 17328 2854 17356 22170
rect 17420 22098 17448 22358
rect 17408 22092 17460 22098
rect 17408 22034 17460 22040
rect 17512 21978 17540 25894
rect 17880 25894 18000 25922
rect 18052 25968 18104 25974
rect 18052 25910 18104 25916
rect 17880 25226 17908 25894
rect 17868 25220 17920 25226
rect 17868 25162 17920 25168
rect 17610 25052 17918 25061
rect 17610 25050 17616 25052
rect 17672 25050 17696 25052
rect 17752 25050 17776 25052
rect 17832 25050 17856 25052
rect 17912 25050 17918 25052
rect 17672 24998 17674 25050
rect 17854 24998 17856 25050
rect 17610 24996 17616 24998
rect 17672 24996 17696 24998
rect 17752 24996 17776 24998
rect 17832 24996 17856 24998
rect 17912 24996 17918 24998
rect 17610 24987 17918 24996
rect 18156 24206 18184 45834
rect 18236 33584 18288 33590
rect 18236 33526 18288 33532
rect 18248 31754 18276 33526
rect 18340 32230 18368 67050
rect 18616 60722 18644 67186
rect 18972 66564 19024 66570
rect 18972 66506 19024 66512
rect 18880 66020 18932 66026
rect 18880 65962 18932 65968
rect 18788 61600 18840 61606
rect 18788 61542 18840 61548
rect 18604 60716 18656 60722
rect 18604 60658 18656 60664
rect 18512 59492 18564 59498
rect 18512 59434 18564 59440
rect 18524 42294 18552 59434
rect 18616 59430 18644 60658
rect 18604 59424 18656 59430
rect 18604 59366 18656 59372
rect 18696 44532 18748 44538
rect 18696 44474 18748 44480
rect 18604 42628 18656 42634
rect 18604 42570 18656 42576
rect 18512 42288 18564 42294
rect 18512 42230 18564 42236
rect 18616 42090 18644 42570
rect 18604 42084 18656 42090
rect 18604 42026 18656 42032
rect 18616 37466 18644 42026
rect 18604 37460 18656 37466
rect 18604 37402 18656 37408
rect 18420 33312 18472 33318
rect 18420 33254 18472 33260
rect 18328 32224 18380 32230
rect 18328 32166 18380 32172
rect 18340 32026 18368 32166
rect 18328 32020 18380 32026
rect 18328 31962 18380 31968
rect 18432 31906 18460 33254
rect 18432 31878 18552 31906
rect 18248 31726 18460 31754
rect 18328 31340 18380 31346
rect 18328 31282 18380 31288
rect 18236 30796 18288 30802
rect 18236 30738 18288 30744
rect 18144 24200 18196 24206
rect 18144 24142 18196 24148
rect 17610 23964 17918 23973
rect 17610 23962 17616 23964
rect 17672 23962 17696 23964
rect 17752 23962 17776 23964
rect 17832 23962 17856 23964
rect 17912 23962 17918 23964
rect 17672 23910 17674 23962
rect 17854 23910 17856 23962
rect 17610 23908 17616 23910
rect 17672 23908 17696 23910
rect 17752 23908 17776 23910
rect 17832 23908 17856 23910
rect 17912 23908 17918 23910
rect 17610 23899 17918 23908
rect 17960 23112 18012 23118
rect 17960 23054 18012 23060
rect 17610 22876 17918 22885
rect 17610 22874 17616 22876
rect 17672 22874 17696 22876
rect 17752 22874 17776 22876
rect 17832 22874 17856 22876
rect 17912 22874 17918 22876
rect 17672 22822 17674 22874
rect 17854 22822 17856 22874
rect 17610 22820 17616 22822
rect 17672 22820 17696 22822
rect 17752 22820 17776 22822
rect 17832 22820 17856 22822
rect 17912 22820 17918 22822
rect 17610 22811 17918 22820
rect 17972 22778 18000 23054
rect 17868 22772 17920 22778
rect 17868 22714 17920 22720
rect 17960 22772 18012 22778
rect 17960 22714 18012 22720
rect 17592 22636 17644 22642
rect 17592 22578 17644 22584
rect 17604 22234 17632 22578
rect 17592 22228 17644 22234
rect 17592 22170 17644 22176
rect 17420 21950 17540 21978
rect 17420 19786 17448 21950
rect 17880 21894 17908 22714
rect 17500 21888 17552 21894
rect 17500 21830 17552 21836
rect 17868 21888 17920 21894
rect 17868 21830 17920 21836
rect 17408 19780 17460 19786
rect 17408 19722 17460 19728
rect 17420 9450 17448 19722
rect 17408 9444 17460 9450
rect 17408 9386 17460 9392
rect 17512 6390 17540 21830
rect 17610 21788 17918 21797
rect 17610 21786 17616 21788
rect 17672 21786 17696 21788
rect 17752 21786 17776 21788
rect 17832 21786 17856 21788
rect 17912 21786 17918 21788
rect 17672 21734 17674 21786
rect 17854 21734 17856 21786
rect 17610 21732 17616 21734
rect 17672 21732 17696 21734
rect 17752 21732 17776 21734
rect 17832 21732 17856 21734
rect 17912 21732 17918 21734
rect 17610 21723 17918 21732
rect 17610 20700 17918 20709
rect 17610 20698 17616 20700
rect 17672 20698 17696 20700
rect 17752 20698 17776 20700
rect 17832 20698 17856 20700
rect 17912 20698 17918 20700
rect 17672 20646 17674 20698
rect 17854 20646 17856 20698
rect 17610 20644 17616 20646
rect 17672 20644 17696 20646
rect 17752 20644 17776 20646
rect 17832 20644 17856 20646
rect 17912 20644 17918 20646
rect 17610 20635 17918 20644
rect 17610 19612 17918 19621
rect 17610 19610 17616 19612
rect 17672 19610 17696 19612
rect 17752 19610 17776 19612
rect 17832 19610 17856 19612
rect 17912 19610 17918 19612
rect 17672 19558 17674 19610
rect 17854 19558 17856 19610
rect 17610 19556 17616 19558
rect 17672 19556 17696 19558
rect 17752 19556 17776 19558
rect 17832 19556 17856 19558
rect 17912 19556 17918 19558
rect 17610 19547 17918 19556
rect 17868 19168 17920 19174
rect 17868 19110 17920 19116
rect 17880 18766 17908 19110
rect 17868 18760 17920 18766
rect 17868 18702 17920 18708
rect 17610 18524 17918 18533
rect 17610 18522 17616 18524
rect 17672 18522 17696 18524
rect 17752 18522 17776 18524
rect 17832 18522 17856 18524
rect 17912 18522 17918 18524
rect 17672 18470 17674 18522
rect 17854 18470 17856 18522
rect 17610 18468 17616 18470
rect 17672 18468 17696 18470
rect 17752 18468 17776 18470
rect 17832 18468 17856 18470
rect 17912 18468 17918 18470
rect 17610 18459 17918 18468
rect 17610 17436 17918 17445
rect 17610 17434 17616 17436
rect 17672 17434 17696 17436
rect 17752 17434 17776 17436
rect 17832 17434 17856 17436
rect 17912 17434 17918 17436
rect 17672 17382 17674 17434
rect 17854 17382 17856 17434
rect 17610 17380 17616 17382
rect 17672 17380 17696 17382
rect 17752 17380 17776 17382
rect 17832 17380 17856 17382
rect 17912 17380 17918 17382
rect 17610 17371 17918 17380
rect 18156 17338 18184 24142
rect 18248 23118 18276 30738
rect 18340 29714 18368 31282
rect 18328 29708 18380 29714
rect 18328 29650 18380 29656
rect 18328 23316 18380 23322
rect 18328 23258 18380 23264
rect 18236 23112 18288 23118
rect 18236 23054 18288 23060
rect 18236 22976 18288 22982
rect 18236 22918 18288 22924
rect 18248 19922 18276 22918
rect 18340 22710 18368 23258
rect 18328 22704 18380 22710
rect 18328 22646 18380 22652
rect 18236 19916 18288 19922
rect 18236 19858 18288 19864
rect 18144 17332 18196 17338
rect 18144 17274 18196 17280
rect 17610 16348 17918 16357
rect 17610 16346 17616 16348
rect 17672 16346 17696 16348
rect 17752 16346 17776 16348
rect 17832 16346 17856 16348
rect 17912 16346 17918 16348
rect 17672 16294 17674 16346
rect 17854 16294 17856 16346
rect 17610 16292 17616 16294
rect 17672 16292 17696 16294
rect 17752 16292 17776 16294
rect 17832 16292 17856 16294
rect 17912 16292 17918 16294
rect 17610 16283 17918 16292
rect 17610 15260 17918 15269
rect 17610 15258 17616 15260
rect 17672 15258 17696 15260
rect 17752 15258 17776 15260
rect 17832 15258 17856 15260
rect 17912 15258 17918 15260
rect 17672 15206 17674 15258
rect 17854 15206 17856 15258
rect 17610 15204 17616 15206
rect 17672 15204 17696 15206
rect 17752 15204 17776 15206
rect 17832 15204 17856 15206
rect 17912 15204 17918 15206
rect 17610 15195 17918 15204
rect 17610 14172 17918 14181
rect 17610 14170 17616 14172
rect 17672 14170 17696 14172
rect 17752 14170 17776 14172
rect 17832 14170 17856 14172
rect 17912 14170 17918 14172
rect 17672 14118 17674 14170
rect 17854 14118 17856 14170
rect 17610 14116 17616 14118
rect 17672 14116 17696 14118
rect 17752 14116 17776 14118
rect 17832 14116 17856 14118
rect 17912 14116 17918 14118
rect 17610 14107 17918 14116
rect 17610 13084 17918 13093
rect 17610 13082 17616 13084
rect 17672 13082 17696 13084
rect 17752 13082 17776 13084
rect 17832 13082 17856 13084
rect 17912 13082 17918 13084
rect 17672 13030 17674 13082
rect 17854 13030 17856 13082
rect 17610 13028 17616 13030
rect 17672 13028 17696 13030
rect 17752 13028 17776 13030
rect 17832 13028 17856 13030
rect 17912 13028 17918 13030
rect 17610 13019 17918 13028
rect 17610 11996 17918 12005
rect 17610 11994 17616 11996
rect 17672 11994 17696 11996
rect 17752 11994 17776 11996
rect 17832 11994 17856 11996
rect 17912 11994 17918 11996
rect 17672 11942 17674 11994
rect 17854 11942 17856 11994
rect 17610 11940 17616 11942
rect 17672 11940 17696 11942
rect 17752 11940 17776 11942
rect 17832 11940 17856 11942
rect 17912 11940 17918 11942
rect 17610 11931 17918 11940
rect 17610 10908 17918 10917
rect 17610 10906 17616 10908
rect 17672 10906 17696 10908
rect 17752 10906 17776 10908
rect 17832 10906 17856 10908
rect 17912 10906 17918 10908
rect 17672 10854 17674 10906
rect 17854 10854 17856 10906
rect 17610 10852 17616 10854
rect 17672 10852 17696 10854
rect 17752 10852 17776 10854
rect 17832 10852 17856 10854
rect 17912 10852 17918 10854
rect 17610 10843 17918 10852
rect 17960 10532 18012 10538
rect 17960 10474 18012 10480
rect 17610 9820 17918 9829
rect 17610 9818 17616 9820
rect 17672 9818 17696 9820
rect 17752 9818 17776 9820
rect 17832 9818 17856 9820
rect 17912 9818 17918 9820
rect 17672 9766 17674 9818
rect 17854 9766 17856 9818
rect 17610 9764 17616 9766
rect 17672 9764 17696 9766
rect 17752 9764 17776 9766
rect 17832 9764 17856 9766
rect 17912 9764 17918 9766
rect 17610 9755 17918 9764
rect 17972 9586 18000 10474
rect 17960 9580 18012 9586
rect 17960 9522 18012 9528
rect 17610 8732 17918 8741
rect 17610 8730 17616 8732
rect 17672 8730 17696 8732
rect 17752 8730 17776 8732
rect 17832 8730 17856 8732
rect 17912 8730 17918 8732
rect 17672 8678 17674 8730
rect 17854 8678 17856 8730
rect 17610 8676 17616 8678
rect 17672 8676 17696 8678
rect 17752 8676 17776 8678
rect 17832 8676 17856 8678
rect 17912 8676 17918 8678
rect 17610 8667 17918 8676
rect 17610 7644 17918 7653
rect 17610 7642 17616 7644
rect 17672 7642 17696 7644
rect 17752 7642 17776 7644
rect 17832 7642 17856 7644
rect 17912 7642 17918 7644
rect 17672 7590 17674 7642
rect 17854 7590 17856 7642
rect 17610 7588 17616 7590
rect 17672 7588 17696 7590
rect 17752 7588 17776 7590
rect 17832 7588 17856 7590
rect 17912 7588 17918 7590
rect 17610 7579 17918 7588
rect 18340 6914 18368 22646
rect 18432 20058 18460 31726
rect 18524 31142 18552 31878
rect 18512 31136 18564 31142
rect 18512 31078 18564 31084
rect 18616 26926 18644 37402
rect 18708 36582 18736 44474
rect 18696 36576 18748 36582
rect 18696 36518 18748 36524
rect 18696 34740 18748 34746
rect 18696 34682 18748 34688
rect 18708 33318 18736 34682
rect 18696 33312 18748 33318
rect 18696 33254 18748 33260
rect 18696 31952 18748 31958
rect 18696 31894 18748 31900
rect 18708 28762 18736 31894
rect 18696 28756 18748 28762
rect 18696 28698 18748 28704
rect 18604 26920 18656 26926
rect 18604 26862 18656 26868
rect 18604 24812 18656 24818
rect 18604 24754 18656 24760
rect 18616 22166 18644 24754
rect 18696 24200 18748 24206
rect 18696 24142 18748 24148
rect 18604 22160 18656 22166
rect 18604 22102 18656 22108
rect 18420 20052 18472 20058
rect 18420 19994 18472 20000
rect 18432 19446 18460 19994
rect 18512 19780 18564 19786
rect 18512 19722 18564 19728
rect 18420 19440 18472 19446
rect 18420 19382 18472 19388
rect 18420 18760 18472 18766
rect 18420 18702 18472 18708
rect 18432 17218 18460 18702
rect 18524 18442 18552 19722
rect 18616 18766 18644 22102
rect 18708 19786 18736 24142
rect 18696 19780 18748 19786
rect 18696 19722 18748 19728
rect 18696 19372 18748 19378
rect 18696 19314 18748 19320
rect 18708 18766 18736 19314
rect 18604 18760 18656 18766
rect 18604 18702 18656 18708
rect 18696 18760 18748 18766
rect 18696 18702 18748 18708
rect 18524 18414 18736 18442
rect 18432 17190 18644 17218
rect 18420 15156 18472 15162
rect 18420 15098 18472 15104
rect 18432 11082 18460 15098
rect 18420 11076 18472 11082
rect 18420 11018 18472 11024
rect 18248 6886 18368 6914
rect 17610 6556 17918 6565
rect 17610 6554 17616 6556
rect 17672 6554 17696 6556
rect 17752 6554 17776 6556
rect 17832 6554 17856 6556
rect 17912 6554 17918 6556
rect 17672 6502 17674 6554
rect 17854 6502 17856 6554
rect 17610 6500 17616 6502
rect 17672 6500 17696 6502
rect 17752 6500 17776 6502
rect 17832 6500 17856 6502
rect 17912 6500 17918 6502
rect 17610 6491 17918 6500
rect 17500 6384 17552 6390
rect 17500 6326 17552 6332
rect 17610 5468 17918 5477
rect 17610 5466 17616 5468
rect 17672 5466 17696 5468
rect 17752 5466 17776 5468
rect 17832 5466 17856 5468
rect 17912 5466 17918 5468
rect 17672 5414 17674 5466
rect 17854 5414 17856 5466
rect 17610 5412 17616 5414
rect 17672 5412 17696 5414
rect 17752 5412 17776 5414
rect 17832 5412 17856 5414
rect 17912 5412 17918 5414
rect 17610 5403 17918 5412
rect 18248 4554 18276 6886
rect 18616 4622 18644 17190
rect 18708 10674 18736 18414
rect 18696 10668 18748 10674
rect 18696 10610 18748 10616
rect 18800 6254 18828 61542
rect 18892 33454 18920 65962
rect 18984 37330 19012 66506
rect 19616 65408 19668 65414
rect 19616 65350 19668 65356
rect 19248 64456 19300 64462
rect 19248 64398 19300 64404
rect 19260 61266 19288 64398
rect 19248 61260 19300 61266
rect 19248 61202 19300 61208
rect 19628 60314 19656 65350
rect 19708 60512 19760 60518
rect 19708 60454 19760 60460
rect 19616 60308 19668 60314
rect 19616 60250 19668 60256
rect 19248 60104 19300 60110
rect 19248 60046 19300 60052
rect 19064 59424 19116 59430
rect 19064 59366 19116 59372
rect 19076 44538 19104 59366
rect 19260 58682 19288 60046
rect 19248 58676 19300 58682
rect 19248 58618 19300 58624
rect 19432 55888 19484 55894
rect 19432 55830 19484 55836
rect 19248 55752 19300 55758
rect 19248 55694 19300 55700
rect 19156 54188 19208 54194
rect 19156 54130 19208 54136
rect 19168 48142 19196 54130
rect 19260 49094 19288 55694
rect 19248 49088 19300 49094
rect 19248 49030 19300 49036
rect 19156 48136 19208 48142
rect 19156 48078 19208 48084
rect 19156 48000 19208 48006
rect 19156 47942 19208 47948
rect 19064 44532 19116 44538
rect 19064 44474 19116 44480
rect 19168 44418 19196 47942
rect 19076 44402 19196 44418
rect 19064 44396 19196 44402
rect 19116 44390 19196 44396
rect 19064 44338 19116 44344
rect 19156 44328 19208 44334
rect 19156 44270 19208 44276
rect 19168 42634 19196 44270
rect 19156 42628 19208 42634
rect 19156 42570 19208 42576
rect 18972 37324 19024 37330
rect 18972 37266 19024 37272
rect 19260 35562 19288 49030
rect 19444 44742 19472 55830
rect 19524 45008 19576 45014
rect 19524 44950 19576 44956
rect 19432 44736 19484 44742
rect 19432 44678 19484 44684
rect 19444 39438 19472 44678
rect 19536 42770 19564 44950
rect 19628 43994 19656 60250
rect 19720 59974 19748 60454
rect 19708 59968 19760 59974
rect 19708 59910 19760 59916
rect 19720 59430 19748 59910
rect 19708 59424 19760 59430
rect 19708 59366 19760 59372
rect 19812 56914 19840 68274
rect 20076 67040 20128 67046
rect 20076 66982 20128 66988
rect 19984 62892 20036 62898
rect 19984 62834 20036 62840
rect 19892 58540 19944 58546
rect 19892 58482 19944 58488
rect 19904 58002 19932 58482
rect 19892 57996 19944 58002
rect 19892 57938 19944 57944
rect 19800 56908 19852 56914
rect 19800 56850 19852 56856
rect 19812 44946 19840 56850
rect 19904 50522 19932 57938
rect 19996 56710 20024 62834
rect 20088 62218 20116 66982
rect 20180 64530 20208 68614
rect 21950 68028 22258 68037
rect 21950 68026 21956 68028
rect 22012 68026 22036 68028
rect 22092 68026 22116 68028
rect 22172 68026 22196 68028
rect 22252 68026 22258 68028
rect 22012 67974 22014 68026
rect 22194 67974 22196 68026
rect 21950 67972 21956 67974
rect 22012 67972 22036 67974
rect 22092 67972 22116 67974
rect 22172 67972 22196 67974
rect 22252 67972 22258 67974
rect 21950 67963 22258 67972
rect 20536 67584 20588 67590
rect 20536 67526 20588 67532
rect 20548 65618 20576 67526
rect 21950 66940 22258 66949
rect 21950 66938 21956 66940
rect 22012 66938 22036 66940
rect 22092 66938 22116 66940
rect 22172 66938 22196 66940
rect 22252 66938 22258 66940
rect 22012 66886 22014 66938
rect 22194 66886 22196 66938
rect 21950 66884 21956 66886
rect 22012 66884 22036 66886
rect 22092 66884 22116 66886
rect 22172 66884 22196 66886
rect 22252 66884 22258 66886
rect 21950 66875 22258 66884
rect 20628 66496 20680 66502
rect 20628 66438 20680 66444
rect 20536 65612 20588 65618
rect 20536 65554 20588 65560
rect 20640 64666 20668 66438
rect 21950 65852 22258 65861
rect 21950 65850 21956 65852
rect 22012 65850 22036 65852
rect 22092 65850 22116 65852
rect 22172 65850 22196 65852
rect 22252 65850 22258 65852
rect 22012 65798 22014 65850
rect 22194 65798 22196 65850
rect 21950 65796 21956 65798
rect 22012 65796 22036 65798
rect 22092 65796 22116 65798
rect 22172 65796 22196 65798
rect 22252 65796 22258 65798
rect 21950 65787 22258 65796
rect 21732 65612 21784 65618
rect 21732 65554 21784 65560
rect 20628 64660 20680 64666
rect 20628 64602 20680 64608
rect 20812 64660 20864 64666
rect 20812 64602 20864 64608
rect 20168 64524 20220 64530
rect 20168 64466 20220 64472
rect 20076 62212 20128 62218
rect 20076 62154 20128 62160
rect 20076 57928 20128 57934
rect 20076 57870 20128 57876
rect 19984 56704 20036 56710
rect 19984 56646 20036 56652
rect 19892 50516 19944 50522
rect 19892 50458 19944 50464
rect 19996 48822 20024 56646
rect 19984 48816 20036 48822
rect 19984 48758 20036 48764
rect 19996 45554 20024 48758
rect 19904 45526 20024 45554
rect 19800 44940 19852 44946
rect 19800 44882 19852 44888
rect 19616 43988 19668 43994
rect 19616 43930 19668 43936
rect 19628 43110 19656 43930
rect 19616 43104 19668 43110
rect 19616 43046 19668 43052
rect 19524 42764 19576 42770
rect 19524 42706 19576 42712
rect 19812 39438 19840 44882
rect 19904 42226 19932 45526
rect 19892 42220 19944 42226
rect 19892 42162 19944 42168
rect 19432 39432 19484 39438
rect 19432 39374 19484 39380
rect 19616 39432 19668 39438
rect 19616 39374 19668 39380
rect 19800 39432 19852 39438
rect 19800 39374 19852 39380
rect 19524 38548 19576 38554
rect 19524 38490 19576 38496
rect 19248 35556 19300 35562
rect 19248 35498 19300 35504
rect 19260 33658 19288 35498
rect 19248 33652 19300 33658
rect 19248 33594 19300 33600
rect 19340 33584 19392 33590
rect 19340 33526 19392 33532
rect 18880 33448 18932 33454
rect 18880 33390 18932 33396
rect 18892 31890 18920 33390
rect 19064 32564 19116 32570
rect 19064 32506 19116 32512
rect 19076 32298 19104 32506
rect 19248 32360 19300 32366
rect 19248 32302 19300 32308
rect 18972 32292 19024 32298
rect 18972 32234 19024 32240
rect 19064 32292 19116 32298
rect 19064 32234 19116 32240
rect 18880 31884 18932 31890
rect 18880 31826 18932 31832
rect 18984 26874 19012 32234
rect 18892 26846 19012 26874
rect 19156 26920 19208 26926
rect 19156 26862 19208 26868
rect 18892 17678 18920 26846
rect 18972 25832 19024 25838
rect 18972 25774 19024 25780
rect 18984 24274 19012 25774
rect 18972 24268 19024 24274
rect 18972 24210 19024 24216
rect 18984 19514 19012 24210
rect 19168 24070 19196 26862
rect 19260 26450 19288 32302
rect 19352 31958 19380 33526
rect 19340 31952 19392 31958
rect 19340 31894 19392 31900
rect 19248 26444 19300 26450
rect 19248 26386 19300 26392
rect 19536 25158 19564 38490
rect 19628 34474 19656 39374
rect 19800 38344 19852 38350
rect 19800 38286 19852 38292
rect 19616 34468 19668 34474
rect 19616 34410 19668 34416
rect 19812 28422 19840 38286
rect 19904 35222 19932 42162
rect 19984 41268 20036 41274
rect 19984 41210 20036 41216
rect 19892 35216 19944 35222
rect 19892 35158 19944 35164
rect 19904 33590 19932 35158
rect 19892 33584 19944 33590
rect 19892 33526 19944 33532
rect 19996 33386 20024 41210
rect 20088 36242 20116 57870
rect 20180 49298 20208 64466
rect 20352 64456 20404 64462
rect 20352 64398 20404 64404
rect 20720 64456 20772 64462
rect 20720 64398 20772 64404
rect 20260 64320 20312 64326
rect 20260 64262 20312 64268
rect 20168 49292 20220 49298
rect 20168 49234 20220 49240
rect 20180 45558 20208 49234
rect 20168 45552 20220 45558
rect 20168 45494 20220 45500
rect 20180 45286 20208 45494
rect 20168 45280 20220 45286
rect 20168 45222 20220 45228
rect 20166 38992 20222 39001
rect 20166 38927 20222 38936
rect 20180 38826 20208 38927
rect 20168 38820 20220 38826
rect 20168 38762 20220 38768
rect 20076 36236 20128 36242
rect 20076 36178 20128 36184
rect 19984 33380 20036 33386
rect 19984 33322 20036 33328
rect 19800 28416 19852 28422
rect 19800 28358 19852 28364
rect 19812 27674 19840 28358
rect 19800 27668 19852 27674
rect 19800 27610 19852 27616
rect 19524 25152 19576 25158
rect 19524 25094 19576 25100
rect 19156 24064 19208 24070
rect 19156 24006 19208 24012
rect 18972 19508 19024 19514
rect 18972 19450 19024 19456
rect 18880 17672 18932 17678
rect 18880 17614 18932 17620
rect 19168 13938 19196 24006
rect 19536 19990 19564 25094
rect 19996 24818 20024 33322
rect 19984 24812 20036 24818
rect 19984 24754 20036 24760
rect 19996 24698 20024 24754
rect 19812 24670 20024 24698
rect 19524 19984 19576 19990
rect 19524 19926 19576 19932
rect 19524 18624 19576 18630
rect 19524 18566 19576 18572
rect 19156 13932 19208 13938
rect 19156 13874 19208 13880
rect 19168 9110 19196 13874
rect 19156 9104 19208 9110
rect 19156 9046 19208 9052
rect 18788 6248 18840 6254
rect 18788 6190 18840 6196
rect 19536 4622 19564 18566
rect 19812 7410 19840 24670
rect 19984 24608 20036 24614
rect 19984 24550 20036 24556
rect 19892 23044 19944 23050
rect 19892 22986 19944 22992
rect 19800 7404 19852 7410
rect 19800 7346 19852 7352
rect 19904 7342 19932 22986
rect 19892 7336 19944 7342
rect 19892 7278 19944 7284
rect 19616 5092 19668 5098
rect 19616 5034 19668 5040
rect 18604 4616 18656 4622
rect 18604 4558 18656 4564
rect 19524 4616 19576 4622
rect 19524 4558 19576 4564
rect 19628 4554 19656 5034
rect 19996 4690 20024 24550
rect 20088 15162 20116 36178
rect 20076 15156 20128 15162
rect 20076 15098 20128 15104
rect 20272 8906 20300 64262
rect 20364 63617 20392 64398
rect 20732 64054 20760 64398
rect 20720 64048 20772 64054
rect 20720 63990 20772 63996
rect 20350 63608 20406 63617
rect 20350 63543 20406 63552
rect 20352 62212 20404 62218
rect 20352 62154 20404 62160
rect 20364 54194 20392 62154
rect 20824 60734 20852 64602
rect 21744 64462 21772 65554
rect 21950 64764 22258 64773
rect 21950 64762 21956 64764
rect 22012 64762 22036 64764
rect 22092 64762 22116 64764
rect 22172 64762 22196 64764
rect 22252 64762 22258 64764
rect 22012 64710 22014 64762
rect 22194 64710 22196 64762
rect 21950 64708 21956 64710
rect 22012 64708 22036 64710
rect 22092 64708 22116 64710
rect 22172 64708 22196 64710
rect 22252 64708 22258 64710
rect 21950 64699 22258 64708
rect 21088 64456 21140 64462
rect 21088 64398 21140 64404
rect 21732 64456 21784 64462
rect 21732 64398 21784 64404
rect 20904 62212 20956 62218
rect 20904 62154 20956 62160
rect 20732 60706 20852 60734
rect 20732 57934 20760 60706
rect 20812 58948 20864 58954
rect 20812 58890 20864 58896
rect 20720 57928 20772 57934
rect 20720 57870 20772 57876
rect 20732 57594 20760 57870
rect 20720 57588 20772 57594
rect 20720 57530 20772 57536
rect 20352 54188 20404 54194
rect 20352 54130 20404 54136
rect 20536 52556 20588 52562
rect 20536 52498 20588 52504
rect 20548 52086 20576 52498
rect 20536 52080 20588 52086
rect 20536 52022 20588 52028
rect 20626 52048 20682 52057
rect 20626 51983 20682 51992
rect 20640 51950 20668 51983
rect 20628 51944 20680 51950
rect 20824 51898 20852 58890
rect 20628 51886 20680 51892
rect 20732 51870 20852 51898
rect 20628 50448 20680 50454
rect 20628 50390 20680 50396
rect 20536 50312 20588 50318
rect 20536 50254 20588 50260
rect 20352 46436 20404 46442
rect 20352 46378 20404 46384
rect 20364 38894 20392 46378
rect 20444 39092 20496 39098
rect 20444 39034 20496 39040
rect 20456 38962 20484 39034
rect 20444 38956 20496 38962
rect 20444 38898 20496 38904
rect 20352 38888 20404 38894
rect 20350 38856 20352 38865
rect 20404 38856 20406 38865
rect 20350 38791 20406 38800
rect 20456 10742 20484 38898
rect 20548 24818 20576 50254
rect 20640 46510 20668 50390
rect 20628 46504 20680 46510
rect 20628 46446 20680 46452
rect 20732 31754 20760 51870
rect 20732 31726 20852 31754
rect 20720 28552 20772 28558
rect 20720 28494 20772 28500
rect 20628 27668 20680 27674
rect 20628 27610 20680 27616
rect 20536 24812 20588 24818
rect 20536 24754 20588 24760
rect 20640 20602 20668 27610
rect 20732 24750 20760 28494
rect 20824 27878 20852 31726
rect 20916 29714 20944 62154
rect 20996 57928 21048 57934
rect 20996 57870 21048 57876
rect 21008 52630 21036 57870
rect 20996 52624 21048 52630
rect 20996 52566 21048 52572
rect 20904 29708 20956 29714
rect 20904 29650 20956 29656
rect 20812 27872 20864 27878
rect 20812 27814 20864 27820
rect 20720 24744 20772 24750
rect 20720 24686 20772 24692
rect 20628 20596 20680 20602
rect 20628 20538 20680 20544
rect 21100 18834 21128 64398
rect 21744 63617 21772 64398
rect 21950 63676 22258 63685
rect 21950 63674 21956 63676
rect 22012 63674 22036 63676
rect 22092 63674 22116 63676
rect 22172 63674 22196 63676
rect 22252 63674 22258 63676
rect 22012 63622 22014 63674
rect 22194 63622 22196 63674
rect 21950 63620 21956 63622
rect 22012 63620 22036 63622
rect 22092 63620 22116 63622
rect 22172 63620 22196 63622
rect 22252 63620 22258 63622
rect 21730 63608 21786 63617
rect 21950 63611 22258 63620
rect 21730 63543 21786 63552
rect 22388 63442 22416 69294
rect 26950 69116 27258 69125
rect 26950 69114 26956 69116
rect 27012 69114 27036 69116
rect 27092 69114 27116 69116
rect 27172 69114 27196 69116
rect 27252 69114 27258 69116
rect 27012 69062 27014 69114
rect 27194 69062 27196 69114
rect 26950 69060 26956 69062
rect 27012 69060 27036 69062
rect 27092 69060 27116 69062
rect 27172 69060 27196 69062
rect 27252 69060 27258 69062
rect 26950 69051 27258 69060
rect 31950 69116 32258 69125
rect 31950 69114 31956 69116
rect 32012 69114 32036 69116
rect 32092 69114 32116 69116
rect 32172 69114 32196 69116
rect 32252 69114 32258 69116
rect 32012 69062 32014 69114
rect 32194 69062 32196 69114
rect 31950 69060 31956 69062
rect 32012 69060 32036 69062
rect 32092 69060 32116 69062
rect 32172 69060 32196 69062
rect 32252 69060 32258 69062
rect 31950 69051 32258 69060
rect 28724 68808 28776 68814
rect 28724 68750 28776 68756
rect 31484 68808 31536 68814
rect 31484 68750 31536 68756
rect 22610 68572 22918 68581
rect 22610 68570 22616 68572
rect 22672 68570 22696 68572
rect 22752 68570 22776 68572
rect 22832 68570 22856 68572
rect 22912 68570 22918 68572
rect 22672 68518 22674 68570
rect 22854 68518 22856 68570
rect 22610 68516 22616 68518
rect 22672 68516 22696 68518
rect 22752 68516 22776 68518
rect 22832 68516 22856 68518
rect 22912 68516 22918 68518
rect 22610 68507 22918 68516
rect 27610 68572 27918 68581
rect 27610 68570 27616 68572
rect 27672 68570 27696 68572
rect 27752 68570 27776 68572
rect 27832 68570 27856 68572
rect 27912 68570 27918 68572
rect 27672 68518 27674 68570
rect 27854 68518 27856 68570
rect 27610 68516 27616 68518
rect 27672 68516 27696 68518
rect 27752 68516 27776 68518
rect 27832 68516 27856 68518
rect 27912 68516 27918 68518
rect 27610 68507 27918 68516
rect 23848 68400 23900 68406
rect 23848 68342 23900 68348
rect 23112 68332 23164 68338
rect 23112 68274 23164 68280
rect 22610 67484 22918 67493
rect 22610 67482 22616 67484
rect 22672 67482 22696 67484
rect 22752 67482 22776 67484
rect 22832 67482 22856 67484
rect 22912 67482 22918 67484
rect 22672 67430 22674 67482
rect 22854 67430 22856 67482
rect 22610 67428 22616 67430
rect 22672 67428 22696 67430
rect 22752 67428 22776 67430
rect 22832 67428 22856 67430
rect 22912 67428 22918 67430
rect 22610 67419 22918 67428
rect 22610 66396 22918 66405
rect 22610 66394 22616 66396
rect 22672 66394 22696 66396
rect 22752 66394 22776 66396
rect 22832 66394 22856 66396
rect 22912 66394 22918 66396
rect 22672 66342 22674 66394
rect 22854 66342 22856 66394
rect 22610 66340 22616 66342
rect 22672 66340 22696 66342
rect 22752 66340 22776 66342
rect 22832 66340 22856 66342
rect 22912 66340 22918 66342
rect 22610 66331 22918 66340
rect 22610 65308 22918 65317
rect 22610 65306 22616 65308
rect 22672 65306 22696 65308
rect 22752 65306 22776 65308
rect 22832 65306 22856 65308
rect 22912 65306 22918 65308
rect 22672 65254 22674 65306
rect 22854 65254 22856 65306
rect 22610 65252 22616 65254
rect 22672 65252 22696 65254
rect 22752 65252 22776 65254
rect 22832 65252 22856 65254
rect 22912 65252 22918 65254
rect 22610 65243 22918 65252
rect 23124 64874 23152 68274
rect 23296 67244 23348 67250
rect 23296 67186 23348 67192
rect 23032 64846 23152 64874
rect 22610 64220 22918 64229
rect 22610 64218 22616 64220
rect 22672 64218 22696 64220
rect 22752 64218 22776 64220
rect 22832 64218 22856 64220
rect 22912 64218 22918 64220
rect 22672 64166 22674 64218
rect 22854 64166 22856 64218
rect 22610 64164 22616 64166
rect 22672 64164 22696 64166
rect 22752 64164 22776 64166
rect 22832 64164 22856 64166
rect 22912 64164 22918 64166
rect 22610 64155 22918 64164
rect 22376 63436 22428 63442
rect 22376 63378 22428 63384
rect 21950 62588 22258 62597
rect 21950 62586 21956 62588
rect 22012 62586 22036 62588
rect 22092 62586 22116 62588
rect 22172 62586 22196 62588
rect 22252 62586 22258 62588
rect 22012 62534 22014 62586
rect 22194 62534 22196 62586
rect 21950 62532 21956 62534
rect 22012 62532 22036 62534
rect 22092 62532 22116 62534
rect 22172 62532 22196 62534
rect 22252 62532 22258 62534
rect 21950 62523 22258 62532
rect 21950 61500 22258 61509
rect 21950 61498 21956 61500
rect 22012 61498 22036 61500
rect 22092 61498 22116 61500
rect 22172 61498 22196 61500
rect 22252 61498 22258 61500
rect 22012 61446 22014 61498
rect 22194 61446 22196 61498
rect 21950 61444 21956 61446
rect 22012 61444 22036 61446
rect 22092 61444 22116 61446
rect 22172 61444 22196 61446
rect 22252 61444 22258 61446
rect 21950 61435 22258 61444
rect 21950 60412 22258 60421
rect 21950 60410 21956 60412
rect 22012 60410 22036 60412
rect 22092 60410 22116 60412
rect 22172 60410 22196 60412
rect 22252 60410 22258 60412
rect 22012 60358 22014 60410
rect 22194 60358 22196 60410
rect 21950 60356 21956 60358
rect 22012 60356 22036 60358
rect 22092 60356 22116 60358
rect 22172 60356 22196 60358
rect 22252 60356 22258 60358
rect 21950 60347 22258 60356
rect 22100 60104 22152 60110
rect 22100 60046 22152 60052
rect 21272 60036 21324 60042
rect 21272 59978 21324 59984
rect 21284 59702 21312 59978
rect 21272 59696 21324 59702
rect 21272 59638 21324 59644
rect 21180 42628 21232 42634
rect 21180 42570 21232 42576
rect 21088 18828 21140 18834
rect 21088 18770 21140 18776
rect 21100 11218 21128 18770
rect 21088 11212 21140 11218
rect 21088 11154 21140 11160
rect 21192 11014 21220 42570
rect 21284 41414 21312 59638
rect 22112 59537 22140 60046
rect 22098 59528 22154 59537
rect 22098 59463 22154 59472
rect 21364 59424 21416 59430
rect 21364 59366 21416 59372
rect 21376 45014 21404 59366
rect 21950 59324 22258 59333
rect 21950 59322 21956 59324
rect 22012 59322 22036 59324
rect 22092 59322 22116 59324
rect 22172 59322 22196 59324
rect 22252 59322 22258 59324
rect 22012 59270 22014 59322
rect 22194 59270 22196 59322
rect 21950 59268 21956 59270
rect 22012 59268 22036 59270
rect 22092 59268 22116 59270
rect 22172 59268 22196 59270
rect 22252 59268 22258 59270
rect 21950 59259 22258 59268
rect 22388 59090 22416 63378
rect 22610 63132 22918 63141
rect 22610 63130 22616 63132
rect 22672 63130 22696 63132
rect 22752 63130 22776 63132
rect 22832 63130 22856 63132
rect 22912 63130 22918 63132
rect 22672 63078 22674 63130
rect 22854 63078 22856 63130
rect 22610 63076 22616 63078
rect 22672 63076 22696 63078
rect 22752 63076 22776 63078
rect 22832 63076 22856 63078
rect 22912 63076 22918 63078
rect 22610 63067 22918 63076
rect 22610 62044 22918 62053
rect 22610 62042 22616 62044
rect 22672 62042 22696 62044
rect 22752 62042 22776 62044
rect 22832 62042 22856 62044
rect 22912 62042 22918 62044
rect 22672 61990 22674 62042
rect 22854 61990 22856 62042
rect 22610 61988 22616 61990
rect 22672 61988 22696 61990
rect 22752 61988 22776 61990
rect 22832 61988 22856 61990
rect 22912 61988 22918 61990
rect 22610 61979 22918 61988
rect 22610 60956 22918 60965
rect 22610 60954 22616 60956
rect 22672 60954 22696 60956
rect 22752 60954 22776 60956
rect 22832 60954 22856 60956
rect 22912 60954 22918 60956
rect 22672 60902 22674 60954
rect 22854 60902 22856 60954
rect 22610 60900 22616 60902
rect 22672 60900 22696 60902
rect 22752 60900 22776 60902
rect 22832 60900 22856 60902
rect 22912 60900 22918 60902
rect 22610 60891 22918 60900
rect 22468 59968 22520 59974
rect 22468 59910 22520 59916
rect 22376 59084 22428 59090
rect 22376 59026 22428 59032
rect 22284 59016 22336 59022
rect 22284 58958 22336 58964
rect 21950 58236 22258 58245
rect 21950 58234 21956 58236
rect 22012 58234 22036 58236
rect 22092 58234 22116 58236
rect 22172 58234 22196 58236
rect 22252 58234 22258 58236
rect 22012 58182 22014 58234
rect 22194 58182 22196 58234
rect 21950 58180 21956 58182
rect 22012 58180 22036 58182
rect 22092 58180 22116 58182
rect 22172 58180 22196 58182
rect 22252 58180 22258 58182
rect 21950 58171 22258 58180
rect 21548 57452 21600 57458
rect 21548 57394 21600 57400
rect 21560 54262 21588 57394
rect 22296 57322 22324 58958
rect 22376 57384 22428 57390
rect 22376 57326 22428 57332
rect 22284 57316 22336 57322
rect 22284 57258 22336 57264
rect 21950 57148 22258 57157
rect 21950 57146 21956 57148
rect 22012 57146 22036 57148
rect 22092 57146 22116 57148
rect 22172 57146 22196 57148
rect 22252 57146 22258 57148
rect 22012 57094 22014 57146
rect 22194 57094 22196 57146
rect 21950 57092 21956 57094
rect 22012 57092 22036 57094
rect 22092 57092 22116 57094
rect 22172 57092 22196 57094
rect 22252 57092 22258 57094
rect 21950 57083 22258 57092
rect 22388 56250 22416 57326
rect 22296 56222 22416 56250
rect 21950 56060 22258 56069
rect 21950 56058 21956 56060
rect 22012 56058 22036 56060
rect 22092 56058 22116 56060
rect 22172 56058 22196 56060
rect 22252 56058 22258 56060
rect 22012 56006 22014 56058
rect 22194 56006 22196 56058
rect 21950 56004 21956 56006
rect 22012 56004 22036 56006
rect 22092 56004 22116 56006
rect 22172 56004 22196 56006
rect 22252 56004 22258 56006
rect 21950 55995 22258 56004
rect 21950 54972 22258 54981
rect 21950 54970 21956 54972
rect 22012 54970 22036 54972
rect 22092 54970 22116 54972
rect 22172 54970 22196 54972
rect 22252 54970 22258 54972
rect 22012 54918 22014 54970
rect 22194 54918 22196 54970
rect 21950 54916 21956 54918
rect 22012 54916 22036 54918
rect 22092 54916 22116 54918
rect 22172 54916 22196 54918
rect 22252 54916 22258 54918
rect 21950 54907 22258 54916
rect 21548 54256 21600 54262
rect 21548 54198 21600 54204
rect 21456 52080 21508 52086
rect 21454 52048 21456 52057
rect 21508 52048 21510 52057
rect 21560 52018 21588 54198
rect 21950 53884 22258 53893
rect 21950 53882 21956 53884
rect 22012 53882 22036 53884
rect 22092 53882 22116 53884
rect 22172 53882 22196 53884
rect 22252 53882 22258 53884
rect 22012 53830 22014 53882
rect 22194 53830 22196 53882
rect 21950 53828 21956 53830
rect 22012 53828 22036 53830
rect 22092 53828 22116 53830
rect 22172 53828 22196 53830
rect 22252 53828 22258 53830
rect 21950 53819 22258 53828
rect 21732 53168 21784 53174
rect 21732 53110 21784 53116
rect 21744 52494 21772 53110
rect 21950 52796 22258 52805
rect 21950 52794 21956 52796
rect 22012 52794 22036 52796
rect 22092 52794 22116 52796
rect 22172 52794 22196 52796
rect 22252 52794 22258 52796
rect 22012 52742 22014 52794
rect 22194 52742 22196 52794
rect 21950 52740 21956 52742
rect 22012 52740 22036 52742
rect 22092 52740 22116 52742
rect 22172 52740 22196 52742
rect 22252 52740 22258 52742
rect 21950 52731 22258 52740
rect 21732 52488 21784 52494
rect 21732 52430 21784 52436
rect 21640 52148 21692 52154
rect 21640 52090 21692 52096
rect 21454 51983 21510 51992
rect 21548 52012 21600 52018
rect 21548 51954 21600 51960
rect 21652 51950 21680 52090
rect 21640 51944 21692 51950
rect 21640 51886 21692 51892
rect 21744 51814 21772 52430
rect 21732 51808 21784 51814
rect 21732 51750 21784 51756
rect 21950 51708 22258 51717
rect 21950 51706 21956 51708
rect 22012 51706 22036 51708
rect 22092 51706 22116 51708
rect 22172 51706 22196 51708
rect 22252 51706 22258 51708
rect 22012 51654 22014 51706
rect 22194 51654 22196 51706
rect 21950 51652 21956 51654
rect 22012 51652 22036 51654
rect 22092 51652 22116 51654
rect 22172 51652 22196 51654
rect 22252 51652 22258 51654
rect 21950 51643 22258 51652
rect 22296 51066 22324 56222
rect 22376 55820 22428 55826
rect 22376 55762 22428 55768
rect 22284 51060 22336 51066
rect 22284 51002 22336 51008
rect 22388 50998 22416 55762
rect 22376 50992 22428 50998
rect 22376 50934 22428 50940
rect 21824 50924 21876 50930
rect 21824 50866 21876 50872
rect 22284 50924 22336 50930
rect 22284 50866 22336 50872
rect 21732 50856 21784 50862
rect 21732 50798 21784 50804
rect 21364 45008 21416 45014
rect 21364 44950 21416 44956
rect 21548 42832 21600 42838
rect 21548 42774 21600 42780
rect 21284 41386 21496 41414
rect 21364 40724 21416 40730
rect 21364 40666 21416 40672
rect 21376 12238 21404 40666
rect 21468 39370 21496 41386
rect 21560 41206 21588 42774
rect 21744 41414 21772 50798
rect 21836 47666 21864 50866
rect 21950 50620 22258 50629
rect 21950 50618 21956 50620
rect 22012 50618 22036 50620
rect 22092 50618 22116 50620
rect 22172 50618 22196 50620
rect 22252 50618 22258 50620
rect 22012 50566 22014 50618
rect 22194 50566 22196 50618
rect 21950 50564 21956 50566
rect 22012 50564 22036 50566
rect 22092 50564 22116 50566
rect 22172 50564 22196 50566
rect 22252 50564 22258 50566
rect 21950 50555 22258 50564
rect 21950 49532 22258 49541
rect 21950 49530 21956 49532
rect 22012 49530 22036 49532
rect 22092 49530 22116 49532
rect 22172 49530 22196 49532
rect 22252 49530 22258 49532
rect 22012 49478 22014 49530
rect 22194 49478 22196 49530
rect 21950 49476 21956 49478
rect 22012 49476 22036 49478
rect 22092 49476 22116 49478
rect 22172 49476 22196 49478
rect 22252 49476 22258 49478
rect 21950 49467 22258 49476
rect 22296 49366 22324 50866
rect 22388 49774 22416 50934
rect 22376 49768 22428 49774
rect 22376 49710 22428 49716
rect 22284 49360 22336 49366
rect 22284 49302 22336 49308
rect 22376 48748 22428 48754
rect 22376 48690 22428 48696
rect 22284 48544 22336 48550
rect 22284 48486 22336 48492
rect 21950 48444 22258 48453
rect 21950 48442 21956 48444
rect 22012 48442 22036 48444
rect 22092 48442 22116 48444
rect 22172 48442 22196 48444
rect 22252 48442 22258 48444
rect 22012 48390 22014 48442
rect 22194 48390 22196 48442
rect 21950 48388 21956 48390
rect 22012 48388 22036 48390
rect 22092 48388 22116 48390
rect 22172 48388 22196 48390
rect 22252 48388 22258 48390
rect 21950 48379 22258 48388
rect 21824 47660 21876 47666
rect 21824 47602 21876 47608
rect 21950 47356 22258 47365
rect 21950 47354 21956 47356
rect 22012 47354 22036 47356
rect 22092 47354 22116 47356
rect 22172 47354 22196 47356
rect 22252 47354 22258 47356
rect 22012 47302 22014 47354
rect 22194 47302 22196 47354
rect 21950 47300 21956 47302
rect 22012 47300 22036 47302
rect 22092 47300 22116 47302
rect 22172 47300 22196 47302
rect 22252 47300 22258 47302
rect 21950 47291 22258 47300
rect 21950 46268 22258 46277
rect 21950 46266 21956 46268
rect 22012 46266 22036 46268
rect 22092 46266 22116 46268
rect 22172 46266 22196 46268
rect 22252 46266 22258 46268
rect 22012 46214 22014 46266
rect 22194 46214 22196 46266
rect 21950 46212 21956 46214
rect 22012 46212 22036 46214
rect 22092 46212 22116 46214
rect 22172 46212 22196 46214
rect 22252 46212 22258 46214
rect 21950 46203 22258 46212
rect 21950 45180 22258 45189
rect 21950 45178 21956 45180
rect 22012 45178 22036 45180
rect 22092 45178 22116 45180
rect 22172 45178 22196 45180
rect 22252 45178 22258 45180
rect 22012 45126 22014 45178
rect 22194 45126 22196 45178
rect 21950 45124 21956 45126
rect 22012 45124 22036 45126
rect 22092 45124 22116 45126
rect 22172 45124 22196 45126
rect 22252 45124 22258 45126
rect 21950 45115 22258 45124
rect 21950 44092 22258 44101
rect 21950 44090 21956 44092
rect 22012 44090 22036 44092
rect 22092 44090 22116 44092
rect 22172 44090 22196 44092
rect 22252 44090 22258 44092
rect 22012 44038 22014 44090
rect 22194 44038 22196 44090
rect 21950 44036 21956 44038
rect 22012 44036 22036 44038
rect 22092 44036 22116 44038
rect 22172 44036 22196 44038
rect 22252 44036 22258 44038
rect 21950 44027 22258 44036
rect 21950 43004 22258 43013
rect 21950 43002 21956 43004
rect 22012 43002 22036 43004
rect 22092 43002 22116 43004
rect 22172 43002 22196 43004
rect 22252 43002 22258 43004
rect 22012 42950 22014 43002
rect 22194 42950 22196 43002
rect 21950 42948 21956 42950
rect 22012 42948 22036 42950
rect 22092 42948 22116 42950
rect 22172 42948 22196 42950
rect 22252 42948 22258 42950
rect 21950 42939 22258 42948
rect 22192 42900 22244 42906
rect 22192 42842 22244 42848
rect 22098 42800 22154 42809
rect 22098 42735 22154 42744
rect 22112 42702 22140 42735
rect 22100 42696 22152 42702
rect 22100 42638 22152 42644
rect 22204 42106 22232 42842
rect 22296 42770 22324 48486
rect 22388 46578 22416 48690
rect 22376 46572 22428 46578
rect 22376 46514 22428 46520
rect 22376 46436 22428 46442
rect 22376 46378 22428 46384
rect 22388 44878 22416 46378
rect 22376 44872 22428 44878
rect 22376 44814 22428 44820
rect 22284 42764 22336 42770
rect 22284 42706 22336 42712
rect 22388 42650 22416 44814
rect 22480 42809 22508 59910
rect 22610 59868 22918 59877
rect 22610 59866 22616 59868
rect 22672 59866 22696 59868
rect 22752 59866 22776 59868
rect 22832 59866 22856 59868
rect 22912 59866 22918 59868
rect 22672 59814 22674 59866
rect 22854 59814 22856 59866
rect 22610 59812 22616 59814
rect 22672 59812 22696 59814
rect 22752 59812 22776 59814
rect 22832 59812 22856 59814
rect 22912 59812 22918 59814
rect 22610 59803 22918 59812
rect 22610 58780 22918 58789
rect 22610 58778 22616 58780
rect 22672 58778 22696 58780
rect 22752 58778 22776 58780
rect 22832 58778 22856 58780
rect 22912 58778 22918 58780
rect 22672 58726 22674 58778
rect 22854 58726 22856 58778
rect 22610 58724 22616 58726
rect 22672 58724 22696 58726
rect 22752 58724 22776 58726
rect 22832 58724 22856 58726
rect 22912 58724 22918 58726
rect 22610 58715 22918 58724
rect 22610 57692 22918 57701
rect 22610 57690 22616 57692
rect 22672 57690 22696 57692
rect 22752 57690 22776 57692
rect 22832 57690 22856 57692
rect 22912 57690 22918 57692
rect 22672 57638 22674 57690
rect 22854 57638 22856 57690
rect 22610 57636 22616 57638
rect 22672 57636 22696 57638
rect 22752 57636 22776 57638
rect 22832 57636 22856 57638
rect 22912 57636 22918 57638
rect 22610 57627 22918 57636
rect 22610 56604 22918 56613
rect 22610 56602 22616 56604
rect 22672 56602 22696 56604
rect 22752 56602 22776 56604
rect 22832 56602 22856 56604
rect 22912 56602 22918 56604
rect 22672 56550 22674 56602
rect 22854 56550 22856 56602
rect 22610 56548 22616 56550
rect 22672 56548 22696 56550
rect 22752 56548 22776 56550
rect 22832 56548 22856 56550
rect 22912 56548 22918 56550
rect 22610 56539 22918 56548
rect 22610 55516 22918 55525
rect 22610 55514 22616 55516
rect 22672 55514 22696 55516
rect 22752 55514 22776 55516
rect 22832 55514 22856 55516
rect 22912 55514 22918 55516
rect 22672 55462 22674 55514
rect 22854 55462 22856 55514
rect 22610 55460 22616 55462
rect 22672 55460 22696 55462
rect 22752 55460 22776 55462
rect 22832 55460 22856 55462
rect 22912 55460 22918 55462
rect 22610 55451 22918 55460
rect 22610 54428 22918 54437
rect 22610 54426 22616 54428
rect 22672 54426 22696 54428
rect 22752 54426 22776 54428
rect 22832 54426 22856 54428
rect 22912 54426 22918 54428
rect 22672 54374 22674 54426
rect 22854 54374 22856 54426
rect 22610 54372 22616 54374
rect 22672 54372 22696 54374
rect 22752 54372 22776 54374
rect 22832 54372 22856 54374
rect 22912 54372 22918 54374
rect 22610 54363 22918 54372
rect 22610 53340 22918 53349
rect 22610 53338 22616 53340
rect 22672 53338 22696 53340
rect 22752 53338 22776 53340
rect 22832 53338 22856 53340
rect 22912 53338 22918 53340
rect 22672 53286 22674 53338
rect 22854 53286 22856 53338
rect 22610 53284 22616 53286
rect 22672 53284 22696 53286
rect 22752 53284 22776 53286
rect 22832 53284 22856 53286
rect 22912 53284 22918 53286
rect 22610 53275 22918 53284
rect 22610 52252 22918 52261
rect 22610 52250 22616 52252
rect 22672 52250 22696 52252
rect 22752 52250 22776 52252
rect 22832 52250 22856 52252
rect 22912 52250 22918 52252
rect 22672 52198 22674 52250
rect 22854 52198 22856 52250
rect 22610 52196 22616 52198
rect 22672 52196 22696 52198
rect 22752 52196 22776 52198
rect 22832 52196 22856 52198
rect 22912 52196 22918 52198
rect 22610 52187 22918 52196
rect 22610 51164 22918 51173
rect 22610 51162 22616 51164
rect 22672 51162 22696 51164
rect 22752 51162 22776 51164
rect 22832 51162 22856 51164
rect 22912 51162 22918 51164
rect 22672 51110 22674 51162
rect 22854 51110 22856 51162
rect 22610 51108 22616 51110
rect 22672 51108 22696 51110
rect 22752 51108 22776 51110
rect 22832 51108 22856 51110
rect 22912 51108 22918 51110
rect 22610 51099 22918 51108
rect 22610 50076 22918 50085
rect 22610 50074 22616 50076
rect 22672 50074 22696 50076
rect 22752 50074 22776 50076
rect 22832 50074 22856 50076
rect 22912 50074 22918 50076
rect 22672 50022 22674 50074
rect 22854 50022 22856 50074
rect 22610 50020 22616 50022
rect 22672 50020 22696 50022
rect 22752 50020 22776 50022
rect 22832 50020 22856 50022
rect 22912 50020 22918 50022
rect 22610 50011 22918 50020
rect 22610 48988 22918 48997
rect 22610 48986 22616 48988
rect 22672 48986 22696 48988
rect 22752 48986 22776 48988
rect 22832 48986 22856 48988
rect 22912 48986 22918 48988
rect 22672 48934 22674 48986
rect 22854 48934 22856 48986
rect 22610 48932 22616 48934
rect 22672 48932 22696 48934
rect 22752 48932 22776 48934
rect 22832 48932 22856 48934
rect 22912 48932 22918 48934
rect 22610 48923 22918 48932
rect 22610 47900 22918 47909
rect 22610 47898 22616 47900
rect 22672 47898 22696 47900
rect 22752 47898 22776 47900
rect 22832 47898 22856 47900
rect 22912 47898 22918 47900
rect 22672 47846 22674 47898
rect 22854 47846 22856 47898
rect 22610 47844 22616 47846
rect 22672 47844 22696 47846
rect 22752 47844 22776 47846
rect 22832 47844 22856 47846
rect 22912 47844 22918 47846
rect 22610 47835 22918 47844
rect 22610 46812 22918 46821
rect 22610 46810 22616 46812
rect 22672 46810 22696 46812
rect 22752 46810 22776 46812
rect 22832 46810 22856 46812
rect 22912 46810 22918 46812
rect 22672 46758 22674 46810
rect 22854 46758 22856 46810
rect 22610 46756 22616 46758
rect 22672 46756 22696 46758
rect 22752 46756 22776 46758
rect 22832 46756 22856 46758
rect 22912 46756 22918 46758
rect 22610 46747 22918 46756
rect 23032 46442 23060 64846
rect 23204 62144 23256 62150
rect 23204 62086 23256 62092
rect 23112 60104 23164 60110
rect 23112 60046 23164 60052
rect 23124 53446 23152 60046
rect 23216 55826 23244 62086
rect 23204 55820 23256 55826
rect 23204 55762 23256 55768
rect 23112 53440 23164 53446
rect 23112 53382 23164 53388
rect 23112 51060 23164 51066
rect 23112 51002 23164 51008
rect 23124 49978 23152 51002
rect 23204 50720 23256 50726
rect 23204 50662 23256 50668
rect 23112 49972 23164 49978
rect 23112 49914 23164 49920
rect 23112 49768 23164 49774
rect 23112 49710 23164 49716
rect 23020 46436 23072 46442
rect 23020 46378 23072 46384
rect 23020 46164 23072 46170
rect 23020 46106 23072 46112
rect 22610 45724 22918 45733
rect 22610 45722 22616 45724
rect 22672 45722 22696 45724
rect 22752 45722 22776 45724
rect 22832 45722 22856 45724
rect 22912 45722 22918 45724
rect 22672 45670 22674 45722
rect 22854 45670 22856 45722
rect 22610 45668 22616 45670
rect 22672 45668 22696 45670
rect 22752 45668 22776 45670
rect 22832 45668 22856 45670
rect 22912 45668 22918 45670
rect 22610 45659 22918 45668
rect 22610 44636 22918 44645
rect 22610 44634 22616 44636
rect 22672 44634 22696 44636
rect 22752 44634 22776 44636
rect 22832 44634 22856 44636
rect 22912 44634 22918 44636
rect 22672 44582 22674 44634
rect 22854 44582 22856 44634
rect 22610 44580 22616 44582
rect 22672 44580 22696 44582
rect 22752 44580 22776 44582
rect 22832 44580 22856 44582
rect 22912 44580 22918 44582
rect 22610 44571 22918 44580
rect 22610 43548 22918 43557
rect 22610 43546 22616 43548
rect 22672 43546 22696 43548
rect 22752 43546 22776 43548
rect 22832 43546 22856 43548
rect 22912 43546 22918 43548
rect 22672 43494 22674 43546
rect 22854 43494 22856 43546
rect 22610 43492 22616 43494
rect 22672 43492 22696 43494
rect 22752 43492 22776 43494
rect 22832 43492 22856 43494
rect 22912 43492 22918 43494
rect 22610 43483 22918 43492
rect 22466 42800 22522 42809
rect 22466 42735 22522 42744
rect 22744 42764 22796 42770
rect 22744 42706 22796 42712
rect 22388 42622 22508 42650
rect 22376 42560 22428 42566
rect 22376 42502 22428 42508
rect 22388 42226 22416 42502
rect 22376 42220 22428 42226
rect 22376 42162 22428 42168
rect 22204 42078 22324 42106
rect 21950 41916 22258 41925
rect 21950 41914 21956 41916
rect 22012 41914 22036 41916
rect 22092 41914 22116 41916
rect 22172 41914 22196 41916
rect 22252 41914 22258 41916
rect 22012 41862 22014 41914
rect 22194 41862 22196 41914
rect 21950 41860 21956 41862
rect 22012 41860 22036 41862
rect 22092 41860 22116 41862
rect 22172 41860 22196 41862
rect 22252 41860 22258 41862
rect 21950 41851 22258 41860
rect 21744 41386 21864 41414
rect 21548 41200 21600 41206
rect 21548 41142 21600 41148
rect 21456 39364 21508 39370
rect 21456 39306 21508 39312
rect 21468 12850 21496 39306
rect 21836 34762 21864 41386
rect 21950 40828 22258 40837
rect 21950 40826 21956 40828
rect 22012 40826 22036 40828
rect 22092 40826 22116 40828
rect 22172 40826 22196 40828
rect 22252 40826 22258 40828
rect 22012 40774 22014 40826
rect 22194 40774 22196 40826
rect 21950 40772 21956 40774
rect 22012 40772 22036 40774
rect 22092 40772 22116 40774
rect 22172 40772 22196 40774
rect 22252 40772 22258 40774
rect 21950 40763 22258 40772
rect 21950 39740 22258 39749
rect 21950 39738 21956 39740
rect 22012 39738 22036 39740
rect 22092 39738 22116 39740
rect 22172 39738 22196 39740
rect 22252 39738 22258 39740
rect 22012 39686 22014 39738
rect 22194 39686 22196 39738
rect 21950 39684 21956 39686
rect 22012 39684 22036 39686
rect 22092 39684 22116 39686
rect 22172 39684 22196 39686
rect 22252 39684 22258 39686
rect 21950 39675 22258 39684
rect 22190 39400 22246 39409
rect 22190 39335 22246 39344
rect 22204 39302 22232 39335
rect 22192 39296 22244 39302
rect 22192 39238 22244 39244
rect 21950 38652 22258 38661
rect 21950 38650 21956 38652
rect 22012 38650 22036 38652
rect 22092 38650 22116 38652
rect 22172 38650 22196 38652
rect 22252 38650 22258 38652
rect 22012 38598 22014 38650
rect 22194 38598 22196 38650
rect 21950 38596 21956 38598
rect 22012 38596 22036 38598
rect 22092 38596 22116 38598
rect 22172 38596 22196 38598
rect 22252 38596 22258 38598
rect 21950 38587 22258 38596
rect 21950 37564 22258 37573
rect 21950 37562 21956 37564
rect 22012 37562 22036 37564
rect 22092 37562 22116 37564
rect 22172 37562 22196 37564
rect 22252 37562 22258 37564
rect 22012 37510 22014 37562
rect 22194 37510 22196 37562
rect 21950 37508 21956 37510
rect 22012 37508 22036 37510
rect 22092 37508 22116 37510
rect 22172 37508 22196 37510
rect 22252 37508 22258 37510
rect 21950 37499 22258 37508
rect 21950 36476 22258 36485
rect 21950 36474 21956 36476
rect 22012 36474 22036 36476
rect 22092 36474 22116 36476
rect 22172 36474 22196 36476
rect 22252 36474 22258 36476
rect 22012 36422 22014 36474
rect 22194 36422 22196 36474
rect 21950 36420 21956 36422
rect 22012 36420 22036 36422
rect 22092 36420 22116 36422
rect 22172 36420 22196 36422
rect 22252 36420 22258 36422
rect 21950 36411 22258 36420
rect 21950 35388 22258 35397
rect 21950 35386 21956 35388
rect 22012 35386 22036 35388
rect 22092 35386 22116 35388
rect 22172 35386 22196 35388
rect 22252 35386 22258 35388
rect 22012 35334 22014 35386
rect 22194 35334 22196 35386
rect 21950 35332 21956 35334
rect 22012 35332 22036 35334
rect 22092 35332 22116 35334
rect 22172 35332 22196 35334
rect 22252 35332 22258 35334
rect 21950 35323 22258 35332
rect 21652 34734 21864 34762
rect 21652 34610 21680 34734
rect 21640 34604 21692 34610
rect 21640 34546 21692 34552
rect 21732 34604 21784 34610
rect 21732 34546 21784 34552
rect 21640 29640 21692 29646
rect 21640 29582 21692 29588
rect 21548 27872 21600 27878
rect 21548 27814 21600 27820
rect 21456 12844 21508 12850
rect 21456 12786 21508 12792
rect 21560 12306 21588 27814
rect 21652 13190 21680 29582
rect 21744 23322 21772 34546
rect 21836 34134 21864 34734
rect 21950 34300 22258 34309
rect 21950 34298 21956 34300
rect 22012 34298 22036 34300
rect 22092 34298 22116 34300
rect 22172 34298 22196 34300
rect 22252 34298 22258 34300
rect 22012 34246 22014 34298
rect 22194 34246 22196 34298
rect 21950 34244 21956 34246
rect 22012 34244 22036 34246
rect 22092 34244 22116 34246
rect 22172 34244 22196 34246
rect 22252 34244 22258 34246
rect 21950 34235 22258 34244
rect 21824 34128 21876 34134
rect 21824 34070 21876 34076
rect 21836 29646 21864 34070
rect 21950 33212 22258 33221
rect 21950 33210 21956 33212
rect 22012 33210 22036 33212
rect 22092 33210 22116 33212
rect 22172 33210 22196 33212
rect 22252 33210 22258 33212
rect 22012 33158 22014 33210
rect 22194 33158 22196 33210
rect 21950 33156 21956 33158
rect 22012 33156 22036 33158
rect 22092 33156 22116 33158
rect 22172 33156 22196 33158
rect 22252 33156 22258 33158
rect 21950 33147 22258 33156
rect 21950 32124 22258 32133
rect 21950 32122 21956 32124
rect 22012 32122 22036 32124
rect 22092 32122 22116 32124
rect 22172 32122 22196 32124
rect 22252 32122 22258 32124
rect 22012 32070 22014 32122
rect 22194 32070 22196 32122
rect 21950 32068 21956 32070
rect 22012 32068 22036 32070
rect 22092 32068 22116 32070
rect 22172 32068 22196 32070
rect 22252 32068 22258 32070
rect 21950 32059 22258 32068
rect 21950 31036 22258 31045
rect 21950 31034 21956 31036
rect 22012 31034 22036 31036
rect 22092 31034 22116 31036
rect 22172 31034 22196 31036
rect 22252 31034 22258 31036
rect 22012 30982 22014 31034
rect 22194 30982 22196 31034
rect 21950 30980 21956 30982
rect 22012 30980 22036 30982
rect 22092 30980 22116 30982
rect 22172 30980 22196 30982
rect 22252 30980 22258 30982
rect 21950 30971 22258 30980
rect 21950 29948 22258 29957
rect 21950 29946 21956 29948
rect 22012 29946 22036 29948
rect 22092 29946 22116 29948
rect 22172 29946 22196 29948
rect 22252 29946 22258 29948
rect 22012 29894 22014 29946
rect 22194 29894 22196 29946
rect 21950 29892 21956 29894
rect 22012 29892 22036 29894
rect 22092 29892 22116 29894
rect 22172 29892 22196 29894
rect 22252 29892 22258 29894
rect 21950 29883 22258 29892
rect 21824 29640 21876 29646
rect 21824 29582 21876 29588
rect 21950 28860 22258 28869
rect 21950 28858 21956 28860
rect 22012 28858 22036 28860
rect 22092 28858 22116 28860
rect 22172 28858 22196 28860
rect 22252 28858 22258 28860
rect 22012 28806 22014 28858
rect 22194 28806 22196 28858
rect 21950 28804 21956 28806
rect 22012 28804 22036 28806
rect 22092 28804 22116 28806
rect 22172 28804 22196 28806
rect 22252 28804 22258 28806
rect 21950 28795 22258 28804
rect 21950 27772 22258 27781
rect 21950 27770 21956 27772
rect 22012 27770 22036 27772
rect 22092 27770 22116 27772
rect 22172 27770 22196 27772
rect 22252 27770 22258 27772
rect 22012 27718 22014 27770
rect 22194 27718 22196 27770
rect 21950 27716 21956 27718
rect 22012 27716 22036 27718
rect 22092 27716 22116 27718
rect 22172 27716 22196 27718
rect 22252 27716 22258 27718
rect 21950 27707 22258 27716
rect 21950 26684 22258 26693
rect 21950 26682 21956 26684
rect 22012 26682 22036 26684
rect 22092 26682 22116 26684
rect 22172 26682 22196 26684
rect 22252 26682 22258 26684
rect 22012 26630 22014 26682
rect 22194 26630 22196 26682
rect 21950 26628 21956 26630
rect 22012 26628 22036 26630
rect 22092 26628 22116 26630
rect 22172 26628 22196 26630
rect 22252 26628 22258 26630
rect 21950 26619 22258 26628
rect 21950 25596 22258 25605
rect 21950 25594 21956 25596
rect 22012 25594 22036 25596
rect 22092 25594 22116 25596
rect 22172 25594 22196 25596
rect 22252 25594 22258 25596
rect 22012 25542 22014 25594
rect 22194 25542 22196 25594
rect 21950 25540 21956 25542
rect 22012 25540 22036 25542
rect 22092 25540 22116 25542
rect 22172 25540 22196 25542
rect 22252 25540 22258 25542
rect 21950 25531 22258 25540
rect 21950 24508 22258 24517
rect 21950 24506 21956 24508
rect 22012 24506 22036 24508
rect 22092 24506 22116 24508
rect 22172 24506 22196 24508
rect 22252 24506 22258 24508
rect 22012 24454 22014 24506
rect 22194 24454 22196 24506
rect 21950 24452 21956 24454
rect 22012 24452 22036 24454
rect 22092 24452 22116 24454
rect 22172 24452 22196 24454
rect 22252 24452 22258 24454
rect 21950 24443 22258 24452
rect 21950 23420 22258 23429
rect 21950 23418 21956 23420
rect 22012 23418 22036 23420
rect 22092 23418 22116 23420
rect 22172 23418 22196 23420
rect 22252 23418 22258 23420
rect 22012 23366 22014 23418
rect 22194 23366 22196 23418
rect 21950 23364 21956 23366
rect 22012 23364 22036 23366
rect 22092 23364 22116 23366
rect 22172 23364 22196 23366
rect 22252 23364 22258 23366
rect 21950 23355 22258 23364
rect 21732 23316 21784 23322
rect 21732 23258 21784 23264
rect 21950 22332 22258 22341
rect 21950 22330 21956 22332
rect 22012 22330 22036 22332
rect 22092 22330 22116 22332
rect 22172 22330 22196 22332
rect 22252 22330 22258 22332
rect 22012 22278 22014 22330
rect 22194 22278 22196 22330
rect 21950 22276 21956 22278
rect 22012 22276 22036 22278
rect 22092 22276 22116 22278
rect 22172 22276 22196 22278
rect 22252 22276 22258 22278
rect 21950 22267 22258 22276
rect 21950 21244 22258 21253
rect 21950 21242 21956 21244
rect 22012 21242 22036 21244
rect 22092 21242 22116 21244
rect 22172 21242 22196 21244
rect 22252 21242 22258 21244
rect 22012 21190 22014 21242
rect 22194 21190 22196 21242
rect 21950 21188 21956 21190
rect 22012 21188 22036 21190
rect 22092 21188 22116 21190
rect 22172 21188 22196 21190
rect 22252 21188 22258 21190
rect 21950 21179 22258 21188
rect 22296 21010 22324 42078
rect 22480 41414 22508 42622
rect 22756 42566 22784 42706
rect 22744 42560 22796 42566
rect 22744 42502 22796 42508
rect 22610 42460 22918 42469
rect 22610 42458 22616 42460
rect 22672 42458 22696 42460
rect 22752 42458 22776 42460
rect 22832 42458 22856 42460
rect 22912 42458 22918 42460
rect 22672 42406 22674 42458
rect 22854 42406 22856 42458
rect 22610 42404 22616 42406
rect 22672 42404 22696 42406
rect 22752 42404 22776 42406
rect 22832 42404 22856 42406
rect 22912 42404 22918 42406
rect 22610 42395 22918 42404
rect 22388 41386 22508 41414
rect 22388 33590 22416 41386
rect 22610 41372 22918 41381
rect 22610 41370 22616 41372
rect 22672 41370 22696 41372
rect 22752 41370 22776 41372
rect 22832 41370 22856 41372
rect 22912 41370 22918 41372
rect 22672 41318 22674 41370
rect 22854 41318 22856 41370
rect 22610 41316 22616 41318
rect 22672 41316 22696 41318
rect 22752 41316 22776 41318
rect 22832 41316 22856 41318
rect 22912 41316 22918 41318
rect 22610 41307 22918 41316
rect 22836 41132 22888 41138
rect 22836 41074 22888 41080
rect 22744 40996 22796 41002
rect 22744 40938 22796 40944
rect 22468 40520 22520 40526
rect 22468 40462 22520 40468
rect 22376 33584 22428 33590
rect 22376 33526 22428 33532
rect 22480 30002 22508 40462
rect 22756 40390 22784 40938
rect 22848 40474 22876 41074
rect 23032 40730 23060 46106
rect 23124 41478 23152 49710
rect 23216 46442 23244 50662
rect 23204 46436 23256 46442
rect 23204 46378 23256 46384
rect 23204 45552 23256 45558
rect 23204 45494 23256 45500
rect 23216 42906 23244 45494
rect 23204 42900 23256 42906
rect 23204 42842 23256 42848
rect 23204 42628 23256 42634
rect 23204 42570 23256 42576
rect 23112 41472 23164 41478
rect 23112 41414 23164 41420
rect 23112 40928 23164 40934
rect 23112 40870 23164 40876
rect 23020 40724 23072 40730
rect 23020 40666 23072 40672
rect 23124 40526 23152 40870
rect 23112 40520 23164 40526
rect 22848 40446 23060 40474
rect 23112 40462 23164 40468
rect 22744 40384 22796 40390
rect 22744 40326 22796 40332
rect 22610 40284 22918 40293
rect 22610 40282 22616 40284
rect 22672 40282 22696 40284
rect 22752 40282 22776 40284
rect 22832 40282 22856 40284
rect 22912 40282 22918 40284
rect 22672 40230 22674 40282
rect 22854 40230 22856 40282
rect 22610 40228 22616 40230
rect 22672 40228 22696 40230
rect 22752 40228 22776 40230
rect 22832 40228 22856 40230
rect 22912 40228 22918 40230
rect 22610 40219 22918 40228
rect 23032 39386 23060 40446
rect 23216 39438 23244 42570
rect 23308 39438 23336 67186
rect 23388 66156 23440 66162
rect 23388 66098 23440 66104
rect 23400 62150 23428 66098
rect 23388 62144 23440 62150
rect 23388 62086 23440 62092
rect 23860 60178 23888 68342
rect 26950 68028 27258 68037
rect 26950 68026 26956 68028
rect 27012 68026 27036 68028
rect 27092 68026 27116 68028
rect 27172 68026 27196 68028
rect 27252 68026 27258 68028
rect 27012 67974 27014 68026
rect 27194 67974 27196 68026
rect 26950 67972 26956 67974
rect 27012 67972 27036 67974
rect 27092 67972 27116 67974
rect 27172 67972 27196 67974
rect 27252 67972 27258 67974
rect 26950 67963 27258 67972
rect 26148 67788 26200 67794
rect 26148 67730 26200 67736
rect 24124 67244 24176 67250
rect 24124 67186 24176 67192
rect 23848 60172 23900 60178
rect 23848 60114 23900 60120
rect 23388 59016 23440 59022
rect 23388 58958 23440 58964
rect 23400 46170 23428 58958
rect 23664 58948 23716 58954
rect 23664 58890 23716 58896
rect 23676 57322 23704 58890
rect 23664 57316 23716 57322
rect 23664 57258 23716 57264
rect 23480 52624 23532 52630
rect 23480 52566 23532 52572
rect 23492 50454 23520 52566
rect 23480 50448 23532 50454
rect 23480 50390 23532 50396
rect 23664 49836 23716 49842
rect 23664 49778 23716 49784
rect 23756 49836 23808 49842
rect 23756 49778 23808 49784
rect 23572 49768 23624 49774
rect 23572 49710 23624 49716
rect 23480 49360 23532 49366
rect 23480 49302 23532 49308
rect 23388 46164 23440 46170
rect 23388 46106 23440 46112
rect 23492 46050 23520 49302
rect 23400 46022 23520 46050
rect 23400 42702 23428 46022
rect 23388 42696 23440 42702
rect 23388 42638 23440 42644
rect 23388 42560 23440 42566
rect 23388 42502 23440 42508
rect 23400 41138 23428 42502
rect 23584 42226 23612 49710
rect 23676 42226 23704 49778
rect 23768 45558 23796 49778
rect 23756 45552 23808 45558
rect 23756 45494 23808 45500
rect 23572 42220 23624 42226
rect 23572 42162 23624 42168
rect 23664 42220 23716 42226
rect 23664 42162 23716 42168
rect 23388 41132 23440 41138
rect 23388 41074 23440 41080
rect 23676 41002 23704 42162
rect 23756 41472 23808 41478
rect 23756 41414 23808 41420
rect 23664 40996 23716 41002
rect 23664 40938 23716 40944
rect 23768 40882 23796 41414
rect 23400 40854 23796 40882
rect 23400 39846 23428 40854
rect 23570 40624 23626 40633
rect 23570 40559 23626 40568
rect 23584 40526 23612 40559
rect 23572 40520 23624 40526
rect 23572 40462 23624 40468
rect 23388 39840 23440 39846
rect 23388 39782 23440 39788
rect 23664 39840 23716 39846
rect 23664 39782 23716 39788
rect 23400 39574 23428 39782
rect 23572 39636 23624 39642
rect 23572 39578 23624 39584
rect 23388 39568 23440 39574
rect 23388 39510 23440 39516
rect 23584 39438 23612 39578
rect 23676 39438 23704 39782
rect 23204 39432 23256 39438
rect 23032 39358 23152 39386
rect 23204 39374 23256 39380
rect 23296 39432 23348 39438
rect 23296 39374 23348 39380
rect 23572 39432 23624 39438
rect 23572 39374 23624 39380
rect 23664 39432 23716 39438
rect 23860 39409 23888 60114
rect 24136 55690 24164 67186
rect 26160 66638 26188 67730
rect 27610 67484 27918 67493
rect 27610 67482 27616 67484
rect 27672 67482 27696 67484
rect 27752 67482 27776 67484
rect 27832 67482 27856 67484
rect 27912 67482 27918 67484
rect 27672 67430 27674 67482
rect 27854 67430 27856 67482
rect 27610 67428 27616 67430
rect 27672 67428 27696 67430
rect 27752 67428 27776 67430
rect 27832 67428 27856 67430
rect 27912 67428 27918 67430
rect 27610 67419 27918 67428
rect 26950 66940 27258 66949
rect 26950 66938 26956 66940
rect 27012 66938 27036 66940
rect 27092 66938 27116 66940
rect 27172 66938 27196 66940
rect 27252 66938 27258 66940
rect 27012 66886 27014 66938
rect 27194 66886 27196 66938
rect 26950 66884 26956 66886
rect 27012 66884 27036 66886
rect 27092 66884 27116 66886
rect 27172 66884 27196 66886
rect 27252 66884 27258 66886
rect 26950 66875 27258 66884
rect 26148 66632 26200 66638
rect 26148 66574 26200 66580
rect 26332 66632 26384 66638
rect 26332 66574 26384 66580
rect 26424 66632 26476 66638
rect 26424 66574 26476 66580
rect 24676 65952 24728 65958
rect 24676 65894 24728 65900
rect 24400 64320 24452 64326
rect 24400 64262 24452 64268
rect 24216 56228 24268 56234
rect 24216 56170 24268 56176
rect 24124 55684 24176 55690
rect 24124 55626 24176 55632
rect 24124 48748 24176 48754
rect 24124 48690 24176 48696
rect 23940 42764 23992 42770
rect 23940 42706 23992 42712
rect 23952 42090 23980 42706
rect 24032 42220 24084 42226
rect 24032 42162 24084 42168
rect 23940 42084 23992 42090
rect 23940 42026 23992 42032
rect 23664 39374 23716 39380
rect 23846 39400 23902 39409
rect 23020 39296 23072 39302
rect 23020 39238 23072 39244
rect 22610 39196 22918 39205
rect 22610 39194 22616 39196
rect 22672 39194 22696 39196
rect 22752 39194 22776 39196
rect 22832 39194 22856 39196
rect 22912 39194 22918 39196
rect 22672 39142 22674 39194
rect 22854 39142 22856 39194
rect 22610 39140 22616 39142
rect 22672 39140 22696 39142
rect 22752 39140 22776 39142
rect 22832 39140 22856 39142
rect 22912 39140 22918 39142
rect 22610 39131 22918 39140
rect 22610 38108 22918 38117
rect 22610 38106 22616 38108
rect 22672 38106 22696 38108
rect 22752 38106 22776 38108
rect 22832 38106 22856 38108
rect 22912 38106 22918 38108
rect 22672 38054 22674 38106
rect 22854 38054 22856 38106
rect 22610 38052 22616 38054
rect 22672 38052 22696 38054
rect 22752 38052 22776 38054
rect 22832 38052 22856 38054
rect 22912 38052 22918 38054
rect 22610 38043 22918 38052
rect 22610 37020 22918 37029
rect 22610 37018 22616 37020
rect 22672 37018 22696 37020
rect 22752 37018 22776 37020
rect 22832 37018 22856 37020
rect 22912 37018 22918 37020
rect 22672 36966 22674 37018
rect 22854 36966 22856 37018
rect 22610 36964 22616 36966
rect 22672 36964 22696 36966
rect 22752 36964 22776 36966
rect 22832 36964 22856 36966
rect 22912 36964 22918 36966
rect 22610 36955 22918 36964
rect 22610 35932 22918 35941
rect 22610 35930 22616 35932
rect 22672 35930 22696 35932
rect 22752 35930 22776 35932
rect 22832 35930 22856 35932
rect 22912 35930 22918 35932
rect 22672 35878 22674 35930
rect 22854 35878 22856 35930
rect 22610 35876 22616 35878
rect 22672 35876 22696 35878
rect 22752 35876 22776 35878
rect 22832 35876 22856 35878
rect 22912 35876 22918 35878
rect 22610 35867 22918 35876
rect 22610 34844 22918 34853
rect 22610 34842 22616 34844
rect 22672 34842 22696 34844
rect 22752 34842 22776 34844
rect 22832 34842 22856 34844
rect 22912 34842 22918 34844
rect 22672 34790 22674 34842
rect 22854 34790 22856 34842
rect 22610 34788 22616 34790
rect 22672 34788 22696 34790
rect 22752 34788 22776 34790
rect 22832 34788 22856 34790
rect 22912 34788 22918 34790
rect 22610 34779 22918 34788
rect 22610 33756 22918 33765
rect 22610 33754 22616 33756
rect 22672 33754 22696 33756
rect 22752 33754 22776 33756
rect 22832 33754 22856 33756
rect 22912 33754 22918 33756
rect 22672 33702 22674 33754
rect 22854 33702 22856 33754
rect 22610 33700 22616 33702
rect 22672 33700 22696 33702
rect 22752 33700 22776 33702
rect 22832 33700 22856 33702
rect 22912 33700 22918 33702
rect 22610 33691 22918 33700
rect 22610 32668 22918 32677
rect 22610 32666 22616 32668
rect 22672 32666 22696 32668
rect 22752 32666 22776 32668
rect 22832 32666 22856 32668
rect 22912 32666 22918 32668
rect 22672 32614 22674 32666
rect 22854 32614 22856 32666
rect 22610 32612 22616 32614
rect 22672 32612 22696 32614
rect 22752 32612 22776 32614
rect 22832 32612 22856 32614
rect 22912 32612 22918 32614
rect 22610 32603 22918 32612
rect 22610 31580 22918 31589
rect 22610 31578 22616 31580
rect 22672 31578 22696 31580
rect 22752 31578 22776 31580
rect 22832 31578 22856 31580
rect 22912 31578 22918 31580
rect 22672 31526 22674 31578
rect 22854 31526 22856 31578
rect 22610 31524 22616 31526
rect 22672 31524 22696 31526
rect 22752 31524 22776 31526
rect 22832 31524 22856 31526
rect 22912 31524 22918 31526
rect 22610 31515 22918 31524
rect 22610 30492 22918 30501
rect 22610 30490 22616 30492
rect 22672 30490 22696 30492
rect 22752 30490 22776 30492
rect 22832 30490 22856 30492
rect 22912 30490 22918 30492
rect 22672 30438 22674 30490
rect 22854 30438 22856 30490
rect 22610 30436 22616 30438
rect 22672 30436 22696 30438
rect 22752 30436 22776 30438
rect 22832 30436 22856 30438
rect 22912 30436 22918 30438
rect 22610 30427 22918 30436
rect 22388 29974 22508 30002
rect 22388 27946 22416 29974
rect 22468 29708 22520 29714
rect 22468 29650 22520 29656
rect 22376 27940 22428 27946
rect 22376 27882 22428 27888
rect 22388 24682 22416 27882
rect 22376 24676 22428 24682
rect 22376 24618 22428 24624
rect 22480 21078 22508 29650
rect 22610 29404 22918 29413
rect 22610 29402 22616 29404
rect 22672 29402 22696 29404
rect 22752 29402 22776 29404
rect 22832 29402 22856 29404
rect 22912 29402 22918 29404
rect 22672 29350 22674 29402
rect 22854 29350 22856 29402
rect 22610 29348 22616 29350
rect 22672 29348 22696 29350
rect 22752 29348 22776 29350
rect 22832 29348 22856 29350
rect 22912 29348 22918 29350
rect 22610 29339 22918 29348
rect 22610 28316 22918 28325
rect 22610 28314 22616 28316
rect 22672 28314 22696 28316
rect 22752 28314 22776 28316
rect 22832 28314 22856 28316
rect 22912 28314 22918 28316
rect 22672 28262 22674 28314
rect 22854 28262 22856 28314
rect 22610 28260 22616 28262
rect 22672 28260 22696 28262
rect 22752 28260 22776 28262
rect 22832 28260 22856 28262
rect 22912 28260 22918 28262
rect 22610 28251 22918 28260
rect 22610 27228 22918 27237
rect 22610 27226 22616 27228
rect 22672 27226 22696 27228
rect 22752 27226 22776 27228
rect 22832 27226 22856 27228
rect 22912 27226 22918 27228
rect 22672 27174 22674 27226
rect 22854 27174 22856 27226
rect 22610 27172 22616 27174
rect 22672 27172 22696 27174
rect 22752 27172 22776 27174
rect 22832 27172 22856 27174
rect 22912 27172 22918 27174
rect 22610 27163 22918 27172
rect 22610 26140 22918 26149
rect 22610 26138 22616 26140
rect 22672 26138 22696 26140
rect 22752 26138 22776 26140
rect 22832 26138 22856 26140
rect 22912 26138 22918 26140
rect 22672 26086 22674 26138
rect 22854 26086 22856 26138
rect 22610 26084 22616 26086
rect 22672 26084 22696 26086
rect 22752 26084 22776 26086
rect 22832 26084 22856 26086
rect 22912 26084 22918 26086
rect 22610 26075 22918 26084
rect 22610 25052 22918 25061
rect 22610 25050 22616 25052
rect 22672 25050 22696 25052
rect 22752 25050 22776 25052
rect 22832 25050 22856 25052
rect 22912 25050 22918 25052
rect 22672 24998 22674 25050
rect 22854 24998 22856 25050
rect 22610 24996 22616 24998
rect 22672 24996 22696 24998
rect 22752 24996 22776 24998
rect 22832 24996 22856 24998
rect 22912 24996 22918 24998
rect 22610 24987 22918 24996
rect 22610 23964 22918 23973
rect 22610 23962 22616 23964
rect 22672 23962 22696 23964
rect 22752 23962 22776 23964
rect 22832 23962 22856 23964
rect 22912 23962 22918 23964
rect 22672 23910 22674 23962
rect 22854 23910 22856 23962
rect 22610 23908 22616 23910
rect 22672 23908 22696 23910
rect 22752 23908 22776 23910
rect 22832 23908 22856 23910
rect 22912 23908 22918 23910
rect 22610 23899 22918 23908
rect 22610 22876 22918 22885
rect 22610 22874 22616 22876
rect 22672 22874 22696 22876
rect 22752 22874 22776 22876
rect 22832 22874 22856 22876
rect 22912 22874 22918 22876
rect 22672 22822 22674 22874
rect 22854 22822 22856 22874
rect 22610 22820 22616 22822
rect 22672 22820 22696 22822
rect 22752 22820 22776 22822
rect 22832 22820 22856 22822
rect 22912 22820 22918 22822
rect 22610 22811 22918 22820
rect 22610 21788 22918 21797
rect 22610 21786 22616 21788
rect 22672 21786 22696 21788
rect 22752 21786 22776 21788
rect 22832 21786 22856 21788
rect 22912 21786 22918 21788
rect 22672 21734 22674 21786
rect 22854 21734 22856 21786
rect 22610 21732 22616 21734
rect 22672 21732 22696 21734
rect 22752 21732 22776 21734
rect 22832 21732 22856 21734
rect 22912 21732 22918 21734
rect 22610 21723 22918 21732
rect 22468 21072 22520 21078
rect 22468 21014 22520 21020
rect 22284 21004 22336 21010
rect 22284 20946 22336 20952
rect 21824 20936 21876 20942
rect 21824 20878 21876 20884
rect 21836 15162 21864 20878
rect 21950 20156 22258 20165
rect 21950 20154 21956 20156
rect 22012 20154 22036 20156
rect 22092 20154 22116 20156
rect 22172 20154 22196 20156
rect 22252 20154 22258 20156
rect 22012 20102 22014 20154
rect 22194 20102 22196 20154
rect 21950 20100 21956 20102
rect 22012 20100 22036 20102
rect 22092 20100 22116 20102
rect 22172 20100 22196 20102
rect 22252 20100 22258 20102
rect 21950 20091 22258 20100
rect 22296 19174 22324 20946
rect 22376 20936 22428 20942
rect 22376 20878 22428 20884
rect 22388 20398 22416 20878
rect 22376 20392 22428 20398
rect 22376 20334 22428 20340
rect 22284 19168 22336 19174
rect 22284 19110 22336 19116
rect 21950 19068 22258 19077
rect 21950 19066 21956 19068
rect 22012 19066 22036 19068
rect 22092 19066 22116 19068
rect 22172 19066 22196 19068
rect 22252 19066 22258 19068
rect 22012 19014 22014 19066
rect 22194 19014 22196 19066
rect 21950 19012 21956 19014
rect 22012 19012 22036 19014
rect 22092 19012 22116 19014
rect 22172 19012 22196 19014
rect 22252 19012 22258 19014
rect 21950 19003 22258 19012
rect 21950 17980 22258 17989
rect 21950 17978 21956 17980
rect 22012 17978 22036 17980
rect 22092 17978 22116 17980
rect 22172 17978 22196 17980
rect 22252 17978 22258 17980
rect 22012 17926 22014 17978
rect 22194 17926 22196 17978
rect 21950 17924 21956 17926
rect 22012 17924 22036 17926
rect 22092 17924 22116 17926
rect 22172 17924 22196 17926
rect 22252 17924 22258 17926
rect 21950 17915 22258 17924
rect 21950 16892 22258 16901
rect 21950 16890 21956 16892
rect 22012 16890 22036 16892
rect 22092 16890 22116 16892
rect 22172 16890 22196 16892
rect 22252 16890 22258 16892
rect 22012 16838 22014 16890
rect 22194 16838 22196 16890
rect 21950 16836 21956 16838
rect 22012 16836 22036 16838
rect 22092 16836 22116 16838
rect 22172 16836 22196 16838
rect 22252 16836 22258 16838
rect 21950 16827 22258 16836
rect 22296 16794 22324 19110
rect 22284 16788 22336 16794
rect 22284 16730 22336 16736
rect 22388 16726 22416 20334
rect 22376 16720 22428 16726
rect 22376 16662 22428 16668
rect 21950 15804 22258 15813
rect 21950 15802 21956 15804
rect 22012 15802 22036 15804
rect 22092 15802 22116 15804
rect 22172 15802 22196 15804
rect 22252 15802 22258 15804
rect 22012 15750 22014 15802
rect 22194 15750 22196 15802
rect 21950 15748 21956 15750
rect 22012 15748 22036 15750
rect 22092 15748 22116 15750
rect 22172 15748 22196 15750
rect 22252 15748 22258 15750
rect 21950 15739 22258 15748
rect 21824 15156 21876 15162
rect 21824 15098 21876 15104
rect 21640 13184 21692 13190
rect 21640 13126 21692 13132
rect 21836 12434 21864 15098
rect 22374 15056 22430 15065
rect 22374 14991 22430 15000
rect 21950 14716 22258 14725
rect 21950 14714 21956 14716
rect 22012 14714 22036 14716
rect 22092 14714 22116 14716
rect 22172 14714 22196 14716
rect 22252 14714 22258 14716
rect 22012 14662 22014 14714
rect 22194 14662 22196 14714
rect 21950 14660 21956 14662
rect 22012 14660 22036 14662
rect 22092 14660 22116 14662
rect 22172 14660 22196 14662
rect 22252 14660 22258 14662
rect 21950 14651 22258 14660
rect 21950 13628 22258 13637
rect 21950 13626 21956 13628
rect 22012 13626 22036 13628
rect 22092 13626 22116 13628
rect 22172 13626 22196 13628
rect 22252 13626 22258 13628
rect 22012 13574 22014 13626
rect 22194 13574 22196 13626
rect 21950 13572 21956 13574
rect 22012 13572 22036 13574
rect 22092 13572 22116 13574
rect 22172 13572 22196 13574
rect 22252 13572 22258 13574
rect 21950 13563 22258 13572
rect 21950 12540 22258 12549
rect 21950 12538 21956 12540
rect 22012 12538 22036 12540
rect 22092 12538 22116 12540
rect 22172 12538 22196 12540
rect 22252 12538 22258 12540
rect 22012 12486 22014 12538
rect 22194 12486 22196 12538
rect 21950 12484 21956 12486
rect 22012 12484 22036 12486
rect 22092 12484 22116 12486
rect 22172 12484 22196 12486
rect 22252 12484 22258 12486
rect 21950 12475 22258 12484
rect 21744 12406 21864 12434
rect 21548 12300 21600 12306
rect 21548 12242 21600 12248
rect 21364 12232 21416 12238
rect 21364 12174 21416 12180
rect 21180 11008 21232 11014
rect 21180 10950 21232 10956
rect 20444 10736 20496 10742
rect 20444 10678 20496 10684
rect 20260 8900 20312 8906
rect 20260 8842 20312 8848
rect 20076 7404 20128 7410
rect 20076 7346 20128 7352
rect 19984 4684 20036 4690
rect 19984 4626 20036 4632
rect 18236 4548 18288 4554
rect 18236 4490 18288 4496
rect 19616 4548 19668 4554
rect 19616 4490 19668 4496
rect 17610 4380 17918 4389
rect 17610 4378 17616 4380
rect 17672 4378 17696 4380
rect 17752 4378 17776 4380
rect 17832 4378 17856 4380
rect 17912 4378 17918 4380
rect 17672 4326 17674 4378
rect 17854 4326 17856 4378
rect 17610 4324 17616 4326
rect 17672 4324 17696 4326
rect 17752 4324 17776 4326
rect 17832 4324 17856 4326
rect 17912 4324 17918 4326
rect 17610 4315 17918 4324
rect 17610 3292 17918 3301
rect 17610 3290 17616 3292
rect 17672 3290 17696 3292
rect 17752 3290 17776 3292
rect 17832 3290 17856 3292
rect 17912 3290 17918 3292
rect 17672 3238 17674 3290
rect 17854 3238 17856 3290
rect 17610 3236 17616 3238
rect 17672 3236 17696 3238
rect 17752 3236 17776 3238
rect 17832 3236 17856 3238
rect 17912 3236 17918 3238
rect 17610 3227 17918 3236
rect 20088 2990 20116 7346
rect 21744 6730 21772 12406
rect 21950 11452 22258 11461
rect 21950 11450 21956 11452
rect 22012 11450 22036 11452
rect 22092 11450 22116 11452
rect 22172 11450 22196 11452
rect 22252 11450 22258 11452
rect 22012 11398 22014 11450
rect 22194 11398 22196 11450
rect 21950 11396 21956 11398
rect 22012 11396 22036 11398
rect 22092 11396 22116 11398
rect 22172 11396 22196 11398
rect 22252 11396 22258 11398
rect 21950 11387 22258 11396
rect 21950 10364 22258 10373
rect 21950 10362 21956 10364
rect 22012 10362 22036 10364
rect 22092 10362 22116 10364
rect 22172 10362 22196 10364
rect 22252 10362 22258 10364
rect 22012 10310 22014 10362
rect 22194 10310 22196 10362
rect 21950 10308 21956 10310
rect 22012 10308 22036 10310
rect 22092 10308 22116 10310
rect 22172 10308 22196 10310
rect 22252 10308 22258 10310
rect 21950 10299 22258 10308
rect 21950 9276 22258 9285
rect 21950 9274 21956 9276
rect 22012 9274 22036 9276
rect 22092 9274 22116 9276
rect 22172 9274 22196 9276
rect 22252 9274 22258 9276
rect 22012 9222 22014 9274
rect 22194 9222 22196 9274
rect 21950 9220 21956 9222
rect 22012 9220 22036 9222
rect 22092 9220 22116 9222
rect 22172 9220 22196 9222
rect 22252 9220 22258 9222
rect 21950 9211 22258 9220
rect 21950 8188 22258 8197
rect 21950 8186 21956 8188
rect 22012 8186 22036 8188
rect 22092 8186 22116 8188
rect 22172 8186 22196 8188
rect 22252 8186 22258 8188
rect 22012 8134 22014 8186
rect 22194 8134 22196 8186
rect 21950 8132 21956 8134
rect 22012 8132 22036 8134
rect 22092 8132 22116 8134
rect 22172 8132 22196 8134
rect 22252 8132 22258 8134
rect 21950 8123 22258 8132
rect 22388 7818 22416 14991
rect 22480 7954 22508 21014
rect 22610 20700 22918 20709
rect 22610 20698 22616 20700
rect 22672 20698 22696 20700
rect 22752 20698 22776 20700
rect 22832 20698 22856 20700
rect 22912 20698 22918 20700
rect 22672 20646 22674 20698
rect 22854 20646 22856 20698
rect 22610 20644 22616 20646
rect 22672 20644 22696 20646
rect 22752 20644 22776 20646
rect 22832 20644 22856 20646
rect 22912 20644 22918 20646
rect 22610 20635 22918 20644
rect 23032 20534 23060 39238
rect 23124 35222 23152 39358
rect 23216 35834 23244 39374
rect 23204 35828 23256 35834
rect 23204 35770 23256 35776
rect 23112 35216 23164 35222
rect 23112 35158 23164 35164
rect 23124 34746 23152 35158
rect 23112 34740 23164 34746
rect 23112 34682 23164 34688
rect 23308 33522 23336 39374
rect 23388 38752 23440 38758
rect 23386 38720 23388 38729
rect 23440 38720 23442 38729
rect 23386 38655 23442 38664
rect 23480 36780 23532 36786
rect 23480 36722 23532 36728
rect 23388 35828 23440 35834
rect 23388 35770 23440 35776
rect 23296 33516 23348 33522
rect 23296 33458 23348 33464
rect 23308 32450 23336 33458
rect 23124 32422 23336 32450
rect 23124 26926 23152 32422
rect 23400 31754 23428 35770
rect 23216 31726 23428 31754
rect 23216 29646 23244 31726
rect 23386 31104 23442 31113
rect 23386 31039 23442 31048
rect 23204 29640 23256 29646
rect 23204 29582 23256 29588
rect 23296 29504 23348 29510
rect 23296 29446 23348 29452
rect 23308 27606 23336 29446
rect 23296 27600 23348 27606
rect 23296 27542 23348 27548
rect 23112 26920 23164 26926
rect 23112 26862 23164 26868
rect 23296 24200 23348 24206
rect 23296 24142 23348 24148
rect 23020 20528 23072 20534
rect 23020 20470 23072 20476
rect 23308 20398 23336 24142
rect 23296 20392 23348 20398
rect 23296 20334 23348 20340
rect 23296 20256 23348 20262
rect 23296 20198 23348 20204
rect 22610 19612 22918 19621
rect 22610 19610 22616 19612
rect 22672 19610 22696 19612
rect 22752 19610 22776 19612
rect 22832 19610 22856 19612
rect 22912 19610 22918 19612
rect 22672 19558 22674 19610
rect 22854 19558 22856 19610
rect 22610 19556 22616 19558
rect 22672 19556 22696 19558
rect 22752 19556 22776 19558
rect 22832 19556 22856 19558
rect 22912 19556 22918 19558
rect 22610 19547 22918 19556
rect 22610 18524 22918 18533
rect 22610 18522 22616 18524
rect 22672 18522 22696 18524
rect 22752 18522 22776 18524
rect 22832 18522 22856 18524
rect 22912 18522 22918 18524
rect 22672 18470 22674 18522
rect 22854 18470 22856 18522
rect 22610 18468 22616 18470
rect 22672 18468 22696 18470
rect 22752 18468 22776 18470
rect 22832 18468 22856 18470
rect 22912 18468 22918 18470
rect 22610 18459 22918 18468
rect 22610 17436 22918 17445
rect 22610 17434 22616 17436
rect 22672 17434 22696 17436
rect 22752 17434 22776 17436
rect 22832 17434 22856 17436
rect 22912 17434 22918 17436
rect 22672 17382 22674 17434
rect 22854 17382 22856 17434
rect 22610 17380 22616 17382
rect 22672 17380 22696 17382
rect 22752 17380 22776 17382
rect 22832 17380 22856 17382
rect 22912 17380 22918 17382
rect 22610 17371 22918 17380
rect 22610 16348 22918 16357
rect 22610 16346 22616 16348
rect 22672 16346 22696 16348
rect 22752 16346 22776 16348
rect 22832 16346 22856 16348
rect 22912 16346 22918 16348
rect 22672 16294 22674 16346
rect 22854 16294 22856 16346
rect 22610 16292 22616 16294
rect 22672 16292 22696 16294
rect 22752 16292 22776 16294
rect 22832 16292 22856 16294
rect 22912 16292 22918 16294
rect 22610 16283 22918 16292
rect 22610 15260 22918 15269
rect 22610 15258 22616 15260
rect 22672 15258 22696 15260
rect 22752 15258 22776 15260
rect 22832 15258 22856 15260
rect 22912 15258 22918 15260
rect 22672 15206 22674 15258
rect 22854 15206 22856 15258
rect 22610 15204 22616 15206
rect 22672 15204 22696 15206
rect 22752 15204 22776 15206
rect 22832 15204 22856 15206
rect 22912 15204 22918 15206
rect 22610 15195 22918 15204
rect 22610 14172 22918 14181
rect 22610 14170 22616 14172
rect 22672 14170 22696 14172
rect 22752 14170 22776 14172
rect 22832 14170 22856 14172
rect 22912 14170 22918 14172
rect 22672 14118 22674 14170
rect 22854 14118 22856 14170
rect 22610 14116 22616 14118
rect 22672 14116 22696 14118
rect 22752 14116 22776 14118
rect 22832 14116 22856 14118
rect 22912 14116 22918 14118
rect 22610 14107 22918 14116
rect 22610 13084 22918 13093
rect 22610 13082 22616 13084
rect 22672 13082 22696 13084
rect 22752 13082 22776 13084
rect 22832 13082 22856 13084
rect 22912 13082 22918 13084
rect 22672 13030 22674 13082
rect 22854 13030 22856 13082
rect 22610 13028 22616 13030
rect 22672 13028 22696 13030
rect 22752 13028 22776 13030
rect 22832 13028 22856 13030
rect 22912 13028 22918 13030
rect 22610 13019 22918 13028
rect 23308 12986 23336 20198
rect 23296 12980 23348 12986
rect 23296 12922 23348 12928
rect 23400 12850 23428 31039
rect 23492 16574 23520 36722
rect 23584 33930 23612 39374
rect 23846 39335 23902 39344
rect 23756 39296 23808 39302
rect 23756 39238 23808 39244
rect 23768 36689 23796 39238
rect 23860 38894 23888 39335
rect 23848 38888 23900 38894
rect 23848 38830 23900 38836
rect 23848 38412 23900 38418
rect 23848 38354 23900 38360
rect 23754 36680 23810 36689
rect 23754 36615 23810 36624
rect 23572 33924 23624 33930
rect 23572 33866 23624 33872
rect 23860 31754 23888 38354
rect 23952 36786 23980 42026
rect 23940 36780 23992 36786
rect 23940 36722 23992 36728
rect 23860 31726 23980 31754
rect 23572 29844 23624 29850
rect 23572 29786 23624 29792
rect 23584 29306 23612 29786
rect 23572 29300 23624 29306
rect 23572 29242 23624 29248
rect 23952 28762 23980 31726
rect 23940 28756 23992 28762
rect 23940 28698 23992 28704
rect 24044 21010 24072 42162
rect 24136 38554 24164 48690
rect 24124 38548 24176 38554
rect 24124 38490 24176 38496
rect 24124 33924 24176 33930
rect 24124 33866 24176 33872
rect 24032 21004 24084 21010
rect 24032 20946 24084 20952
rect 24136 20466 24164 33866
rect 24228 33590 24256 56170
rect 24308 49836 24360 49842
rect 24308 49778 24360 49784
rect 24320 42226 24348 49778
rect 24412 49230 24440 64262
rect 24688 49842 24716 65894
rect 25504 65680 25556 65686
rect 25504 65622 25556 65628
rect 25596 65680 25648 65686
rect 25596 65622 25648 65628
rect 25044 62756 25096 62762
rect 25044 62698 25096 62704
rect 24860 57588 24912 57594
rect 24860 57530 24912 57536
rect 24872 54738 24900 57530
rect 24860 54732 24912 54738
rect 24860 54674 24912 54680
rect 24676 49836 24728 49842
rect 24676 49778 24728 49784
rect 24400 49224 24452 49230
rect 24400 49166 24452 49172
rect 24492 45280 24544 45286
rect 24492 45222 24544 45228
rect 24308 42220 24360 42226
rect 24308 42162 24360 42168
rect 24400 40452 24452 40458
rect 24400 40394 24452 40400
rect 24308 38888 24360 38894
rect 24306 38856 24308 38865
rect 24360 38856 24362 38865
rect 24306 38791 24362 38800
rect 24216 33584 24268 33590
rect 24216 33526 24268 33532
rect 24308 32360 24360 32366
rect 24308 32302 24360 32308
rect 24216 27600 24268 27606
rect 24216 27542 24268 27548
rect 24124 20460 24176 20466
rect 24124 20402 24176 20408
rect 24228 17746 24256 27542
rect 24320 25770 24348 32302
rect 24412 28626 24440 40394
rect 24504 33114 24532 45222
rect 24688 42294 24716 49778
rect 25056 49774 25084 62698
rect 25044 49768 25096 49774
rect 25044 49710 25096 49716
rect 24860 49088 24912 49094
rect 24860 49030 24912 49036
rect 24872 48346 24900 49030
rect 24860 48340 24912 48346
rect 24860 48282 24912 48288
rect 24676 42288 24728 42294
rect 24676 42230 24728 42236
rect 24676 40520 24728 40526
rect 24676 40462 24728 40468
rect 24582 38992 24638 39001
rect 24582 38927 24638 38936
rect 24596 38826 24624 38927
rect 24584 38820 24636 38826
rect 24584 38762 24636 38768
rect 24584 38344 24636 38350
rect 24584 38286 24636 38292
rect 24492 33108 24544 33114
rect 24492 33050 24544 33056
rect 24596 31890 24624 38286
rect 24584 31884 24636 31890
rect 24584 31826 24636 31832
rect 24584 31272 24636 31278
rect 24584 31214 24636 31220
rect 24492 29300 24544 29306
rect 24492 29242 24544 29248
rect 24400 28620 24452 28626
rect 24400 28562 24452 28568
rect 24412 28082 24440 28562
rect 24400 28076 24452 28082
rect 24400 28018 24452 28024
rect 24308 25764 24360 25770
rect 24308 25706 24360 25712
rect 24216 17740 24268 17746
rect 24216 17682 24268 17688
rect 24504 16658 24532 29242
rect 24596 23730 24624 31214
rect 24688 28082 24716 40462
rect 24860 40112 24912 40118
rect 24860 40054 24912 40060
rect 24766 38448 24822 38457
rect 24766 38383 24768 38392
rect 24820 38383 24822 38392
rect 24768 38354 24820 38360
rect 24872 34218 24900 40054
rect 24952 35692 25004 35698
rect 24952 35634 25004 35640
rect 24964 35494 24992 35634
rect 24952 35488 25004 35494
rect 24952 35430 25004 35436
rect 24872 34190 24992 34218
rect 24860 34060 24912 34066
rect 24860 34002 24912 34008
rect 24872 33590 24900 34002
rect 24860 33584 24912 33590
rect 24860 33526 24912 33532
rect 24964 31754 24992 34190
rect 24872 31726 24992 31754
rect 24768 31272 24820 31278
rect 24768 31214 24820 31220
rect 24780 30938 24808 31214
rect 24768 30932 24820 30938
rect 24768 30874 24820 30880
rect 24872 28218 24900 31726
rect 24952 31204 25004 31210
rect 24952 31146 25004 31152
rect 24860 28212 24912 28218
rect 24860 28154 24912 28160
rect 24676 28076 24728 28082
rect 24676 28018 24728 28024
rect 24688 24410 24716 28018
rect 24964 26518 24992 31146
rect 24952 26512 25004 26518
rect 24952 26454 25004 26460
rect 24950 26344 25006 26353
rect 24950 26279 25006 26288
rect 24676 24404 24728 24410
rect 24676 24346 24728 24352
rect 24584 23724 24636 23730
rect 24584 23666 24636 23672
rect 24964 20602 24992 26279
rect 25056 22098 25084 49710
rect 25136 41132 25188 41138
rect 25136 41074 25188 41080
rect 25148 40526 25176 41074
rect 25136 40520 25188 40526
rect 25136 40462 25188 40468
rect 25226 38040 25282 38049
rect 25226 37975 25282 37984
rect 25240 37942 25268 37975
rect 25516 37942 25544 65622
rect 25608 50182 25636 65622
rect 25688 58948 25740 58954
rect 25688 58890 25740 58896
rect 25700 52086 25728 58890
rect 26160 57798 26188 66574
rect 26344 65754 26372 66574
rect 26436 66026 26464 66574
rect 27610 66396 27918 66405
rect 27610 66394 27616 66396
rect 27672 66394 27696 66396
rect 27752 66394 27776 66396
rect 27832 66394 27856 66396
rect 27912 66394 27918 66396
rect 27672 66342 27674 66394
rect 27854 66342 27856 66394
rect 27610 66340 27616 66342
rect 27672 66340 27696 66342
rect 27752 66340 27776 66342
rect 27832 66340 27856 66342
rect 27912 66340 27918 66342
rect 27610 66331 27918 66340
rect 26424 66020 26476 66026
rect 26424 65962 26476 65968
rect 26950 65852 27258 65861
rect 26950 65850 26956 65852
rect 27012 65850 27036 65852
rect 27092 65850 27116 65852
rect 27172 65850 27196 65852
rect 27252 65850 27258 65852
rect 27012 65798 27014 65850
rect 27194 65798 27196 65850
rect 26950 65796 26956 65798
rect 27012 65796 27036 65798
rect 27092 65796 27116 65798
rect 27172 65796 27196 65798
rect 27252 65796 27258 65798
rect 26950 65787 27258 65796
rect 26332 65748 26384 65754
rect 26332 65690 26384 65696
rect 27610 65308 27918 65317
rect 27610 65306 27616 65308
rect 27672 65306 27696 65308
rect 27752 65306 27776 65308
rect 27832 65306 27856 65308
rect 27912 65306 27918 65308
rect 27672 65254 27674 65306
rect 27854 65254 27856 65306
rect 27610 65252 27616 65254
rect 27672 65252 27696 65254
rect 27752 65252 27776 65254
rect 27832 65252 27856 65254
rect 27912 65252 27918 65254
rect 27610 65243 27918 65252
rect 26950 64764 27258 64773
rect 26950 64762 26956 64764
rect 27012 64762 27036 64764
rect 27092 64762 27116 64764
rect 27172 64762 27196 64764
rect 27252 64762 27258 64764
rect 27012 64710 27014 64762
rect 27194 64710 27196 64762
rect 26950 64708 26956 64710
rect 27012 64708 27036 64710
rect 27092 64708 27116 64710
rect 27172 64708 27196 64710
rect 27252 64708 27258 64710
rect 26950 64699 27258 64708
rect 27610 64220 27918 64229
rect 27610 64218 27616 64220
rect 27672 64218 27696 64220
rect 27752 64218 27776 64220
rect 27832 64218 27856 64220
rect 27912 64218 27918 64220
rect 27672 64166 27674 64218
rect 27854 64166 27856 64218
rect 27610 64164 27616 64166
rect 27672 64164 27696 64166
rect 27752 64164 27776 64166
rect 27832 64164 27856 64166
rect 27912 64164 27918 64166
rect 27610 64155 27918 64164
rect 26950 63676 27258 63685
rect 26950 63674 26956 63676
rect 27012 63674 27036 63676
rect 27092 63674 27116 63676
rect 27172 63674 27196 63676
rect 27252 63674 27258 63676
rect 27012 63622 27014 63674
rect 27194 63622 27196 63674
rect 26950 63620 26956 63622
rect 27012 63620 27036 63622
rect 27092 63620 27116 63622
rect 27172 63620 27196 63622
rect 27252 63620 27258 63622
rect 26950 63611 27258 63620
rect 26700 63300 26752 63306
rect 26700 63242 26752 63248
rect 26712 59226 26740 63242
rect 27988 63232 28040 63238
rect 27988 63174 28040 63180
rect 27610 63132 27918 63141
rect 27610 63130 27616 63132
rect 27672 63130 27696 63132
rect 27752 63130 27776 63132
rect 27832 63130 27856 63132
rect 27912 63130 27918 63132
rect 27672 63078 27674 63130
rect 27854 63078 27856 63130
rect 27610 63076 27616 63078
rect 27672 63076 27696 63078
rect 27752 63076 27776 63078
rect 27832 63076 27856 63078
rect 27912 63076 27918 63078
rect 27610 63067 27918 63076
rect 26950 62588 27258 62597
rect 26950 62586 26956 62588
rect 27012 62586 27036 62588
rect 27092 62586 27116 62588
rect 27172 62586 27196 62588
rect 27252 62586 27258 62588
rect 27012 62534 27014 62586
rect 27194 62534 27196 62586
rect 26950 62532 26956 62534
rect 27012 62532 27036 62534
rect 27092 62532 27116 62534
rect 27172 62532 27196 62534
rect 27252 62532 27258 62534
rect 26950 62523 27258 62532
rect 27436 62484 27488 62490
rect 27436 62426 27488 62432
rect 26950 61500 27258 61509
rect 26950 61498 26956 61500
rect 27012 61498 27036 61500
rect 27092 61498 27116 61500
rect 27172 61498 27196 61500
rect 27252 61498 27258 61500
rect 27012 61446 27014 61498
rect 27194 61446 27196 61498
rect 26950 61444 26956 61446
rect 27012 61444 27036 61446
rect 27092 61444 27116 61446
rect 27172 61444 27196 61446
rect 27252 61444 27258 61446
rect 26950 61435 27258 61444
rect 26950 60412 27258 60421
rect 26950 60410 26956 60412
rect 27012 60410 27036 60412
rect 27092 60410 27116 60412
rect 27172 60410 27196 60412
rect 27252 60410 27258 60412
rect 27012 60358 27014 60410
rect 27194 60358 27196 60410
rect 26950 60356 26956 60358
rect 27012 60356 27036 60358
rect 27092 60356 27116 60358
rect 27172 60356 27196 60358
rect 27252 60356 27258 60358
rect 26950 60347 27258 60356
rect 26950 59324 27258 59333
rect 26950 59322 26956 59324
rect 27012 59322 27036 59324
rect 27092 59322 27116 59324
rect 27172 59322 27196 59324
rect 27252 59322 27258 59324
rect 27012 59270 27014 59322
rect 27194 59270 27196 59322
rect 26950 59268 26956 59270
rect 27012 59268 27036 59270
rect 27092 59268 27116 59270
rect 27172 59268 27196 59270
rect 27252 59268 27258 59270
rect 26950 59259 27258 59268
rect 26700 59220 26752 59226
rect 26700 59162 26752 59168
rect 27448 58954 27476 62426
rect 27610 62044 27918 62053
rect 27610 62042 27616 62044
rect 27672 62042 27696 62044
rect 27752 62042 27776 62044
rect 27832 62042 27856 62044
rect 27912 62042 27918 62044
rect 27672 61990 27674 62042
rect 27854 61990 27856 62042
rect 27610 61988 27616 61990
rect 27672 61988 27696 61990
rect 27752 61988 27776 61990
rect 27832 61988 27856 61990
rect 27912 61988 27918 61990
rect 27610 61979 27918 61988
rect 27610 60956 27918 60965
rect 27610 60954 27616 60956
rect 27672 60954 27696 60956
rect 27752 60954 27776 60956
rect 27832 60954 27856 60956
rect 27912 60954 27918 60956
rect 27672 60902 27674 60954
rect 27854 60902 27856 60954
rect 27610 60900 27616 60902
rect 27672 60900 27696 60902
rect 27752 60900 27776 60902
rect 27832 60900 27856 60902
rect 27912 60900 27918 60902
rect 27610 60891 27918 60900
rect 27528 59968 27580 59974
rect 27528 59910 27580 59916
rect 27436 58948 27488 58954
rect 27436 58890 27488 58896
rect 26950 58236 27258 58245
rect 26950 58234 26956 58236
rect 27012 58234 27036 58236
rect 27092 58234 27116 58236
rect 27172 58234 27196 58236
rect 27252 58234 27258 58236
rect 27012 58182 27014 58234
rect 27194 58182 27196 58234
rect 26950 58180 26956 58182
rect 27012 58180 27036 58182
rect 27092 58180 27116 58182
rect 27172 58180 27196 58182
rect 27252 58180 27258 58182
rect 26950 58171 27258 58180
rect 26148 57792 26200 57798
rect 26148 57734 26200 57740
rect 26950 57148 27258 57157
rect 26950 57146 26956 57148
rect 27012 57146 27036 57148
rect 27092 57146 27116 57148
rect 27172 57146 27196 57148
rect 27252 57146 27258 57148
rect 27012 57094 27014 57146
rect 27194 57094 27196 57146
rect 26950 57092 26956 57094
rect 27012 57092 27036 57094
rect 27092 57092 27116 57094
rect 27172 57092 27196 57094
rect 27252 57092 27258 57094
rect 26950 57083 27258 57092
rect 26240 57044 26292 57050
rect 26240 56986 26292 56992
rect 26252 56846 26280 56986
rect 26148 56840 26200 56846
rect 26148 56782 26200 56788
rect 26240 56840 26292 56846
rect 26240 56782 26292 56788
rect 25688 52080 25740 52086
rect 25688 52022 25740 52028
rect 25596 50176 25648 50182
rect 25596 50118 25648 50124
rect 25700 48314 25728 52022
rect 26160 50862 26188 56782
rect 26950 56060 27258 56069
rect 26950 56058 26956 56060
rect 27012 56058 27036 56060
rect 27092 56058 27116 56060
rect 27172 56058 27196 56060
rect 27252 56058 27258 56060
rect 27012 56006 27014 56058
rect 27194 56006 27196 56058
rect 26950 56004 26956 56006
rect 27012 56004 27036 56006
rect 27092 56004 27116 56006
rect 27172 56004 27196 56006
rect 27252 56004 27258 56006
rect 26950 55995 27258 56004
rect 26950 54972 27258 54981
rect 26950 54970 26956 54972
rect 27012 54970 27036 54972
rect 27092 54970 27116 54972
rect 27172 54970 27196 54972
rect 27252 54970 27258 54972
rect 27012 54918 27014 54970
rect 27194 54918 27196 54970
rect 26950 54916 26956 54918
rect 27012 54916 27036 54918
rect 27092 54916 27116 54918
rect 27172 54916 27196 54918
rect 27252 54916 27258 54918
rect 26950 54907 27258 54916
rect 26950 53884 27258 53893
rect 26950 53882 26956 53884
rect 27012 53882 27036 53884
rect 27092 53882 27116 53884
rect 27172 53882 27196 53884
rect 27252 53882 27258 53884
rect 27012 53830 27014 53882
rect 27194 53830 27196 53882
rect 26950 53828 26956 53830
rect 27012 53828 27036 53830
rect 27092 53828 27116 53830
rect 27172 53828 27196 53830
rect 27252 53828 27258 53830
rect 26950 53819 27258 53828
rect 26792 53508 26844 53514
rect 26792 53450 26844 53456
rect 26148 50856 26200 50862
rect 26148 50798 26200 50804
rect 25700 48286 26096 48314
rect 25872 46980 25924 46986
rect 25872 46922 25924 46928
rect 25688 42356 25740 42362
rect 25688 42298 25740 42304
rect 25228 37936 25280 37942
rect 25228 37878 25280 37884
rect 25504 37936 25556 37942
rect 25504 37878 25556 37884
rect 25136 35556 25188 35562
rect 25136 35498 25188 35504
rect 25148 25906 25176 35498
rect 25136 25900 25188 25906
rect 25136 25842 25188 25848
rect 25044 22092 25096 22098
rect 25044 22034 25096 22040
rect 24952 20596 25004 20602
rect 24952 20538 25004 20544
rect 25148 20482 25176 25842
rect 24872 20454 25176 20482
rect 24676 20392 24728 20398
rect 24676 20334 24728 20340
rect 24584 20324 24636 20330
rect 24584 20266 24636 20272
rect 24492 16652 24544 16658
rect 24492 16594 24544 16600
rect 23492 16546 23612 16574
rect 23584 15026 23612 16546
rect 23572 15020 23624 15026
rect 23572 14962 23624 14968
rect 23480 14544 23532 14550
rect 23480 14486 23532 14492
rect 23388 12844 23440 12850
rect 23388 12786 23440 12792
rect 22610 11996 22918 12005
rect 22610 11994 22616 11996
rect 22672 11994 22696 11996
rect 22752 11994 22776 11996
rect 22832 11994 22856 11996
rect 22912 11994 22918 11996
rect 22672 11942 22674 11994
rect 22854 11942 22856 11994
rect 22610 11940 22616 11942
rect 22672 11940 22696 11942
rect 22752 11940 22776 11942
rect 22832 11940 22856 11942
rect 22912 11940 22918 11942
rect 22610 11931 22918 11940
rect 22610 10908 22918 10917
rect 22610 10906 22616 10908
rect 22672 10906 22696 10908
rect 22752 10906 22776 10908
rect 22832 10906 22856 10908
rect 22912 10906 22918 10908
rect 22672 10854 22674 10906
rect 22854 10854 22856 10906
rect 22610 10852 22616 10854
rect 22672 10852 22696 10854
rect 22752 10852 22776 10854
rect 22832 10852 22856 10854
rect 22912 10852 22918 10854
rect 22610 10843 22918 10852
rect 22610 9820 22918 9829
rect 22610 9818 22616 9820
rect 22672 9818 22696 9820
rect 22752 9818 22776 9820
rect 22832 9818 22856 9820
rect 22912 9818 22918 9820
rect 22672 9766 22674 9818
rect 22854 9766 22856 9818
rect 22610 9764 22616 9766
rect 22672 9764 22696 9766
rect 22752 9764 22776 9766
rect 22832 9764 22856 9766
rect 22912 9764 22918 9766
rect 22610 9755 22918 9764
rect 23400 9110 23428 12786
rect 23492 9518 23520 14486
rect 23584 11218 23612 14962
rect 23572 11212 23624 11218
rect 23572 11154 23624 11160
rect 23480 9512 23532 9518
rect 23480 9454 23532 9460
rect 23388 9104 23440 9110
rect 23388 9046 23440 9052
rect 22610 8732 22918 8741
rect 22610 8730 22616 8732
rect 22672 8730 22696 8732
rect 22752 8730 22776 8732
rect 22832 8730 22856 8732
rect 22912 8730 22918 8732
rect 22672 8678 22674 8730
rect 22854 8678 22856 8730
rect 22610 8676 22616 8678
rect 22672 8676 22696 8678
rect 22752 8676 22776 8678
rect 22832 8676 22856 8678
rect 22912 8676 22918 8678
rect 22610 8667 22918 8676
rect 22468 7948 22520 7954
rect 22468 7890 22520 7896
rect 22376 7812 22428 7818
rect 22376 7754 22428 7760
rect 21950 7100 22258 7109
rect 21950 7098 21956 7100
rect 22012 7098 22036 7100
rect 22092 7098 22116 7100
rect 22172 7098 22196 7100
rect 22252 7098 22258 7100
rect 22012 7046 22014 7098
rect 22194 7046 22196 7098
rect 21950 7044 21956 7046
rect 22012 7044 22036 7046
rect 22092 7044 22116 7046
rect 22172 7044 22196 7046
rect 22252 7044 22258 7046
rect 21950 7035 22258 7044
rect 21732 6724 21784 6730
rect 21732 6666 21784 6672
rect 21950 6012 22258 6021
rect 21950 6010 21956 6012
rect 22012 6010 22036 6012
rect 22092 6010 22116 6012
rect 22172 6010 22196 6012
rect 22252 6010 22258 6012
rect 22012 5958 22014 6010
rect 22194 5958 22196 6010
rect 21950 5956 21956 5958
rect 22012 5956 22036 5958
rect 22092 5956 22116 5958
rect 22172 5956 22196 5958
rect 22252 5956 22258 5958
rect 21950 5947 22258 5956
rect 22480 5234 22508 7890
rect 22610 7644 22918 7653
rect 22610 7642 22616 7644
rect 22672 7642 22696 7644
rect 22752 7642 22776 7644
rect 22832 7642 22856 7644
rect 22912 7642 22918 7644
rect 22672 7590 22674 7642
rect 22854 7590 22856 7642
rect 22610 7588 22616 7590
rect 22672 7588 22696 7590
rect 22752 7588 22776 7590
rect 22832 7588 22856 7590
rect 22912 7588 22918 7590
rect 22610 7579 22918 7588
rect 22610 6556 22918 6565
rect 22610 6554 22616 6556
rect 22672 6554 22696 6556
rect 22752 6554 22776 6556
rect 22832 6554 22856 6556
rect 22912 6554 22918 6556
rect 22672 6502 22674 6554
rect 22854 6502 22856 6554
rect 22610 6500 22616 6502
rect 22672 6500 22696 6502
rect 22752 6500 22776 6502
rect 22832 6500 22856 6502
rect 22912 6500 22918 6502
rect 22610 6491 22918 6500
rect 22610 5468 22918 5477
rect 22610 5466 22616 5468
rect 22672 5466 22696 5468
rect 22752 5466 22776 5468
rect 22832 5466 22856 5468
rect 22912 5466 22918 5468
rect 22672 5414 22674 5466
rect 22854 5414 22856 5466
rect 22610 5412 22616 5414
rect 22672 5412 22696 5414
rect 22752 5412 22776 5414
rect 22832 5412 22856 5414
rect 22912 5412 22918 5414
rect 22610 5403 22918 5412
rect 22468 5228 22520 5234
rect 22468 5170 22520 5176
rect 21950 4924 22258 4933
rect 21950 4922 21956 4924
rect 22012 4922 22036 4924
rect 22092 4922 22116 4924
rect 22172 4922 22196 4924
rect 22252 4922 22258 4924
rect 22012 4870 22014 4922
rect 22194 4870 22196 4922
rect 21950 4868 21956 4870
rect 22012 4868 22036 4870
rect 22092 4868 22116 4870
rect 22172 4868 22196 4870
rect 22252 4868 22258 4870
rect 21950 4859 22258 4868
rect 22610 4380 22918 4389
rect 22610 4378 22616 4380
rect 22672 4378 22696 4380
rect 22752 4378 22776 4380
rect 22832 4378 22856 4380
rect 22912 4378 22918 4380
rect 22672 4326 22674 4378
rect 22854 4326 22856 4378
rect 22610 4324 22616 4326
rect 22672 4324 22696 4326
rect 22752 4324 22776 4326
rect 22832 4324 22856 4326
rect 22912 4324 22918 4326
rect 22610 4315 22918 4324
rect 21950 3836 22258 3845
rect 21950 3834 21956 3836
rect 22012 3834 22036 3836
rect 22092 3834 22116 3836
rect 22172 3834 22196 3836
rect 22252 3834 22258 3836
rect 22012 3782 22014 3834
rect 22194 3782 22196 3834
rect 21950 3780 21956 3782
rect 22012 3780 22036 3782
rect 22092 3780 22116 3782
rect 22172 3780 22196 3782
rect 22252 3780 22258 3782
rect 21950 3771 22258 3780
rect 22610 3292 22918 3301
rect 22610 3290 22616 3292
rect 22672 3290 22696 3292
rect 22752 3290 22776 3292
rect 22832 3290 22856 3292
rect 22912 3290 22918 3292
rect 22672 3238 22674 3290
rect 22854 3238 22856 3290
rect 22610 3236 22616 3238
rect 22672 3236 22696 3238
rect 22752 3236 22776 3238
rect 22832 3236 22856 3238
rect 22912 3236 22918 3238
rect 22610 3227 22918 3236
rect 20076 2984 20128 2990
rect 20076 2926 20128 2932
rect 17316 2848 17368 2854
rect 17316 2790 17368 2796
rect 16950 2748 17258 2757
rect 16950 2746 16956 2748
rect 17012 2746 17036 2748
rect 17092 2746 17116 2748
rect 17172 2746 17196 2748
rect 17252 2746 17258 2748
rect 17012 2694 17014 2746
rect 17194 2694 17196 2746
rect 16950 2692 16956 2694
rect 17012 2692 17036 2694
rect 17092 2692 17116 2694
rect 17172 2692 17196 2694
rect 17252 2692 17258 2694
rect 16950 2683 17258 2692
rect 21950 2748 22258 2757
rect 21950 2746 21956 2748
rect 22012 2746 22036 2748
rect 22092 2746 22116 2748
rect 22172 2746 22196 2748
rect 22252 2746 22258 2748
rect 22012 2694 22014 2746
rect 22194 2694 22196 2746
rect 21950 2692 21956 2694
rect 22012 2692 22036 2694
rect 22092 2692 22116 2694
rect 22172 2692 22196 2694
rect 22252 2692 22258 2694
rect 21950 2683 22258 2692
rect 24596 2650 24624 20266
rect 24688 19514 24716 20334
rect 24676 19508 24728 19514
rect 24676 19450 24728 19456
rect 24872 16046 24900 20454
rect 24952 16584 25004 16590
rect 24952 16526 25004 16532
rect 24860 16040 24912 16046
rect 24860 15982 24912 15988
rect 24858 12200 24914 12209
rect 24858 12135 24914 12144
rect 24872 7750 24900 12135
rect 24860 7744 24912 7750
rect 24860 7686 24912 7692
rect 24964 7342 24992 16526
rect 24952 7336 25004 7342
rect 24952 7278 25004 7284
rect 25240 6322 25268 37878
rect 25700 37874 25728 42298
rect 25884 41138 25912 46922
rect 25964 43648 26016 43654
rect 25964 43590 26016 43596
rect 25872 41132 25924 41138
rect 25872 41074 25924 41080
rect 25872 39432 25924 39438
rect 25872 39374 25924 39380
rect 25884 38282 25912 39374
rect 25872 38276 25924 38282
rect 25872 38218 25924 38224
rect 25688 37868 25740 37874
rect 25688 37810 25740 37816
rect 25504 37800 25556 37806
rect 25504 37742 25556 37748
rect 25516 37398 25544 37742
rect 25504 37392 25556 37398
rect 25504 37334 25556 37340
rect 25412 34196 25464 34202
rect 25412 34138 25464 34144
rect 25424 33522 25452 34138
rect 25412 33516 25464 33522
rect 25412 33458 25464 33464
rect 25516 31754 25544 37334
rect 25424 31726 25544 31754
rect 25320 28960 25372 28966
rect 25320 28902 25372 28908
rect 25332 28490 25360 28902
rect 25320 28484 25372 28490
rect 25320 28426 25372 28432
rect 25332 25974 25360 28426
rect 25320 25968 25372 25974
rect 25320 25910 25372 25916
rect 25424 18290 25452 31726
rect 25596 29572 25648 29578
rect 25596 29514 25648 29520
rect 25608 18902 25636 29514
rect 25596 18896 25648 18902
rect 25596 18838 25648 18844
rect 25412 18284 25464 18290
rect 25412 18226 25464 18232
rect 25608 16590 25636 18838
rect 25700 18222 25728 37810
rect 25884 35086 25912 38218
rect 25872 35080 25924 35086
rect 25872 35022 25924 35028
rect 25872 33516 25924 33522
rect 25872 33458 25924 33464
rect 25884 23866 25912 33458
rect 25976 28966 26004 43590
rect 26068 42158 26096 48286
rect 26056 42152 26108 42158
rect 26056 42094 26108 42100
rect 26068 29714 26096 42094
rect 26160 39438 26188 50798
rect 26804 42226 26832 53450
rect 26950 52796 27258 52805
rect 26950 52794 26956 52796
rect 27012 52794 27036 52796
rect 27092 52794 27116 52796
rect 27172 52794 27196 52796
rect 27252 52794 27258 52796
rect 27012 52742 27014 52794
rect 27194 52742 27196 52794
rect 26950 52740 26956 52742
rect 27012 52740 27036 52742
rect 27092 52740 27116 52742
rect 27172 52740 27196 52742
rect 27252 52740 27258 52742
rect 26950 52731 27258 52740
rect 26950 51708 27258 51717
rect 26950 51706 26956 51708
rect 27012 51706 27036 51708
rect 27092 51706 27116 51708
rect 27172 51706 27196 51708
rect 27252 51706 27258 51708
rect 27012 51654 27014 51706
rect 27194 51654 27196 51706
rect 26950 51652 26956 51654
rect 27012 51652 27036 51654
rect 27092 51652 27116 51654
rect 27172 51652 27196 51654
rect 27252 51652 27258 51654
rect 26950 51643 27258 51652
rect 26950 50620 27258 50629
rect 26950 50618 26956 50620
rect 27012 50618 27036 50620
rect 27092 50618 27116 50620
rect 27172 50618 27196 50620
rect 27252 50618 27258 50620
rect 27012 50566 27014 50618
rect 27194 50566 27196 50618
rect 26950 50564 26956 50566
rect 27012 50564 27036 50566
rect 27092 50564 27116 50566
rect 27172 50564 27196 50566
rect 27252 50564 27258 50566
rect 26950 50555 27258 50564
rect 26950 49532 27258 49541
rect 26950 49530 26956 49532
rect 27012 49530 27036 49532
rect 27092 49530 27116 49532
rect 27172 49530 27196 49532
rect 27252 49530 27258 49532
rect 27012 49478 27014 49530
rect 27194 49478 27196 49530
rect 26950 49476 26956 49478
rect 27012 49476 27036 49478
rect 27092 49476 27116 49478
rect 27172 49476 27196 49478
rect 27252 49476 27258 49478
rect 26950 49467 27258 49476
rect 26950 48444 27258 48453
rect 26950 48442 26956 48444
rect 27012 48442 27036 48444
rect 27092 48442 27116 48444
rect 27172 48442 27196 48444
rect 27252 48442 27258 48444
rect 27012 48390 27014 48442
rect 27194 48390 27196 48442
rect 26950 48388 26956 48390
rect 27012 48388 27036 48390
rect 27092 48388 27116 48390
rect 27172 48388 27196 48390
rect 27252 48388 27258 48390
rect 26950 48379 27258 48388
rect 26950 47356 27258 47365
rect 26950 47354 26956 47356
rect 27012 47354 27036 47356
rect 27092 47354 27116 47356
rect 27172 47354 27196 47356
rect 27252 47354 27258 47356
rect 27012 47302 27014 47354
rect 27194 47302 27196 47354
rect 26950 47300 26956 47302
rect 27012 47300 27036 47302
rect 27092 47300 27116 47302
rect 27172 47300 27196 47302
rect 27252 47300 27258 47302
rect 26950 47291 27258 47300
rect 26950 46268 27258 46277
rect 26950 46266 26956 46268
rect 27012 46266 27036 46268
rect 27092 46266 27116 46268
rect 27172 46266 27196 46268
rect 27252 46266 27258 46268
rect 27012 46214 27014 46266
rect 27194 46214 27196 46266
rect 26950 46212 26956 46214
rect 27012 46212 27036 46214
rect 27092 46212 27116 46214
rect 27172 46212 27196 46214
rect 27252 46212 27258 46214
rect 26950 46203 27258 46212
rect 26950 45180 27258 45189
rect 26950 45178 26956 45180
rect 27012 45178 27036 45180
rect 27092 45178 27116 45180
rect 27172 45178 27196 45180
rect 27252 45178 27258 45180
rect 27012 45126 27014 45178
rect 27194 45126 27196 45178
rect 26950 45124 26956 45126
rect 27012 45124 27036 45126
rect 27092 45124 27116 45126
rect 27172 45124 27196 45126
rect 27252 45124 27258 45126
rect 26950 45115 27258 45124
rect 26884 44940 26936 44946
rect 26884 44882 26936 44888
rect 26896 44470 26924 44882
rect 26884 44464 26936 44470
rect 26884 44406 26936 44412
rect 26950 44092 27258 44101
rect 26950 44090 26956 44092
rect 27012 44090 27036 44092
rect 27092 44090 27116 44092
rect 27172 44090 27196 44092
rect 27252 44090 27258 44092
rect 27012 44038 27014 44090
rect 27194 44038 27196 44090
rect 26950 44036 26956 44038
rect 27012 44036 27036 44038
rect 27092 44036 27116 44038
rect 27172 44036 27196 44038
rect 27252 44036 27258 44038
rect 26950 44027 27258 44036
rect 26950 43004 27258 43013
rect 26950 43002 26956 43004
rect 27012 43002 27036 43004
rect 27092 43002 27116 43004
rect 27172 43002 27196 43004
rect 27252 43002 27258 43004
rect 27012 42950 27014 43002
rect 27194 42950 27196 43002
rect 26950 42948 26956 42950
rect 27012 42948 27036 42950
rect 27092 42948 27116 42950
rect 27172 42948 27196 42950
rect 27252 42948 27258 42950
rect 26950 42939 27258 42948
rect 26332 42220 26384 42226
rect 26332 42162 26384 42168
rect 26792 42220 26844 42226
rect 26792 42162 26844 42168
rect 27344 42220 27396 42226
rect 27344 42162 27396 42168
rect 26240 39568 26292 39574
rect 26240 39510 26292 39516
rect 26148 39432 26200 39438
rect 26148 39374 26200 39380
rect 26160 35698 26188 39374
rect 26252 39030 26280 39510
rect 26240 39024 26292 39030
rect 26240 38966 26292 38972
rect 26148 35692 26200 35698
rect 26148 35634 26200 35640
rect 26160 33522 26188 35634
rect 26148 33516 26200 33522
rect 26148 33458 26200 33464
rect 26056 29708 26108 29714
rect 26056 29650 26108 29656
rect 25964 28960 26016 28966
rect 25964 28902 26016 28908
rect 26056 25696 26108 25702
rect 26056 25638 26108 25644
rect 26068 24138 26096 25638
rect 26344 24818 26372 42162
rect 26424 42016 26476 42022
rect 26424 41958 26476 41964
rect 26332 24812 26384 24818
rect 26332 24754 26384 24760
rect 26056 24132 26108 24138
rect 26056 24074 26108 24080
rect 26148 24132 26200 24138
rect 26148 24074 26200 24080
rect 25872 23860 25924 23866
rect 25872 23802 25924 23808
rect 25688 18216 25740 18222
rect 25688 18158 25740 18164
rect 25596 16584 25648 16590
rect 25596 16526 25648 16532
rect 25228 6316 25280 6322
rect 25228 6258 25280 6264
rect 26068 3398 26096 24074
rect 26160 24018 26188 24074
rect 26332 24064 26384 24070
rect 26160 23990 26280 24018
rect 26332 24006 26384 24012
rect 26148 23860 26200 23866
rect 26148 23802 26200 23808
rect 26160 22030 26188 23802
rect 26252 23746 26280 23990
rect 26344 23866 26372 24006
rect 26332 23860 26384 23866
rect 26332 23802 26384 23808
rect 26252 23718 26372 23746
rect 26344 23594 26372 23718
rect 26332 23588 26384 23594
rect 26332 23530 26384 23536
rect 26240 22092 26292 22098
rect 26240 22034 26292 22040
rect 26148 22024 26200 22030
rect 26148 21966 26200 21972
rect 26252 18766 26280 22034
rect 26240 18760 26292 18766
rect 26240 18702 26292 18708
rect 26056 3392 26108 3398
rect 26056 3334 26108 3340
rect 26344 2922 26372 23530
rect 26436 18766 26464 41958
rect 26950 41916 27258 41925
rect 26950 41914 26956 41916
rect 27012 41914 27036 41916
rect 27092 41914 27116 41916
rect 27172 41914 27196 41916
rect 27252 41914 27258 41916
rect 27012 41862 27014 41914
rect 27194 41862 27196 41914
rect 26950 41860 26956 41862
rect 27012 41860 27036 41862
rect 27092 41860 27116 41862
rect 27172 41860 27196 41862
rect 27252 41860 27258 41862
rect 26950 41851 27258 41860
rect 27356 41818 27384 42162
rect 27344 41812 27396 41818
rect 27344 41754 27396 41760
rect 26950 40828 27258 40837
rect 26950 40826 26956 40828
rect 27012 40826 27036 40828
rect 27092 40826 27116 40828
rect 27172 40826 27196 40828
rect 27252 40826 27258 40828
rect 27012 40774 27014 40826
rect 27194 40774 27196 40826
rect 26950 40772 26956 40774
rect 27012 40772 27036 40774
rect 27092 40772 27116 40774
rect 27172 40772 27196 40774
rect 27252 40772 27258 40774
rect 26950 40763 27258 40772
rect 26950 39740 27258 39749
rect 26950 39738 26956 39740
rect 27012 39738 27036 39740
rect 27092 39738 27116 39740
rect 27172 39738 27196 39740
rect 27252 39738 27258 39740
rect 27012 39686 27014 39738
rect 27194 39686 27196 39738
rect 26950 39684 26956 39686
rect 27012 39684 27036 39686
rect 27092 39684 27116 39686
rect 27172 39684 27196 39686
rect 27252 39684 27258 39686
rect 26950 39675 27258 39684
rect 26950 38652 27258 38661
rect 26950 38650 26956 38652
rect 27012 38650 27036 38652
rect 27092 38650 27116 38652
rect 27172 38650 27196 38652
rect 27252 38650 27258 38652
rect 27012 38598 27014 38650
rect 27194 38598 27196 38650
rect 26950 38596 26956 38598
rect 27012 38596 27036 38598
rect 27092 38596 27116 38598
rect 27172 38596 27196 38598
rect 27252 38596 27258 38598
rect 26950 38587 27258 38596
rect 27448 37874 27476 58890
rect 27540 58138 27568 59910
rect 27610 59868 27918 59877
rect 27610 59866 27616 59868
rect 27672 59866 27696 59868
rect 27752 59866 27776 59868
rect 27832 59866 27856 59868
rect 27912 59866 27918 59868
rect 27672 59814 27674 59866
rect 27854 59814 27856 59866
rect 27610 59812 27616 59814
rect 27672 59812 27696 59814
rect 27752 59812 27776 59814
rect 27832 59812 27856 59814
rect 27912 59812 27918 59814
rect 27610 59803 27918 59812
rect 27610 58780 27918 58789
rect 27610 58778 27616 58780
rect 27672 58778 27696 58780
rect 27752 58778 27776 58780
rect 27832 58778 27856 58780
rect 27912 58778 27918 58780
rect 27672 58726 27674 58778
rect 27854 58726 27856 58778
rect 27610 58724 27616 58726
rect 27672 58724 27696 58726
rect 27752 58724 27776 58726
rect 27832 58724 27856 58726
rect 27912 58724 27918 58726
rect 27610 58715 27918 58724
rect 27528 58132 27580 58138
rect 27528 58074 27580 58080
rect 27528 57792 27580 57798
rect 27528 57734 27580 57740
rect 26792 37868 26844 37874
rect 26792 37810 26844 37816
rect 27436 37868 27488 37874
rect 27436 37810 27488 37816
rect 26608 37392 26660 37398
rect 26608 37334 26660 37340
rect 26620 36854 26648 37334
rect 26608 36848 26660 36854
rect 26608 36790 26660 36796
rect 26620 36530 26648 36790
rect 26620 36502 26740 36530
rect 26608 35692 26660 35698
rect 26608 35634 26660 35640
rect 26620 34950 26648 35634
rect 26608 34944 26660 34950
rect 26608 34886 26660 34892
rect 26516 26852 26568 26858
rect 26516 26794 26568 26800
rect 26528 24070 26556 26794
rect 26516 24064 26568 24070
rect 26516 24006 26568 24012
rect 26424 18760 26476 18766
rect 26424 18702 26476 18708
rect 26528 14482 26556 24006
rect 26620 18766 26648 34886
rect 26608 18760 26660 18766
rect 26608 18702 26660 18708
rect 26620 14822 26648 18702
rect 26608 14816 26660 14822
rect 26608 14758 26660 14764
rect 26516 14476 26568 14482
rect 26516 14418 26568 14424
rect 26712 8974 26740 36502
rect 26700 8968 26752 8974
rect 26700 8910 26752 8916
rect 26424 8900 26476 8906
rect 26424 8842 26476 8848
rect 26436 4690 26464 8842
rect 26804 8090 26832 37810
rect 26950 37564 27258 37573
rect 26950 37562 26956 37564
rect 27012 37562 27036 37564
rect 27092 37562 27116 37564
rect 27172 37562 27196 37564
rect 27252 37562 27258 37564
rect 27012 37510 27014 37562
rect 27194 37510 27196 37562
rect 26950 37508 26956 37510
rect 27012 37508 27036 37510
rect 27092 37508 27116 37510
rect 27172 37508 27196 37510
rect 27252 37508 27258 37510
rect 26950 37499 27258 37508
rect 26950 36476 27258 36485
rect 26950 36474 26956 36476
rect 27012 36474 27036 36476
rect 27092 36474 27116 36476
rect 27172 36474 27196 36476
rect 27252 36474 27258 36476
rect 27012 36422 27014 36474
rect 27194 36422 27196 36474
rect 26950 36420 26956 36422
rect 27012 36420 27036 36422
rect 27092 36420 27116 36422
rect 27172 36420 27196 36422
rect 27252 36420 27258 36422
rect 26950 36411 27258 36420
rect 26950 35388 27258 35397
rect 26950 35386 26956 35388
rect 27012 35386 27036 35388
rect 27092 35386 27116 35388
rect 27172 35386 27196 35388
rect 27252 35386 27258 35388
rect 27012 35334 27014 35386
rect 27194 35334 27196 35386
rect 26950 35332 26956 35334
rect 27012 35332 27036 35334
rect 27092 35332 27116 35334
rect 27172 35332 27196 35334
rect 27252 35332 27258 35334
rect 26950 35323 27258 35332
rect 26950 34300 27258 34309
rect 26950 34298 26956 34300
rect 27012 34298 27036 34300
rect 27092 34298 27116 34300
rect 27172 34298 27196 34300
rect 27252 34298 27258 34300
rect 27012 34246 27014 34298
rect 27194 34246 27196 34298
rect 26950 34244 26956 34246
rect 27012 34244 27036 34246
rect 27092 34244 27116 34246
rect 27172 34244 27196 34246
rect 27252 34244 27258 34246
rect 26950 34235 27258 34244
rect 26950 33212 27258 33221
rect 26950 33210 26956 33212
rect 27012 33210 27036 33212
rect 27092 33210 27116 33212
rect 27172 33210 27196 33212
rect 27252 33210 27258 33212
rect 27012 33158 27014 33210
rect 27194 33158 27196 33210
rect 26950 33156 26956 33158
rect 27012 33156 27036 33158
rect 27092 33156 27116 33158
rect 27172 33156 27196 33158
rect 27252 33156 27258 33158
rect 26950 33147 27258 33156
rect 26950 32124 27258 32133
rect 26950 32122 26956 32124
rect 27012 32122 27036 32124
rect 27092 32122 27116 32124
rect 27172 32122 27196 32124
rect 27252 32122 27258 32124
rect 27012 32070 27014 32122
rect 27194 32070 27196 32122
rect 26950 32068 26956 32070
rect 27012 32068 27036 32070
rect 27092 32068 27116 32070
rect 27172 32068 27196 32070
rect 27252 32068 27258 32070
rect 26950 32059 27258 32068
rect 27344 31816 27396 31822
rect 27344 31758 27396 31764
rect 26950 31036 27258 31045
rect 26950 31034 26956 31036
rect 27012 31034 27036 31036
rect 27092 31034 27116 31036
rect 27172 31034 27196 31036
rect 27252 31034 27258 31036
rect 27012 30982 27014 31034
rect 27194 30982 27196 31034
rect 26950 30980 26956 30982
rect 27012 30980 27036 30982
rect 27092 30980 27116 30982
rect 27172 30980 27196 30982
rect 27252 30980 27258 30982
rect 26950 30971 27258 30980
rect 26950 29948 27258 29957
rect 26950 29946 26956 29948
rect 27012 29946 27036 29948
rect 27092 29946 27116 29948
rect 27172 29946 27196 29948
rect 27252 29946 27258 29948
rect 27012 29894 27014 29946
rect 27194 29894 27196 29946
rect 26950 29892 26956 29894
rect 27012 29892 27036 29894
rect 27092 29892 27116 29894
rect 27172 29892 27196 29894
rect 27252 29892 27258 29894
rect 26950 29883 27258 29892
rect 26950 28860 27258 28869
rect 26950 28858 26956 28860
rect 27012 28858 27036 28860
rect 27092 28858 27116 28860
rect 27172 28858 27196 28860
rect 27252 28858 27258 28860
rect 27012 28806 27014 28858
rect 27194 28806 27196 28858
rect 26950 28804 26956 28806
rect 27012 28804 27036 28806
rect 27092 28804 27116 28806
rect 27172 28804 27196 28806
rect 27252 28804 27258 28806
rect 26950 28795 27258 28804
rect 26950 27772 27258 27781
rect 26950 27770 26956 27772
rect 27012 27770 27036 27772
rect 27092 27770 27116 27772
rect 27172 27770 27196 27772
rect 27252 27770 27258 27772
rect 27012 27718 27014 27770
rect 27194 27718 27196 27770
rect 26950 27716 26956 27718
rect 27012 27716 27036 27718
rect 27092 27716 27116 27718
rect 27172 27716 27196 27718
rect 27252 27716 27258 27718
rect 26950 27707 27258 27716
rect 26950 26684 27258 26693
rect 26950 26682 26956 26684
rect 27012 26682 27036 26684
rect 27092 26682 27116 26684
rect 27172 26682 27196 26684
rect 27252 26682 27258 26684
rect 27012 26630 27014 26682
rect 27194 26630 27196 26682
rect 26950 26628 26956 26630
rect 27012 26628 27036 26630
rect 27092 26628 27116 26630
rect 27172 26628 27196 26630
rect 27252 26628 27258 26630
rect 26950 26619 27258 26628
rect 26950 25596 27258 25605
rect 26950 25594 26956 25596
rect 27012 25594 27036 25596
rect 27092 25594 27116 25596
rect 27172 25594 27196 25596
rect 27252 25594 27258 25596
rect 27012 25542 27014 25594
rect 27194 25542 27196 25594
rect 26950 25540 26956 25542
rect 27012 25540 27036 25542
rect 27092 25540 27116 25542
rect 27172 25540 27196 25542
rect 27252 25540 27258 25542
rect 26950 25531 27258 25540
rect 27356 25106 27384 31758
rect 27448 30734 27476 37810
rect 27436 30728 27488 30734
rect 27436 30670 27488 30676
rect 27448 29578 27476 30670
rect 27436 29572 27488 29578
rect 27436 29514 27488 29520
rect 27264 25078 27384 25106
rect 27264 24698 27292 25078
rect 27540 24954 27568 57734
rect 27610 57692 27918 57701
rect 27610 57690 27616 57692
rect 27672 57690 27696 57692
rect 27752 57690 27776 57692
rect 27832 57690 27856 57692
rect 27912 57690 27918 57692
rect 27672 57638 27674 57690
rect 27854 57638 27856 57690
rect 27610 57636 27616 57638
rect 27672 57636 27696 57638
rect 27752 57636 27776 57638
rect 27832 57636 27856 57638
rect 27912 57636 27918 57638
rect 27610 57627 27918 57636
rect 27610 56604 27918 56613
rect 27610 56602 27616 56604
rect 27672 56602 27696 56604
rect 27752 56602 27776 56604
rect 27832 56602 27856 56604
rect 27912 56602 27918 56604
rect 27672 56550 27674 56602
rect 27854 56550 27856 56602
rect 27610 56548 27616 56550
rect 27672 56548 27696 56550
rect 27752 56548 27776 56550
rect 27832 56548 27856 56550
rect 27912 56548 27918 56550
rect 27610 56539 27918 56548
rect 27610 55516 27918 55525
rect 27610 55514 27616 55516
rect 27672 55514 27696 55516
rect 27752 55514 27776 55516
rect 27832 55514 27856 55516
rect 27912 55514 27918 55516
rect 27672 55462 27674 55514
rect 27854 55462 27856 55514
rect 27610 55460 27616 55462
rect 27672 55460 27696 55462
rect 27752 55460 27776 55462
rect 27832 55460 27856 55462
rect 27912 55460 27918 55462
rect 27610 55451 27918 55460
rect 27610 54428 27918 54437
rect 27610 54426 27616 54428
rect 27672 54426 27696 54428
rect 27752 54426 27776 54428
rect 27832 54426 27856 54428
rect 27912 54426 27918 54428
rect 27672 54374 27674 54426
rect 27854 54374 27856 54426
rect 27610 54372 27616 54374
rect 27672 54372 27696 54374
rect 27752 54372 27776 54374
rect 27832 54372 27856 54374
rect 27912 54372 27918 54374
rect 27610 54363 27918 54372
rect 27610 53340 27918 53349
rect 27610 53338 27616 53340
rect 27672 53338 27696 53340
rect 27752 53338 27776 53340
rect 27832 53338 27856 53340
rect 27912 53338 27918 53340
rect 27672 53286 27674 53338
rect 27854 53286 27856 53338
rect 27610 53284 27616 53286
rect 27672 53284 27696 53286
rect 27752 53284 27776 53286
rect 27832 53284 27856 53286
rect 27912 53284 27918 53286
rect 27610 53275 27918 53284
rect 27610 52252 27918 52261
rect 27610 52250 27616 52252
rect 27672 52250 27696 52252
rect 27752 52250 27776 52252
rect 27832 52250 27856 52252
rect 27912 52250 27918 52252
rect 27672 52198 27674 52250
rect 27854 52198 27856 52250
rect 27610 52196 27616 52198
rect 27672 52196 27696 52198
rect 27752 52196 27776 52198
rect 27832 52196 27856 52198
rect 27912 52196 27918 52198
rect 27610 52187 27918 52196
rect 27610 51164 27918 51173
rect 27610 51162 27616 51164
rect 27672 51162 27696 51164
rect 27752 51162 27776 51164
rect 27832 51162 27856 51164
rect 27912 51162 27918 51164
rect 27672 51110 27674 51162
rect 27854 51110 27856 51162
rect 27610 51108 27616 51110
rect 27672 51108 27696 51110
rect 27752 51108 27776 51110
rect 27832 51108 27856 51110
rect 27912 51108 27918 51110
rect 27610 51099 27918 51108
rect 27610 50076 27918 50085
rect 27610 50074 27616 50076
rect 27672 50074 27696 50076
rect 27752 50074 27776 50076
rect 27832 50074 27856 50076
rect 27912 50074 27918 50076
rect 27672 50022 27674 50074
rect 27854 50022 27856 50074
rect 27610 50020 27616 50022
rect 27672 50020 27696 50022
rect 27752 50020 27776 50022
rect 27832 50020 27856 50022
rect 27912 50020 27918 50022
rect 27610 50011 27918 50020
rect 27610 48988 27918 48997
rect 27610 48986 27616 48988
rect 27672 48986 27696 48988
rect 27752 48986 27776 48988
rect 27832 48986 27856 48988
rect 27912 48986 27918 48988
rect 27672 48934 27674 48986
rect 27854 48934 27856 48986
rect 27610 48932 27616 48934
rect 27672 48932 27696 48934
rect 27752 48932 27776 48934
rect 27832 48932 27856 48934
rect 27912 48932 27918 48934
rect 27610 48923 27918 48932
rect 27610 47900 27918 47909
rect 27610 47898 27616 47900
rect 27672 47898 27696 47900
rect 27752 47898 27776 47900
rect 27832 47898 27856 47900
rect 27912 47898 27918 47900
rect 27672 47846 27674 47898
rect 27854 47846 27856 47898
rect 27610 47844 27616 47846
rect 27672 47844 27696 47846
rect 27752 47844 27776 47846
rect 27832 47844 27856 47846
rect 27912 47844 27918 47846
rect 27610 47835 27918 47844
rect 28000 47666 28028 63174
rect 28264 62280 28316 62286
rect 28264 62222 28316 62228
rect 28080 57928 28132 57934
rect 28080 57870 28132 57876
rect 28092 55214 28120 57870
rect 28092 55186 28212 55214
rect 28080 54188 28132 54194
rect 28080 54130 28132 54136
rect 27988 47660 28040 47666
rect 27988 47602 28040 47608
rect 27610 46812 27918 46821
rect 27610 46810 27616 46812
rect 27672 46810 27696 46812
rect 27752 46810 27776 46812
rect 27832 46810 27856 46812
rect 27912 46810 27918 46812
rect 27672 46758 27674 46810
rect 27854 46758 27856 46810
rect 27610 46756 27616 46758
rect 27672 46756 27696 46758
rect 27752 46756 27776 46758
rect 27832 46756 27856 46758
rect 27912 46756 27918 46758
rect 27610 46747 27918 46756
rect 27610 45724 27918 45733
rect 27610 45722 27616 45724
rect 27672 45722 27696 45724
rect 27752 45722 27776 45724
rect 27832 45722 27856 45724
rect 27912 45722 27918 45724
rect 27672 45670 27674 45722
rect 27854 45670 27856 45722
rect 27610 45668 27616 45670
rect 27672 45668 27696 45670
rect 27752 45668 27776 45670
rect 27832 45668 27856 45670
rect 27912 45668 27918 45670
rect 27610 45659 27918 45668
rect 27610 44636 27918 44645
rect 27610 44634 27616 44636
rect 27672 44634 27696 44636
rect 27752 44634 27776 44636
rect 27832 44634 27856 44636
rect 27912 44634 27918 44636
rect 27672 44582 27674 44634
rect 27854 44582 27856 44634
rect 27610 44580 27616 44582
rect 27672 44580 27696 44582
rect 27752 44580 27776 44582
rect 27832 44580 27856 44582
rect 27912 44580 27918 44582
rect 27610 44571 27918 44580
rect 27610 43548 27918 43557
rect 27610 43546 27616 43548
rect 27672 43546 27696 43548
rect 27752 43546 27776 43548
rect 27832 43546 27856 43548
rect 27912 43546 27918 43548
rect 27672 43494 27674 43546
rect 27854 43494 27856 43546
rect 27610 43492 27616 43494
rect 27672 43492 27696 43494
rect 27752 43492 27776 43494
rect 27832 43492 27856 43494
rect 27912 43492 27918 43494
rect 27610 43483 27918 43492
rect 27988 43308 28040 43314
rect 27988 43250 28040 43256
rect 27610 42460 27918 42469
rect 27610 42458 27616 42460
rect 27672 42458 27696 42460
rect 27752 42458 27776 42460
rect 27832 42458 27856 42460
rect 27912 42458 27918 42460
rect 27672 42406 27674 42458
rect 27854 42406 27856 42458
rect 27610 42404 27616 42406
rect 27672 42404 27696 42406
rect 27752 42404 27776 42406
rect 27832 42404 27856 42406
rect 27912 42404 27918 42406
rect 27610 42395 27918 42404
rect 28000 42294 28028 43250
rect 27988 42288 28040 42294
rect 27988 42230 28040 42236
rect 27610 41372 27918 41381
rect 27610 41370 27616 41372
rect 27672 41370 27696 41372
rect 27752 41370 27776 41372
rect 27832 41370 27856 41372
rect 27912 41370 27918 41372
rect 27672 41318 27674 41370
rect 27854 41318 27856 41370
rect 27610 41316 27616 41318
rect 27672 41316 27696 41318
rect 27752 41316 27776 41318
rect 27832 41316 27856 41318
rect 27912 41316 27918 41318
rect 27610 41307 27918 41316
rect 27988 41132 28040 41138
rect 27988 41074 28040 41080
rect 27610 40284 27918 40293
rect 27610 40282 27616 40284
rect 27672 40282 27696 40284
rect 27752 40282 27776 40284
rect 27832 40282 27856 40284
rect 27912 40282 27918 40284
rect 27672 40230 27674 40282
rect 27854 40230 27856 40282
rect 27610 40228 27616 40230
rect 27672 40228 27696 40230
rect 27752 40228 27776 40230
rect 27832 40228 27856 40230
rect 27912 40228 27918 40230
rect 27610 40219 27918 40228
rect 27610 39196 27918 39205
rect 27610 39194 27616 39196
rect 27672 39194 27696 39196
rect 27752 39194 27776 39196
rect 27832 39194 27856 39196
rect 27912 39194 27918 39196
rect 27672 39142 27674 39194
rect 27854 39142 27856 39194
rect 27610 39140 27616 39142
rect 27672 39140 27696 39142
rect 27752 39140 27776 39142
rect 27832 39140 27856 39142
rect 27912 39140 27918 39142
rect 27610 39131 27918 39140
rect 27610 38108 27918 38117
rect 27610 38106 27616 38108
rect 27672 38106 27696 38108
rect 27752 38106 27776 38108
rect 27832 38106 27856 38108
rect 27912 38106 27918 38108
rect 27672 38054 27674 38106
rect 27854 38054 27856 38106
rect 27610 38052 27616 38054
rect 27672 38052 27696 38054
rect 27752 38052 27776 38054
rect 27832 38052 27856 38054
rect 27912 38052 27918 38054
rect 27610 38043 27918 38052
rect 27610 37020 27918 37029
rect 27610 37018 27616 37020
rect 27672 37018 27696 37020
rect 27752 37018 27776 37020
rect 27832 37018 27856 37020
rect 27912 37018 27918 37020
rect 27672 36966 27674 37018
rect 27854 36966 27856 37018
rect 27610 36964 27616 36966
rect 27672 36964 27696 36966
rect 27752 36964 27776 36966
rect 27832 36964 27856 36966
rect 27912 36964 27918 36966
rect 27610 36955 27918 36964
rect 27610 35932 27918 35941
rect 27610 35930 27616 35932
rect 27672 35930 27696 35932
rect 27752 35930 27776 35932
rect 27832 35930 27856 35932
rect 27912 35930 27918 35932
rect 27672 35878 27674 35930
rect 27854 35878 27856 35930
rect 27610 35876 27616 35878
rect 27672 35876 27696 35878
rect 27752 35876 27776 35878
rect 27832 35876 27856 35878
rect 27912 35876 27918 35878
rect 27610 35867 27918 35876
rect 27610 34844 27918 34853
rect 27610 34842 27616 34844
rect 27672 34842 27696 34844
rect 27752 34842 27776 34844
rect 27832 34842 27856 34844
rect 27912 34842 27918 34844
rect 27672 34790 27674 34842
rect 27854 34790 27856 34842
rect 27610 34788 27616 34790
rect 27672 34788 27696 34790
rect 27752 34788 27776 34790
rect 27832 34788 27856 34790
rect 27912 34788 27918 34790
rect 27610 34779 27918 34788
rect 28000 33862 28028 41074
rect 28092 37466 28120 54130
rect 28184 47598 28212 55186
rect 28276 54194 28304 62222
rect 28264 54188 28316 54194
rect 28264 54130 28316 54136
rect 28356 53984 28408 53990
rect 28356 53926 28408 53932
rect 28172 47592 28224 47598
rect 28172 47534 28224 47540
rect 28264 41540 28316 41546
rect 28264 41482 28316 41488
rect 28080 37460 28132 37466
rect 28080 37402 28132 37408
rect 28276 36174 28304 41482
rect 28368 41478 28396 53926
rect 28448 53440 28500 53446
rect 28448 53382 28500 53388
rect 28356 41472 28408 41478
rect 28356 41414 28408 41420
rect 28264 36168 28316 36174
rect 28264 36110 28316 36116
rect 27988 33856 28040 33862
rect 27988 33798 28040 33804
rect 27610 33756 27918 33765
rect 27610 33754 27616 33756
rect 27672 33754 27696 33756
rect 27752 33754 27776 33756
rect 27832 33754 27856 33756
rect 27912 33754 27918 33756
rect 27672 33702 27674 33754
rect 27854 33702 27856 33754
rect 27610 33700 27616 33702
rect 27672 33700 27696 33702
rect 27752 33700 27776 33702
rect 27832 33700 27856 33702
rect 27912 33700 27918 33702
rect 27610 33691 27918 33700
rect 27610 32668 27918 32677
rect 27610 32666 27616 32668
rect 27672 32666 27696 32668
rect 27752 32666 27776 32668
rect 27832 32666 27856 32668
rect 27912 32666 27918 32668
rect 27672 32614 27674 32666
rect 27854 32614 27856 32666
rect 27610 32612 27616 32614
rect 27672 32612 27696 32614
rect 27752 32612 27776 32614
rect 27832 32612 27856 32614
rect 27912 32612 27918 32614
rect 27610 32603 27918 32612
rect 27610 31580 27918 31589
rect 27610 31578 27616 31580
rect 27672 31578 27696 31580
rect 27752 31578 27776 31580
rect 27832 31578 27856 31580
rect 27912 31578 27918 31580
rect 27672 31526 27674 31578
rect 27854 31526 27856 31578
rect 27610 31524 27616 31526
rect 27672 31524 27696 31526
rect 27752 31524 27776 31526
rect 27832 31524 27856 31526
rect 27912 31524 27918 31526
rect 27610 31515 27918 31524
rect 27610 30492 27918 30501
rect 27610 30490 27616 30492
rect 27672 30490 27696 30492
rect 27752 30490 27776 30492
rect 27832 30490 27856 30492
rect 27912 30490 27918 30492
rect 27672 30438 27674 30490
rect 27854 30438 27856 30490
rect 27610 30436 27616 30438
rect 27672 30436 27696 30438
rect 27752 30436 27776 30438
rect 27832 30436 27856 30438
rect 27912 30436 27918 30438
rect 27610 30427 27918 30436
rect 27610 29404 27918 29413
rect 27610 29402 27616 29404
rect 27672 29402 27696 29404
rect 27752 29402 27776 29404
rect 27832 29402 27856 29404
rect 27912 29402 27918 29404
rect 27672 29350 27674 29402
rect 27854 29350 27856 29402
rect 27610 29348 27616 29350
rect 27672 29348 27696 29350
rect 27752 29348 27776 29350
rect 27832 29348 27856 29350
rect 27912 29348 27918 29350
rect 27610 29339 27918 29348
rect 27610 28316 27918 28325
rect 27610 28314 27616 28316
rect 27672 28314 27696 28316
rect 27752 28314 27776 28316
rect 27832 28314 27856 28316
rect 27912 28314 27918 28316
rect 27672 28262 27674 28314
rect 27854 28262 27856 28314
rect 27610 28260 27616 28262
rect 27672 28260 27696 28262
rect 27752 28260 27776 28262
rect 27832 28260 27856 28262
rect 27912 28260 27918 28262
rect 27610 28251 27918 28260
rect 27610 27228 27918 27237
rect 27610 27226 27616 27228
rect 27672 27226 27696 27228
rect 27752 27226 27776 27228
rect 27832 27226 27856 27228
rect 27912 27226 27918 27228
rect 27672 27174 27674 27226
rect 27854 27174 27856 27226
rect 27610 27172 27616 27174
rect 27672 27172 27696 27174
rect 27752 27172 27776 27174
rect 27832 27172 27856 27174
rect 27912 27172 27918 27174
rect 27610 27163 27918 27172
rect 27610 26140 27918 26149
rect 27610 26138 27616 26140
rect 27672 26138 27696 26140
rect 27752 26138 27776 26140
rect 27832 26138 27856 26140
rect 27912 26138 27918 26140
rect 27672 26086 27674 26138
rect 27854 26086 27856 26138
rect 27610 26084 27616 26086
rect 27672 26084 27696 26086
rect 27752 26084 27776 26086
rect 27832 26084 27856 26086
rect 27912 26084 27918 26086
rect 27610 26075 27918 26084
rect 27610 25052 27918 25061
rect 27610 25050 27616 25052
rect 27672 25050 27696 25052
rect 27752 25050 27776 25052
rect 27832 25050 27856 25052
rect 27912 25050 27918 25052
rect 27672 24998 27674 25050
rect 27854 24998 27856 25050
rect 27610 24996 27616 24998
rect 27672 24996 27696 24998
rect 27752 24996 27776 24998
rect 27832 24996 27856 24998
rect 27912 24996 27918 24998
rect 27610 24987 27918 24996
rect 27528 24948 27580 24954
rect 27528 24890 27580 24896
rect 27448 24818 27568 24834
rect 27436 24812 27568 24818
rect 27488 24806 27568 24812
rect 27436 24754 27488 24760
rect 27540 24698 27568 24806
rect 27620 24744 27672 24750
rect 27264 24670 27476 24698
rect 27344 24608 27396 24614
rect 27344 24550 27396 24556
rect 26950 24508 27258 24517
rect 26950 24506 26956 24508
rect 27012 24506 27036 24508
rect 27092 24506 27116 24508
rect 27172 24506 27196 24508
rect 27252 24506 27258 24508
rect 27012 24454 27014 24506
rect 27194 24454 27196 24506
rect 26950 24452 26956 24454
rect 27012 24452 27036 24454
rect 27092 24452 27116 24454
rect 27172 24452 27196 24454
rect 27252 24452 27258 24454
rect 26950 24443 27258 24452
rect 26950 23420 27258 23429
rect 26950 23418 26956 23420
rect 27012 23418 27036 23420
rect 27092 23418 27116 23420
rect 27172 23418 27196 23420
rect 27252 23418 27258 23420
rect 27012 23366 27014 23418
rect 27194 23366 27196 23418
rect 26950 23364 26956 23366
rect 27012 23364 27036 23366
rect 27092 23364 27116 23366
rect 27172 23364 27196 23366
rect 27252 23364 27258 23366
rect 26950 23355 27258 23364
rect 26950 22332 27258 22341
rect 26950 22330 26956 22332
rect 27012 22330 27036 22332
rect 27092 22330 27116 22332
rect 27172 22330 27196 22332
rect 27252 22330 27258 22332
rect 27012 22278 27014 22330
rect 27194 22278 27196 22330
rect 26950 22276 26956 22278
rect 27012 22276 27036 22278
rect 27092 22276 27116 22278
rect 27172 22276 27196 22278
rect 27252 22276 27258 22278
rect 26950 22267 27258 22276
rect 26950 21244 27258 21253
rect 26950 21242 26956 21244
rect 27012 21242 27036 21244
rect 27092 21242 27116 21244
rect 27172 21242 27196 21244
rect 27252 21242 27258 21244
rect 27012 21190 27014 21242
rect 27194 21190 27196 21242
rect 26950 21188 26956 21190
rect 27012 21188 27036 21190
rect 27092 21188 27116 21190
rect 27172 21188 27196 21190
rect 27252 21188 27258 21190
rect 26950 21179 27258 21188
rect 27356 20874 27384 24550
rect 27448 23186 27476 24670
rect 27540 24692 27620 24698
rect 27540 24686 27672 24692
rect 27540 24670 27660 24686
rect 27540 23662 27568 24670
rect 27610 23964 27918 23973
rect 27610 23962 27616 23964
rect 27672 23962 27696 23964
rect 27752 23962 27776 23964
rect 27832 23962 27856 23964
rect 27912 23962 27918 23964
rect 27672 23910 27674 23962
rect 27854 23910 27856 23962
rect 27610 23908 27616 23910
rect 27672 23908 27696 23910
rect 27752 23908 27776 23910
rect 27832 23908 27856 23910
rect 27912 23908 27918 23910
rect 27610 23899 27918 23908
rect 27528 23656 27580 23662
rect 27528 23598 27580 23604
rect 27436 23180 27488 23186
rect 27436 23122 27488 23128
rect 27610 22876 27918 22885
rect 27610 22874 27616 22876
rect 27672 22874 27696 22876
rect 27752 22874 27776 22876
rect 27832 22874 27856 22876
rect 27912 22874 27918 22876
rect 27672 22822 27674 22874
rect 27854 22822 27856 22874
rect 27610 22820 27616 22822
rect 27672 22820 27696 22822
rect 27752 22820 27776 22822
rect 27832 22820 27856 22822
rect 27912 22820 27918 22822
rect 27610 22811 27918 22820
rect 27610 21788 27918 21797
rect 27610 21786 27616 21788
rect 27672 21786 27696 21788
rect 27752 21786 27776 21788
rect 27832 21786 27856 21788
rect 27912 21786 27918 21788
rect 27672 21734 27674 21786
rect 27854 21734 27856 21786
rect 27610 21732 27616 21734
rect 27672 21732 27696 21734
rect 27752 21732 27776 21734
rect 27832 21732 27856 21734
rect 27912 21732 27918 21734
rect 27610 21723 27918 21732
rect 27344 20868 27396 20874
rect 27344 20810 27396 20816
rect 27356 20466 27384 20810
rect 27610 20700 27918 20709
rect 27610 20698 27616 20700
rect 27672 20698 27696 20700
rect 27752 20698 27776 20700
rect 27832 20698 27856 20700
rect 27912 20698 27918 20700
rect 27672 20646 27674 20698
rect 27854 20646 27856 20698
rect 27610 20644 27616 20646
rect 27672 20644 27696 20646
rect 27752 20644 27776 20646
rect 27832 20644 27856 20646
rect 27912 20644 27918 20646
rect 27610 20635 27918 20644
rect 27344 20460 27396 20466
rect 27344 20402 27396 20408
rect 26950 20156 27258 20165
rect 26950 20154 26956 20156
rect 27012 20154 27036 20156
rect 27092 20154 27116 20156
rect 27172 20154 27196 20156
rect 27252 20154 27258 20156
rect 27012 20102 27014 20154
rect 27194 20102 27196 20154
rect 26950 20100 26956 20102
rect 27012 20100 27036 20102
rect 27092 20100 27116 20102
rect 27172 20100 27196 20102
rect 27252 20100 27258 20102
rect 26950 20091 27258 20100
rect 27344 20052 27396 20058
rect 27344 19994 27396 20000
rect 26950 19068 27258 19077
rect 26950 19066 26956 19068
rect 27012 19066 27036 19068
rect 27092 19066 27116 19068
rect 27172 19066 27196 19068
rect 27252 19066 27258 19068
rect 27012 19014 27014 19066
rect 27194 19014 27196 19066
rect 26950 19012 26956 19014
rect 27012 19012 27036 19014
rect 27092 19012 27116 19014
rect 27172 19012 27196 19014
rect 27252 19012 27258 19014
rect 26950 19003 27258 19012
rect 26950 17980 27258 17989
rect 26950 17978 26956 17980
rect 27012 17978 27036 17980
rect 27092 17978 27116 17980
rect 27172 17978 27196 17980
rect 27252 17978 27258 17980
rect 27012 17926 27014 17978
rect 27194 17926 27196 17978
rect 26950 17924 26956 17926
rect 27012 17924 27036 17926
rect 27092 17924 27116 17926
rect 27172 17924 27196 17926
rect 27252 17924 27258 17926
rect 26950 17915 27258 17924
rect 26950 16892 27258 16901
rect 26950 16890 26956 16892
rect 27012 16890 27036 16892
rect 27092 16890 27116 16892
rect 27172 16890 27196 16892
rect 27252 16890 27258 16892
rect 27012 16838 27014 16890
rect 27194 16838 27196 16890
rect 26950 16836 26956 16838
rect 27012 16836 27036 16838
rect 27092 16836 27116 16838
rect 27172 16836 27196 16838
rect 27252 16836 27258 16838
rect 26950 16827 27258 16836
rect 26950 15804 27258 15813
rect 26950 15802 26956 15804
rect 27012 15802 27036 15804
rect 27092 15802 27116 15804
rect 27172 15802 27196 15804
rect 27252 15802 27258 15804
rect 27012 15750 27014 15802
rect 27194 15750 27196 15802
rect 26950 15748 26956 15750
rect 27012 15748 27036 15750
rect 27092 15748 27116 15750
rect 27172 15748 27196 15750
rect 27252 15748 27258 15750
rect 26950 15739 27258 15748
rect 26950 14716 27258 14725
rect 26950 14714 26956 14716
rect 27012 14714 27036 14716
rect 27092 14714 27116 14716
rect 27172 14714 27196 14716
rect 27252 14714 27258 14716
rect 27012 14662 27014 14714
rect 27194 14662 27196 14714
rect 26950 14660 26956 14662
rect 27012 14660 27036 14662
rect 27092 14660 27116 14662
rect 27172 14660 27196 14662
rect 27252 14660 27258 14662
rect 26950 14651 27258 14660
rect 26950 13628 27258 13637
rect 26950 13626 26956 13628
rect 27012 13626 27036 13628
rect 27092 13626 27116 13628
rect 27172 13626 27196 13628
rect 27252 13626 27258 13628
rect 27012 13574 27014 13626
rect 27194 13574 27196 13626
rect 26950 13572 26956 13574
rect 27012 13572 27036 13574
rect 27092 13572 27116 13574
rect 27172 13572 27196 13574
rect 27252 13572 27258 13574
rect 26950 13563 27258 13572
rect 26950 12540 27258 12549
rect 26950 12538 26956 12540
rect 27012 12538 27036 12540
rect 27092 12538 27116 12540
rect 27172 12538 27196 12540
rect 27252 12538 27258 12540
rect 27012 12486 27014 12538
rect 27194 12486 27196 12538
rect 26950 12484 26956 12486
rect 27012 12484 27036 12486
rect 27092 12484 27116 12486
rect 27172 12484 27196 12486
rect 27252 12484 27258 12486
rect 26950 12475 27258 12484
rect 26950 11452 27258 11461
rect 26950 11450 26956 11452
rect 27012 11450 27036 11452
rect 27092 11450 27116 11452
rect 27172 11450 27196 11452
rect 27252 11450 27258 11452
rect 27012 11398 27014 11450
rect 27194 11398 27196 11450
rect 26950 11396 26956 11398
rect 27012 11396 27036 11398
rect 27092 11396 27116 11398
rect 27172 11396 27196 11398
rect 27252 11396 27258 11398
rect 26950 11387 27258 11396
rect 26950 10364 27258 10373
rect 26950 10362 26956 10364
rect 27012 10362 27036 10364
rect 27092 10362 27116 10364
rect 27172 10362 27196 10364
rect 27252 10362 27258 10364
rect 27012 10310 27014 10362
rect 27194 10310 27196 10362
rect 26950 10308 26956 10310
rect 27012 10308 27036 10310
rect 27092 10308 27116 10310
rect 27172 10308 27196 10310
rect 27252 10308 27258 10310
rect 26950 10299 27258 10308
rect 26950 9276 27258 9285
rect 26950 9274 26956 9276
rect 27012 9274 27036 9276
rect 27092 9274 27116 9276
rect 27172 9274 27196 9276
rect 27252 9274 27258 9276
rect 27012 9222 27014 9274
rect 27194 9222 27196 9274
rect 26950 9220 26956 9222
rect 27012 9220 27036 9222
rect 27092 9220 27116 9222
rect 27172 9220 27196 9222
rect 27252 9220 27258 9222
rect 26950 9211 27258 9220
rect 27356 8974 27384 19994
rect 27610 19612 27918 19621
rect 27610 19610 27616 19612
rect 27672 19610 27696 19612
rect 27752 19610 27776 19612
rect 27832 19610 27856 19612
rect 27912 19610 27918 19612
rect 27672 19558 27674 19610
rect 27854 19558 27856 19610
rect 27610 19556 27616 19558
rect 27672 19556 27696 19558
rect 27752 19556 27776 19558
rect 27832 19556 27856 19558
rect 27912 19556 27918 19558
rect 27610 19547 27918 19556
rect 27610 18524 27918 18533
rect 27610 18522 27616 18524
rect 27672 18522 27696 18524
rect 27752 18522 27776 18524
rect 27832 18522 27856 18524
rect 27912 18522 27918 18524
rect 27672 18470 27674 18522
rect 27854 18470 27856 18522
rect 27610 18468 27616 18470
rect 27672 18468 27696 18470
rect 27752 18468 27776 18470
rect 27832 18468 27856 18470
rect 27912 18468 27918 18470
rect 27610 18459 27918 18468
rect 27610 17436 27918 17445
rect 27610 17434 27616 17436
rect 27672 17434 27696 17436
rect 27752 17434 27776 17436
rect 27832 17434 27856 17436
rect 27912 17434 27918 17436
rect 27672 17382 27674 17434
rect 27854 17382 27856 17434
rect 27610 17380 27616 17382
rect 27672 17380 27696 17382
rect 27752 17380 27776 17382
rect 27832 17380 27856 17382
rect 27912 17380 27918 17382
rect 27610 17371 27918 17380
rect 28460 16522 28488 53382
rect 28736 41414 28764 68750
rect 31116 68672 31168 68678
rect 31116 68614 31168 68620
rect 29644 66632 29696 66638
rect 29644 66574 29696 66580
rect 30104 66632 30156 66638
rect 30104 66574 30156 66580
rect 30288 66632 30340 66638
rect 30288 66574 30340 66580
rect 29368 66496 29420 66502
rect 29368 66438 29420 66444
rect 29000 62416 29052 62422
rect 29000 62358 29052 62364
rect 28908 60104 28960 60110
rect 28908 60046 28960 60052
rect 28920 57866 28948 60046
rect 28908 57860 28960 57866
rect 28908 57802 28960 57808
rect 29012 54194 29040 62358
rect 29092 60512 29144 60518
rect 29092 60454 29144 60460
rect 29104 56234 29132 60454
rect 29092 56228 29144 56234
rect 29092 56170 29144 56176
rect 29000 54188 29052 54194
rect 29000 54130 29052 54136
rect 28816 41472 28868 41478
rect 28816 41414 28868 41420
rect 28552 41386 28764 41414
rect 28552 37398 28580 41386
rect 28724 39568 28776 39574
rect 28724 39510 28776 39516
rect 28632 39364 28684 39370
rect 28632 39306 28684 39312
rect 28644 38962 28672 39306
rect 28736 39098 28764 39510
rect 28724 39092 28776 39098
rect 28724 39034 28776 39040
rect 28632 38956 28684 38962
rect 28632 38898 28684 38904
rect 28540 37392 28592 37398
rect 28540 37334 28592 37340
rect 28644 32434 28672 38898
rect 28632 32428 28684 32434
rect 28632 32370 28684 32376
rect 28644 29714 28672 32370
rect 28736 32366 28764 39034
rect 28828 39030 28856 41414
rect 29184 41200 29236 41206
rect 29184 41142 29236 41148
rect 29196 40934 29224 41142
rect 29276 41132 29328 41138
rect 29276 41074 29328 41080
rect 29288 41002 29316 41074
rect 29276 40996 29328 41002
rect 29276 40938 29328 40944
rect 29184 40928 29236 40934
rect 29184 40870 29236 40876
rect 28966 39086 29224 39114
rect 28966 39030 28994 39086
rect 28816 39024 28868 39030
rect 28816 38966 28868 38972
rect 28954 39024 29006 39030
rect 28954 38966 29006 38972
rect 29090 38992 29146 39001
rect 28828 38758 28856 38966
rect 29196 38962 29224 39086
rect 29090 38927 29092 38936
rect 29144 38927 29146 38936
rect 29184 38956 29236 38962
rect 29092 38898 29144 38904
rect 29184 38898 29236 38904
rect 29012 38826 29224 38842
rect 29000 38820 29236 38826
rect 29052 38814 29184 38820
rect 29000 38762 29052 38768
rect 29184 38762 29236 38768
rect 28816 38752 28868 38758
rect 29092 38752 29144 38758
rect 28816 38694 28868 38700
rect 28998 38720 29054 38729
rect 28828 32434 28856 38694
rect 29054 38700 29092 38706
rect 29054 38694 29144 38700
rect 29054 38678 29132 38694
rect 28998 38655 29054 38664
rect 29012 32434 29040 38655
rect 28816 32428 28868 32434
rect 28816 32370 28868 32376
rect 29000 32428 29052 32434
rect 29000 32370 29052 32376
rect 28724 32360 28776 32366
rect 28724 32302 28776 32308
rect 29288 31754 29316 40938
rect 29380 40594 29408 66438
rect 29552 60716 29604 60722
rect 29552 60658 29604 60664
rect 29460 52624 29512 52630
rect 29460 52566 29512 52572
rect 29368 40588 29420 40594
rect 29368 40530 29420 40536
rect 29472 40390 29500 52566
rect 29564 49706 29592 60658
rect 29656 60178 29684 66574
rect 30116 65686 30144 66574
rect 30104 65680 30156 65686
rect 30104 65622 30156 65628
rect 30196 63844 30248 63850
rect 30196 63786 30248 63792
rect 29736 63368 29788 63374
rect 29736 63310 29788 63316
rect 29644 60172 29696 60178
rect 29644 60114 29696 60120
rect 29552 49700 29604 49706
rect 29552 49642 29604 49648
rect 29564 42158 29592 49642
rect 29552 42152 29604 42158
rect 29552 42094 29604 42100
rect 29748 41682 29776 63310
rect 30208 62422 30236 63786
rect 30300 62966 30328 66574
rect 31024 66088 31076 66094
rect 31024 66030 31076 66036
rect 30564 65748 30616 65754
rect 30564 65690 30616 65696
rect 30472 65476 30524 65482
rect 30472 65418 30524 65424
rect 30288 62960 30340 62966
rect 30288 62902 30340 62908
rect 30196 62416 30248 62422
rect 30196 62358 30248 62364
rect 30300 62354 30328 62902
rect 30288 62348 30340 62354
rect 30288 62290 30340 62296
rect 29920 59016 29972 59022
rect 29920 58958 29972 58964
rect 29932 55214 29960 58958
rect 30012 58880 30064 58886
rect 30012 58822 30064 58828
rect 29840 55186 29960 55214
rect 29840 51074 29868 55186
rect 29920 54664 29972 54670
rect 29920 54606 29972 54612
rect 29932 54330 29960 54606
rect 29920 54324 29972 54330
rect 29920 54266 29972 54272
rect 29840 51046 29960 51074
rect 29828 50516 29880 50522
rect 29828 50458 29880 50464
rect 29736 41676 29788 41682
rect 29736 41618 29788 41624
rect 29644 41268 29696 41274
rect 29644 41210 29696 41216
rect 29460 40384 29512 40390
rect 29460 40326 29512 40332
rect 29366 38992 29422 39001
rect 29366 38927 29422 38936
rect 29380 38894 29408 38927
rect 29368 38888 29420 38894
rect 29368 38830 29420 38836
rect 29472 35630 29500 40326
rect 29552 38888 29604 38894
rect 29552 38830 29604 38836
rect 29564 38729 29592 38830
rect 29550 38720 29606 38729
rect 29550 38655 29606 38664
rect 29552 37664 29604 37670
rect 29552 37606 29604 37612
rect 29460 35624 29512 35630
rect 29460 35566 29512 35572
rect 29104 31726 29316 31754
rect 28632 29708 28684 29714
rect 28632 29650 28684 29656
rect 28448 16516 28500 16522
rect 28448 16458 28500 16464
rect 27610 16348 27918 16357
rect 27610 16346 27616 16348
rect 27672 16346 27696 16348
rect 27752 16346 27776 16348
rect 27832 16346 27856 16348
rect 27912 16346 27918 16348
rect 27672 16294 27674 16346
rect 27854 16294 27856 16346
rect 27610 16292 27616 16294
rect 27672 16292 27696 16294
rect 27752 16292 27776 16294
rect 27832 16292 27856 16294
rect 27912 16292 27918 16294
rect 27610 16283 27918 16292
rect 27610 15260 27918 15269
rect 27610 15258 27616 15260
rect 27672 15258 27696 15260
rect 27752 15258 27776 15260
rect 27832 15258 27856 15260
rect 27912 15258 27918 15260
rect 27672 15206 27674 15258
rect 27854 15206 27856 15258
rect 27610 15204 27616 15206
rect 27672 15204 27696 15206
rect 27752 15204 27776 15206
rect 27832 15204 27856 15206
rect 27912 15204 27918 15206
rect 27610 15195 27918 15204
rect 29104 14550 29132 31726
rect 29564 18290 29592 37606
rect 29656 34950 29684 41210
rect 29736 39568 29788 39574
rect 29736 39510 29788 39516
rect 29748 38962 29776 39510
rect 29736 38956 29788 38962
rect 29736 38898 29788 38904
rect 29644 34944 29696 34950
rect 29644 34886 29696 34892
rect 29656 24138 29684 34886
rect 29644 24132 29696 24138
rect 29644 24074 29696 24080
rect 29644 18420 29696 18426
rect 29644 18362 29696 18368
rect 29552 18284 29604 18290
rect 29552 18226 29604 18232
rect 29656 16574 29684 18362
rect 29564 16546 29684 16574
rect 29092 14544 29144 14550
rect 29092 14486 29144 14492
rect 27610 14172 27918 14181
rect 27610 14170 27616 14172
rect 27672 14170 27696 14172
rect 27752 14170 27776 14172
rect 27832 14170 27856 14172
rect 27912 14170 27918 14172
rect 27672 14118 27674 14170
rect 27854 14118 27856 14170
rect 27610 14116 27616 14118
rect 27672 14116 27696 14118
rect 27752 14116 27776 14118
rect 27832 14116 27856 14118
rect 27912 14116 27918 14118
rect 27610 14107 27918 14116
rect 27610 13084 27918 13093
rect 27610 13082 27616 13084
rect 27672 13082 27696 13084
rect 27752 13082 27776 13084
rect 27832 13082 27856 13084
rect 27912 13082 27918 13084
rect 27672 13030 27674 13082
rect 27854 13030 27856 13082
rect 27610 13028 27616 13030
rect 27672 13028 27696 13030
rect 27752 13028 27776 13030
rect 27832 13028 27856 13030
rect 27912 13028 27918 13030
rect 27610 13019 27918 13028
rect 27610 11996 27918 12005
rect 27610 11994 27616 11996
rect 27672 11994 27696 11996
rect 27752 11994 27776 11996
rect 27832 11994 27856 11996
rect 27912 11994 27918 11996
rect 27672 11942 27674 11994
rect 27854 11942 27856 11994
rect 27610 11940 27616 11942
rect 27672 11940 27696 11942
rect 27752 11940 27776 11942
rect 27832 11940 27856 11942
rect 27912 11940 27918 11942
rect 27610 11931 27918 11940
rect 28172 11008 28224 11014
rect 28172 10950 28224 10956
rect 27610 10908 27918 10917
rect 27610 10906 27616 10908
rect 27672 10906 27696 10908
rect 27752 10906 27776 10908
rect 27832 10906 27856 10908
rect 27912 10906 27918 10908
rect 27672 10854 27674 10906
rect 27854 10854 27856 10906
rect 27610 10852 27616 10854
rect 27672 10852 27696 10854
rect 27752 10852 27776 10854
rect 27832 10852 27856 10854
rect 27912 10852 27918 10854
rect 27610 10843 27918 10852
rect 27610 9820 27918 9829
rect 27610 9818 27616 9820
rect 27672 9818 27696 9820
rect 27752 9818 27776 9820
rect 27832 9818 27856 9820
rect 27912 9818 27918 9820
rect 27672 9766 27674 9818
rect 27854 9766 27856 9818
rect 27610 9764 27616 9766
rect 27672 9764 27696 9766
rect 27752 9764 27776 9766
rect 27832 9764 27856 9766
rect 27912 9764 27918 9766
rect 27610 9755 27918 9764
rect 27344 8968 27396 8974
rect 27344 8910 27396 8916
rect 27528 8968 27580 8974
rect 27528 8910 27580 8916
rect 26950 8188 27258 8197
rect 26950 8186 26956 8188
rect 27012 8186 27036 8188
rect 27092 8186 27116 8188
rect 27172 8186 27196 8188
rect 27252 8186 27258 8188
rect 27012 8134 27014 8186
rect 27194 8134 27196 8186
rect 26950 8132 26956 8134
rect 27012 8132 27036 8134
rect 27092 8132 27116 8134
rect 27172 8132 27196 8134
rect 27252 8132 27258 8134
rect 26950 8123 27258 8132
rect 26792 8084 26844 8090
rect 26792 8026 26844 8032
rect 26950 7100 27258 7109
rect 26950 7098 26956 7100
rect 27012 7098 27036 7100
rect 27092 7098 27116 7100
rect 27172 7098 27196 7100
rect 27252 7098 27258 7100
rect 27012 7046 27014 7098
rect 27194 7046 27196 7098
rect 26950 7044 26956 7046
rect 27012 7044 27036 7046
rect 27092 7044 27116 7046
rect 27172 7044 27196 7046
rect 27252 7044 27258 7046
rect 26950 7035 27258 7044
rect 26950 6012 27258 6021
rect 26950 6010 26956 6012
rect 27012 6010 27036 6012
rect 27092 6010 27116 6012
rect 27172 6010 27196 6012
rect 27252 6010 27258 6012
rect 27012 5958 27014 6010
rect 27194 5958 27196 6010
rect 26950 5956 26956 5958
rect 27012 5956 27036 5958
rect 27092 5956 27116 5958
rect 27172 5956 27196 5958
rect 27252 5956 27258 5958
rect 26950 5947 27258 5956
rect 26950 4924 27258 4933
rect 26950 4922 26956 4924
rect 27012 4922 27036 4924
rect 27092 4922 27116 4924
rect 27172 4922 27196 4924
rect 27252 4922 27258 4924
rect 27012 4870 27014 4922
rect 27194 4870 27196 4922
rect 26950 4868 26956 4870
rect 27012 4868 27036 4870
rect 27092 4868 27116 4870
rect 27172 4868 27196 4870
rect 27252 4868 27258 4870
rect 26950 4859 27258 4868
rect 26424 4684 26476 4690
rect 26424 4626 26476 4632
rect 26950 3836 27258 3845
rect 26950 3834 26956 3836
rect 27012 3834 27036 3836
rect 27092 3834 27116 3836
rect 27172 3834 27196 3836
rect 27252 3834 27258 3836
rect 27012 3782 27014 3834
rect 27194 3782 27196 3834
rect 26950 3780 26956 3782
rect 27012 3780 27036 3782
rect 27092 3780 27116 3782
rect 27172 3780 27196 3782
rect 27252 3780 27258 3782
rect 26950 3771 27258 3780
rect 27540 3194 27568 8910
rect 27610 8732 27918 8741
rect 27610 8730 27616 8732
rect 27672 8730 27696 8732
rect 27752 8730 27776 8732
rect 27832 8730 27856 8732
rect 27912 8730 27918 8732
rect 27672 8678 27674 8730
rect 27854 8678 27856 8730
rect 27610 8676 27616 8678
rect 27672 8676 27696 8678
rect 27752 8676 27776 8678
rect 27832 8676 27856 8678
rect 27912 8676 27918 8678
rect 27610 8667 27918 8676
rect 27610 7644 27918 7653
rect 27610 7642 27616 7644
rect 27672 7642 27696 7644
rect 27752 7642 27776 7644
rect 27832 7642 27856 7644
rect 27912 7642 27918 7644
rect 27672 7590 27674 7642
rect 27854 7590 27856 7642
rect 27610 7588 27616 7590
rect 27672 7588 27696 7590
rect 27752 7588 27776 7590
rect 27832 7588 27856 7590
rect 27912 7588 27918 7590
rect 27610 7579 27918 7588
rect 27610 6556 27918 6565
rect 27610 6554 27616 6556
rect 27672 6554 27696 6556
rect 27752 6554 27776 6556
rect 27832 6554 27856 6556
rect 27912 6554 27918 6556
rect 27672 6502 27674 6554
rect 27854 6502 27856 6554
rect 27610 6500 27616 6502
rect 27672 6500 27696 6502
rect 27752 6500 27776 6502
rect 27832 6500 27856 6502
rect 27912 6500 27918 6502
rect 27610 6491 27918 6500
rect 27610 5468 27918 5477
rect 27610 5466 27616 5468
rect 27672 5466 27696 5468
rect 27752 5466 27776 5468
rect 27832 5466 27856 5468
rect 27912 5466 27918 5468
rect 27672 5414 27674 5466
rect 27854 5414 27856 5466
rect 27610 5412 27616 5414
rect 27672 5412 27696 5414
rect 27752 5412 27776 5414
rect 27832 5412 27856 5414
rect 27912 5412 27918 5414
rect 27610 5403 27918 5412
rect 27610 4380 27918 4389
rect 27610 4378 27616 4380
rect 27672 4378 27696 4380
rect 27752 4378 27776 4380
rect 27832 4378 27856 4380
rect 27912 4378 27918 4380
rect 27672 4326 27674 4378
rect 27854 4326 27856 4378
rect 27610 4324 27616 4326
rect 27672 4324 27696 4326
rect 27752 4324 27776 4326
rect 27832 4324 27856 4326
rect 27912 4324 27918 4326
rect 27610 4315 27918 4324
rect 27610 3292 27918 3301
rect 27610 3290 27616 3292
rect 27672 3290 27696 3292
rect 27752 3290 27776 3292
rect 27832 3290 27856 3292
rect 27912 3290 27918 3292
rect 27672 3238 27674 3290
rect 27854 3238 27856 3290
rect 27610 3236 27616 3238
rect 27672 3236 27696 3238
rect 27752 3236 27776 3238
rect 27832 3236 27856 3238
rect 27912 3236 27918 3238
rect 27610 3227 27918 3236
rect 27528 3188 27580 3194
rect 27528 3130 27580 3136
rect 28184 3058 28212 10950
rect 29564 6186 29592 16546
rect 29840 14346 29868 50458
rect 29932 47598 29960 51046
rect 29920 47592 29972 47598
rect 29920 47534 29972 47540
rect 29932 41274 29960 47534
rect 29920 41268 29972 41274
rect 29920 41210 29972 41216
rect 29920 41132 29972 41138
rect 29920 41074 29972 41080
rect 29932 39302 29960 41074
rect 29920 39296 29972 39302
rect 29920 39238 29972 39244
rect 29932 34678 29960 39238
rect 29920 34672 29972 34678
rect 29920 34614 29972 34620
rect 30024 17270 30052 58822
rect 30104 58676 30156 58682
rect 30104 58618 30156 58624
rect 30116 44946 30144 58618
rect 30288 54596 30340 54602
rect 30288 54538 30340 54544
rect 30104 44940 30156 44946
rect 30104 44882 30156 44888
rect 30104 40928 30156 40934
rect 30104 40870 30156 40876
rect 30116 39098 30144 40870
rect 30196 39432 30248 39438
rect 30196 39374 30248 39380
rect 30104 39092 30156 39098
rect 30104 39034 30156 39040
rect 30208 38758 30236 39374
rect 30196 38752 30248 38758
rect 30196 38694 30248 38700
rect 30104 30116 30156 30122
rect 30104 30058 30156 30064
rect 30116 29102 30144 30058
rect 30104 29096 30156 29102
rect 30104 29038 30156 29044
rect 30104 18284 30156 18290
rect 30104 18226 30156 18232
rect 30012 17264 30064 17270
rect 30012 17206 30064 17212
rect 30116 14550 30144 18226
rect 30104 14544 30156 14550
rect 30104 14486 30156 14492
rect 29828 14340 29880 14346
rect 29828 14282 29880 14288
rect 29644 11756 29696 11762
rect 29644 11698 29696 11704
rect 29656 6730 29684 11698
rect 29644 6724 29696 6730
rect 29644 6666 29696 6672
rect 30208 6662 30236 38694
rect 30300 36310 30328 54538
rect 30380 46504 30432 46510
rect 30380 46446 30432 46452
rect 30392 46034 30420 46446
rect 30380 46028 30432 46034
rect 30380 45970 30432 45976
rect 30484 39030 30512 65418
rect 30576 41138 30604 65690
rect 30656 62280 30708 62286
rect 30656 62222 30708 62228
rect 30668 55214 30696 62222
rect 30932 60104 30984 60110
rect 30932 60046 30984 60052
rect 30668 55186 30788 55214
rect 30564 41132 30616 41138
rect 30564 41074 30616 41080
rect 30576 40089 30604 41074
rect 30562 40080 30618 40089
rect 30562 40015 30618 40024
rect 30564 39908 30616 39914
rect 30564 39850 30616 39856
rect 30576 39030 30604 39850
rect 30760 39642 30788 55186
rect 30840 41132 30892 41138
rect 30840 41074 30892 41080
rect 30748 39636 30800 39642
rect 30748 39578 30800 39584
rect 30748 39432 30800 39438
rect 30748 39374 30800 39380
rect 30472 39024 30524 39030
rect 30472 38966 30524 38972
rect 30564 39024 30616 39030
rect 30564 38966 30616 38972
rect 30760 38962 30788 39374
rect 30748 38956 30800 38962
rect 30748 38898 30800 38904
rect 30472 37732 30524 37738
rect 30472 37674 30524 37680
rect 30380 36780 30432 36786
rect 30380 36722 30432 36728
rect 30288 36304 30340 36310
rect 30288 36246 30340 36252
rect 30392 33046 30420 36722
rect 30484 35698 30512 37674
rect 30748 36304 30800 36310
rect 30748 36246 30800 36252
rect 30472 35692 30524 35698
rect 30472 35634 30524 35640
rect 30484 35494 30512 35634
rect 30472 35488 30524 35494
rect 30472 35430 30524 35436
rect 30380 33040 30432 33046
rect 30380 32982 30432 32988
rect 30484 32586 30512 35430
rect 30484 32558 30604 32586
rect 30472 32428 30524 32434
rect 30472 32370 30524 32376
rect 30484 30190 30512 32370
rect 30576 31890 30604 32558
rect 30564 31884 30616 31890
rect 30564 31826 30616 31832
rect 30380 30184 30432 30190
rect 30380 30126 30432 30132
rect 30472 30184 30524 30190
rect 30472 30126 30524 30132
rect 30392 27402 30420 30126
rect 30380 27396 30432 27402
rect 30380 27338 30432 27344
rect 30392 23050 30420 27338
rect 30380 23044 30432 23050
rect 30380 22986 30432 22992
rect 30760 14414 30788 36246
rect 30852 19718 30880 41074
rect 30944 38962 30972 60046
rect 31036 59090 31064 66030
rect 31128 64870 31156 68614
rect 31116 64864 31168 64870
rect 31116 64806 31168 64812
rect 31496 64530 31524 68750
rect 32610 68572 32918 68581
rect 32610 68570 32616 68572
rect 32672 68570 32696 68572
rect 32752 68570 32776 68572
rect 32832 68570 32856 68572
rect 32912 68570 32918 68572
rect 32672 68518 32674 68570
rect 32854 68518 32856 68570
rect 32610 68516 32616 68518
rect 32672 68516 32696 68518
rect 32752 68516 32776 68518
rect 32832 68516 32856 68518
rect 32912 68516 32918 68518
rect 32610 68507 32918 68516
rect 31950 68028 32258 68037
rect 31950 68026 31956 68028
rect 32012 68026 32036 68028
rect 32092 68026 32116 68028
rect 32172 68026 32196 68028
rect 32252 68026 32258 68028
rect 32012 67974 32014 68026
rect 32194 67974 32196 68026
rect 31950 67972 31956 67974
rect 32012 67972 32036 67974
rect 32092 67972 32116 67974
rect 32172 67972 32196 67974
rect 32252 67972 32258 67974
rect 31950 67963 32258 67972
rect 35348 67924 35400 67930
rect 35348 67866 35400 67872
rect 35256 67720 35308 67726
rect 35256 67662 35308 67668
rect 33140 67652 33192 67658
rect 33140 67594 33192 67600
rect 32610 67484 32918 67493
rect 32610 67482 32616 67484
rect 32672 67482 32696 67484
rect 32752 67482 32776 67484
rect 32832 67482 32856 67484
rect 32912 67482 32918 67484
rect 32672 67430 32674 67482
rect 32854 67430 32856 67482
rect 32610 67428 32616 67430
rect 32672 67428 32696 67430
rect 32752 67428 32776 67430
rect 32832 67428 32856 67430
rect 32912 67428 32918 67430
rect 32610 67419 32918 67428
rect 31950 66940 32258 66949
rect 31950 66938 31956 66940
rect 32012 66938 32036 66940
rect 32092 66938 32116 66940
rect 32172 66938 32196 66940
rect 32252 66938 32258 66940
rect 32012 66886 32014 66938
rect 32194 66886 32196 66938
rect 31950 66884 31956 66886
rect 32012 66884 32036 66886
rect 32092 66884 32116 66886
rect 32172 66884 32196 66886
rect 32252 66884 32258 66886
rect 31950 66875 32258 66884
rect 32610 66396 32918 66405
rect 32610 66394 32616 66396
rect 32672 66394 32696 66396
rect 32752 66394 32776 66396
rect 32832 66394 32856 66396
rect 32912 66394 32918 66396
rect 32672 66342 32674 66394
rect 32854 66342 32856 66394
rect 32610 66340 32616 66342
rect 32672 66340 32696 66342
rect 32752 66340 32776 66342
rect 32832 66340 32856 66342
rect 32912 66340 32918 66342
rect 32610 66331 32918 66340
rect 31950 65852 32258 65861
rect 31950 65850 31956 65852
rect 32012 65850 32036 65852
rect 32092 65850 32116 65852
rect 32172 65850 32196 65852
rect 32252 65850 32258 65852
rect 32012 65798 32014 65850
rect 32194 65798 32196 65850
rect 31950 65796 31956 65798
rect 32012 65796 32036 65798
rect 32092 65796 32116 65798
rect 32172 65796 32196 65798
rect 32252 65796 32258 65798
rect 31950 65787 32258 65796
rect 33152 65754 33180 67594
rect 34704 66564 34756 66570
rect 34704 66506 34756 66512
rect 33140 65748 33192 65754
rect 33140 65690 33192 65696
rect 32610 65308 32918 65317
rect 32610 65306 32616 65308
rect 32672 65306 32696 65308
rect 32752 65306 32776 65308
rect 32832 65306 32856 65308
rect 32912 65306 32918 65308
rect 32672 65254 32674 65306
rect 32854 65254 32856 65306
rect 32610 65252 32616 65254
rect 32672 65252 32696 65254
rect 32752 65252 32776 65254
rect 32832 65252 32856 65254
rect 32912 65252 32918 65254
rect 32610 65243 32918 65252
rect 31950 64764 32258 64773
rect 31950 64762 31956 64764
rect 32012 64762 32036 64764
rect 32092 64762 32116 64764
rect 32172 64762 32196 64764
rect 32252 64762 32258 64764
rect 32012 64710 32014 64762
rect 32194 64710 32196 64762
rect 31950 64708 31956 64710
rect 32012 64708 32036 64710
rect 32092 64708 32116 64710
rect 32172 64708 32196 64710
rect 32252 64708 32258 64710
rect 31950 64699 32258 64708
rect 32404 64592 32456 64598
rect 32404 64534 32456 64540
rect 31484 64524 31536 64530
rect 31484 64466 31536 64472
rect 31024 59084 31076 59090
rect 31024 59026 31076 59032
rect 31496 59022 31524 64466
rect 31950 63676 32258 63685
rect 31950 63674 31956 63676
rect 32012 63674 32036 63676
rect 32092 63674 32116 63676
rect 32172 63674 32196 63676
rect 32252 63674 32258 63676
rect 32012 63622 32014 63674
rect 32194 63622 32196 63674
rect 31950 63620 31956 63622
rect 32012 63620 32036 63622
rect 32092 63620 32116 63622
rect 32172 63620 32196 63622
rect 32252 63620 32258 63622
rect 31950 63611 32258 63620
rect 31950 62588 32258 62597
rect 31950 62586 31956 62588
rect 32012 62586 32036 62588
rect 32092 62586 32116 62588
rect 32172 62586 32196 62588
rect 32252 62586 32258 62588
rect 32012 62534 32014 62586
rect 32194 62534 32196 62586
rect 31950 62532 31956 62534
rect 32012 62532 32036 62534
rect 32092 62532 32116 62534
rect 32172 62532 32196 62534
rect 32252 62532 32258 62534
rect 31950 62523 32258 62532
rect 31950 61500 32258 61509
rect 31950 61498 31956 61500
rect 32012 61498 32036 61500
rect 32092 61498 32116 61500
rect 32172 61498 32196 61500
rect 32252 61498 32258 61500
rect 32012 61446 32014 61498
rect 32194 61446 32196 61498
rect 31950 61444 31956 61446
rect 32012 61444 32036 61446
rect 32092 61444 32116 61446
rect 32172 61444 32196 61446
rect 32252 61444 32258 61446
rect 31950 61435 32258 61444
rect 31950 60412 32258 60421
rect 31950 60410 31956 60412
rect 32012 60410 32036 60412
rect 32092 60410 32116 60412
rect 32172 60410 32196 60412
rect 32252 60410 32258 60412
rect 32012 60358 32014 60410
rect 32194 60358 32196 60410
rect 31950 60356 31956 60358
rect 32012 60356 32036 60358
rect 32092 60356 32116 60358
rect 32172 60356 32196 60358
rect 32252 60356 32258 60358
rect 31950 60347 32258 60356
rect 31950 59324 32258 59333
rect 31950 59322 31956 59324
rect 32012 59322 32036 59324
rect 32092 59322 32116 59324
rect 32172 59322 32196 59324
rect 32252 59322 32258 59324
rect 32012 59270 32014 59322
rect 32194 59270 32196 59322
rect 31950 59268 31956 59270
rect 32012 59268 32036 59270
rect 32092 59268 32116 59270
rect 32172 59268 32196 59270
rect 32252 59268 32258 59270
rect 31950 59259 32258 59268
rect 31484 59016 31536 59022
rect 31484 58958 31536 58964
rect 31950 58236 32258 58245
rect 31950 58234 31956 58236
rect 32012 58234 32036 58236
rect 32092 58234 32116 58236
rect 32172 58234 32196 58236
rect 32252 58234 32258 58236
rect 32012 58182 32014 58234
rect 32194 58182 32196 58234
rect 31950 58180 31956 58182
rect 32012 58180 32036 58182
rect 32092 58180 32116 58182
rect 32172 58180 32196 58182
rect 32252 58180 32258 58182
rect 31950 58171 32258 58180
rect 31668 57588 31720 57594
rect 31668 57530 31720 57536
rect 31208 57316 31260 57322
rect 31208 57258 31260 57264
rect 31300 57316 31352 57322
rect 31300 57258 31352 57264
rect 31116 56908 31168 56914
rect 31116 56850 31168 56856
rect 31024 45892 31076 45898
rect 31024 45834 31076 45840
rect 31036 41070 31064 45834
rect 31128 41478 31156 56850
rect 31116 41472 31168 41478
rect 31116 41414 31168 41420
rect 31024 41064 31076 41070
rect 31024 41006 31076 41012
rect 30932 38956 30984 38962
rect 30932 38898 30984 38904
rect 30944 32502 30972 38898
rect 30932 32496 30984 32502
rect 30932 32438 30984 32444
rect 30932 29776 30984 29782
rect 30932 29718 30984 29724
rect 30944 29170 30972 29718
rect 30932 29164 30984 29170
rect 30932 29106 30984 29112
rect 30932 28076 30984 28082
rect 30932 28018 30984 28024
rect 30840 19712 30892 19718
rect 30840 19654 30892 19660
rect 30944 18698 30972 28018
rect 31036 25838 31064 41006
rect 31220 37194 31248 57258
rect 31312 46986 31340 57258
rect 31576 49768 31628 49774
rect 31576 49710 31628 49716
rect 31300 46980 31352 46986
rect 31300 46922 31352 46928
rect 31300 46028 31352 46034
rect 31300 45970 31352 45976
rect 31208 37188 31260 37194
rect 31208 37130 31260 37136
rect 31116 31816 31168 31822
rect 31116 31758 31168 31764
rect 31128 26234 31156 31758
rect 31220 31142 31248 37130
rect 31208 31136 31260 31142
rect 31208 31078 31260 31084
rect 31208 30116 31260 30122
rect 31208 30058 31260 30064
rect 31220 29646 31248 30058
rect 31208 29640 31260 29646
rect 31208 29582 31260 29588
rect 31128 26206 31248 26234
rect 31024 25832 31076 25838
rect 31024 25774 31076 25780
rect 30932 18692 30984 18698
rect 30932 18634 30984 18640
rect 30748 14408 30800 14414
rect 30748 14350 30800 14356
rect 30288 12776 30340 12782
rect 30288 12718 30340 12724
rect 30300 9042 30328 12718
rect 30288 9036 30340 9042
rect 30288 8978 30340 8984
rect 30944 8022 30972 18634
rect 31024 15972 31076 15978
rect 31024 15914 31076 15920
rect 31036 15094 31064 15914
rect 31220 15094 31248 26206
rect 31024 15088 31076 15094
rect 31024 15030 31076 15036
rect 31208 15088 31260 15094
rect 31208 15030 31260 15036
rect 31220 14346 31248 15030
rect 31312 14414 31340 45970
rect 31484 33040 31536 33046
rect 31484 32982 31536 32988
rect 31392 31136 31444 31142
rect 31392 31078 31444 31084
rect 31404 15026 31432 31078
rect 31496 25226 31524 32982
rect 31588 31346 31616 49710
rect 31576 31340 31628 31346
rect 31576 31282 31628 31288
rect 31680 29238 31708 57530
rect 31950 57148 32258 57157
rect 31950 57146 31956 57148
rect 32012 57146 32036 57148
rect 32092 57146 32116 57148
rect 32172 57146 32196 57148
rect 32252 57146 32258 57148
rect 32012 57094 32014 57146
rect 32194 57094 32196 57146
rect 31950 57092 31956 57094
rect 32012 57092 32036 57094
rect 32092 57092 32116 57094
rect 32172 57092 32196 57094
rect 32252 57092 32258 57094
rect 31950 57083 32258 57092
rect 31950 56060 32258 56069
rect 31950 56058 31956 56060
rect 32012 56058 32036 56060
rect 32092 56058 32116 56060
rect 32172 56058 32196 56060
rect 32252 56058 32258 56060
rect 32012 56006 32014 56058
rect 32194 56006 32196 56058
rect 31950 56004 31956 56006
rect 32012 56004 32036 56006
rect 32092 56004 32116 56006
rect 32172 56004 32196 56006
rect 32252 56004 32258 56006
rect 31950 55995 32258 56004
rect 31950 54972 32258 54981
rect 31950 54970 31956 54972
rect 32012 54970 32036 54972
rect 32092 54970 32116 54972
rect 32172 54970 32196 54972
rect 32252 54970 32258 54972
rect 32012 54918 32014 54970
rect 32194 54918 32196 54970
rect 31950 54916 31956 54918
rect 32012 54916 32036 54918
rect 32092 54916 32116 54918
rect 32172 54916 32196 54918
rect 32252 54916 32258 54918
rect 31950 54907 32258 54916
rect 31950 53884 32258 53893
rect 31950 53882 31956 53884
rect 32012 53882 32036 53884
rect 32092 53882 32116 53884
rect 32172 53882 32196 53884
rect 32252 53882 32258 53884
rect 32012 53830 32014 53882
rect 32194 53830 32196 53882
rect 31950 53828 31956 53830
rect 32012 53828 32036 53830
rect 32092 53828 32116 53830
rect 32172 53828 32196 53830
rect 32252 53828 32258 53830
rect 31950 53819 32258 53828
rect 31950 52796 32258 52805
rect 31950 52794 31956 52796
rect 32012 52794 32036 52796
rect 32092 52794 32116 52796
rect 32172 52794 32196 52796
rect 32252 52794 32258 52796
rect 32012 52742 32014 52794
rect 32194 52742 32196 52794
rect 31950 52740 31956 52742
rect 32012 52740 32036 52742
rect 32092 52740 32116 52742
rect 32172 52740 32196 52742
rect 32252 52740 32258 52742
rect 31950 52731 32258 52740
rect 31950 51708 32258 51717
rect 31950 51706 31956 51708
rect 32012 51706 32036 51708
rect 32092 51706 32116 51708
rect 32172 51706 32196 51708
rect 32252 51706 32258 51708
rect 32012 51654 32014 51706
rect 32194 51654 32196 51706
rect 31950 51652 31956 51654
rect 32012 51652 32036 51654
rect 32092 51652 32116 51654
rect 32172 51652 32196 51654
rect 32252 51652 32258 51654
rect 31950 51643 32258 51652
rect 31760 51400 31812 51406
rect 31760 51342 31812 51348
rect 31772 35834 31800 51342
rect 32416 51066 32444 64534
rect 33692 64456 33744 64462
rect 33692 64398 33744 64404
rect 33600 64388 33652 64394
rect 33600 64330 33652 64336
rect 32610 64220 32918 64229
rect 32610 64218 32616 64220
rect 32672 64218 32696 64220
rect 32752 64218 32776 64220
rect 32832 64218 32856 64220
rect 32912 64218 32918 64220
rect 32672 64166 32674 64218
rect 32854 64166 32856 64218
rect 32610 64164 32616 64166
rect 32672 64164 32696 64166
rect 32752 64164 32776 64166
rect 32832 64164 32856 64166
rect 32912 64164 32918 64166
rect 32610 64155 32918 64164
rect 32610 63132 32918 63141
rect 32610 63130 32616 63132
rect 32672 63130 32696 63132
rect 32752 63130 32776 63132
rect 32832 63130 32856 63132
rect 32912 63130 32918 63132
rect 32672 63078 32674 63130
rect 32854 63078 32856 63130
rect 32610 63076 32616 63078
rect 32672 63076 32696 63078
rect 32752 63076 32776 63078
rect 32832 63076 32856 63078
rect 32912 63076 32918 63078
rect 32610 63067 32918 63076
rect 33612 62801 33640 64330
rect 33598 62792 33654 62801
rect 33598 62727 33654 62736
rect 32610 62044 32918 62053
rect 32610 62042 32616 62044
rect 32672 62042 32696 62044
rect 32752 62042 32776 62044
rect 32832 62042 32856 62044
rect 32912 62042 32918 62044
rect 32672 61990 32674 62042
rect 32854 61990 32856 62042
rect 32610 61988 32616 61990
rect 32672 61988 32696 61990
rect 32752 61988 32776 61990
rect 32832 61988 32856 61990
rect 32912 61988 32918 61990
rect 32610 61979 32918 61988
rect 32610 60956 32918 60965
rect 32610 60954 32616 60956
rect 32672 60954 32696 60956
rect 32752 60954 32776 60956
rect 32832 60954 32856 60956
rect 32912 60954 32918 60956
rect 32672 60902 32674 60954
rect 32854 60902 32856 60954
rect 32610 60900 32616 60902
rect 32672 60900 32696 60902
rect 32752 60900 32776 60902
rect 32832 60900 32856 60902
rect 32912 60900 32918 60902
rect 32610 60891 32918 60900
rect 33140 60104 33192 60110
rect 33140 60046 33192 60052
rect 33416 60104 33468 60110
rect 33416 60046 33468 60052
rect 32610 59868 32918 59877
rect 32610 59866 32616 59868
rect 32672 59866 32696 59868
rect 32752 59866 32776 59868
rect 32832 59866 32856 59868
rect 32912 59866 32918 59868
rect 32672 59814 32674 59866
rect 32854 59814 32856 59866
rect 32610 59812 32616 59814
rect 32672 59812 32696 59814
rect 32752 59812 32776 59814
rect 32832 59812 32856 59814
rect 32912 59812 32918 59814
rect 32610 59803 32918 59812
rect 32610 58780 32918 58789
rect 32610 58778 32616 58780
rect 32672 58778 32696 58780
rect 32752 58778 32776 58780
rect 32832 58778 32856 58780
rect 32912 58778 32918 58780
rect 32672 58726 32674 58778
rect 32854 58726 32856 58778
rect 32610 58724 32616 58726
rect 32672 58724 32696 58726
rect 32752 58724 32776 58726
rect 32832 58724 32856 58726
rect 32912 58724 32918 58726
rect 32610 58715 32918 58724
rect 32610 57692 32918 57701
rect 32610 57690 32616 57692
rect 32672 57690 32696 57692
rect 32752 57690 32776 57692
rect 32832 57690 32856 57692
rect 32912 57690 32918 57692
rect 32672 57638 32674 57690
rect 32854 57638 32856 57690
rect 32610 57636 32616 57638
rect 32672 57636 32696 57638
rect 32752 57636 32776 57638
rect 32832 57636 32856 57638
rect 32912 57636 32918 57638
rect 32610 57627 32918 57636
rect 32610 56604 32918 56613
rect 32610 56602 32616 56604
rect 32672 56602 32696 56604
rect 32752 56602 32776 56604
rect 32832 56602 32856 56604
rect 32912 56602 32918 56604
rect 32672 56550 32674 56602
rect 32854 56550 32856 56602
rect 32610 56548 32616 56550
rect 32672 56548 32696 56550
rect 32752 56548 32776 56550
rect 32832 56548 32856 56550
rect 32912 56548 32918 56550
rect 32610 56539 32918 56548
rect 32610 55516 32918 55525
rect 32610 55514 32616 55516
rect 32672 55514 32696 55516
rect 32752 55514 32776 55516
rect 32832 55514 32856 55516
rect 32912 55514 32918 55516
rect 32672 55462 32674 55514
rect 32854 55462 32856 55514
rect 32610 55460 32616 55462
rect 32672 55460 32696 55462
rect 32752 55460 32776 55462
rect 32832 55460 32856 55462
rect 32912 55460 32918 55462
rect 32610 55451 32918 55460
rect 32610 54428 32918 54437
rect 32610 54426 32616 54428
rect 32672 54426 32696 54428
rect 32752 54426 32776 54428
rect 32832 54426 32856 54428
rect 32912 54426 32918 54428
rect 32672 54374 32674 54426
rect 32854 54374 32856 54426
rect 32610 54372 32616 54374
rect 32672 54372 32696 54374
rect 32752 54372 32776 54374
rect 32832 54372 32856 54374
rect 32912 54372 32918 54374
rect 32610 54363 32918 54372
rect 32610 53340 32918 53349
rect 32610 53338 32616 53340
rect 32672 53338 32696 53340
rect 32752 53338 32776 53340
rect 32832 53338 32856 53340
rect 32912 53338 32918 53340
rect 32672 53286 32674 53338
rect 32854 53286 32856 53338
rect 32610 53284 32616 53286
rect 32672 53284 32696 53286
rect 32752 53284 32776 53286
rect 32832 53284 32856 53286
rect 32912 53284 32918 53286
rect 32610 53275 32918 53284
rect 32610 52252 32918 52261
rect 32610 52250 32616 52252
rect 32672 52250 32696 52252
rect 32752 52250 32776 52252
rect 32832 52250 32856 52252
rect 32912 52250 32918 52252
rect 32672 52198 32674 52250
rect 32854 52198 32856 52250
rect 32610 52196 32616 52198
rect 32672 52196 32696 52198
rect 32752 52196 32776 52198
rect 32832 52196 32856 52198
rect 32912 52196 32918 52198
rect 32610 52187 32918 52196
rect 32610 51164 32918 51173
rect 32610 51162 32616 51164
rect 32672 51162 32696 51164
rect 32752 51162 32776 51164
rect 32832 51162 32856 51164
rect 32912 51162 32918 51164
rect 32672 51110 32674 51162
rect 32854 51110 32856 51162
rect 32610 51108 32616 51110
rect 32672 51108 32696 51110
rect 32752 51108 32776 51110
rect 32832 51108 32856 51110
rect 32912 51108 32918 51110
rect 32610 51099 32918 51108
rect 32404 51060 32456 51066
rect 32404 51002 32456 51008
rect 31950 50620 32258 50629
rect 31950 50618 31956 50620
rect 32012 50618 32036 50620
rect 32092 50618 32116 50620
rect 32172 50618 32196 50620
rect 32252 50618 32258 50620
rect 32012 50566 32014 50618
rect 32194 50566 32196 50618
rect 31950 50564 31956 50566
rect 32012 50564 32036 50566
rect 32092 50564 32116 50566
rect 32172 50564 32196 50566
rect 32252 50564 32258 50566
rect 31950 50555 32258 50564
rect 32610 50076 32918 50085
rect 32610 50074 32616 50076
rect 32672 50074 32696 50076
rect 32752 50074 32776 50076
rect 32832 50074 32856 50076
rect 32912 50074 32918 50076
rect 32672 50022 32674 50074
rect 32854 50022 32856 50074
rect 32610 50020 32616 50022
rect 32672 50020 32696 50022
rect 32752 50020 32776 50022
rect 32832 50020 32856 50022
rect 32912 50020 32918 50022
rect 32610 50011 32918 50020
rect 31950 49532 32258 49541
rect 31950 49530 31956 49532
rect 32012 49530 32036 49532
rect 32092 49530 32116 49532
rect 32172 49530 32196 49532
rect 32252 49530 32258 49532
rect 32012 49478 32014 49530
rect 32194 49478 32196 49530
rect 31950 49476 31956 49478
rect 32012 49476 32036 49478
rect 32092 49476 32116 49478
rect 32172 49476 32196 49478
rect 32252 49476 32258 49478
rect 31950 49467 32258 49476
rect 32610 48988 32918 48997
rect 32610 48986 32616 48988
rect 32672 48986 32696 48988
rect 32752 48986 32776 48988
rect 32832 48986 32856 48988
rect 32912 48986 32918 48988
rect 32672 48934 32674 48986
rect 32854 48934 32856 48986
rect 32610 48932 32616 48934
rect 32672 48932 32696 48934
rect 32752 48932 32776 48934
rect 32832 48932 32856 48934
rect 32912 48932 32918 48934
rect 32610 48923 32918 48932
rect 32956 48748 33008 48754
rect 32956 48690 33008 48696
rect 31950 48444 32258 48453
rect 31950 48442 31956 48444
rect 32012 48442 32036 48444
rect 32092 48442 32116 48444
rect 32172 48442 32196 48444
rect 32252 48442 32258 48444
rect 32012 48390 32014 48442
rect 32194 48390 32196 48442
rect 31950 48388 31956 48390
rect 32012 48388 32036 48390
rect 32092 48388 32116 48390
rect 32172 48388 32196 48390
rect 32252 48388 32258 48390
rect 31950 48379 32258 48388
rect 32610 47900 32918 47909
rect 32610 47898 32616 47900
rect 32672 47898 32696 47900
rect 32752 47898 32776 47900
rect 32832 47898 32856 47900
rect 32912 47898 32918 47900
rect 32672 47846 32674 47898
rect 32854 47846 32856 47898
rect 32610 47844 32616 47846
rect 32672 47844 32696 47846
rect 32752 47844 32776 47846
rect 32832 47844 32856 47846
rect 32912 47844 32918 47846
rect 32610 47835 32918 47844
rect 31950 47356 32258 47365
rect 31950 47354 31956 47356
rect 32012 47354 32036 47356
rect 32092 47354 32116 47356
rect 32172 47354 32196 47356
rect 32252 47354 32258 47356
rect 32012 47302 32014 47354
rect 32194 47302 32196 47354
rect 31950 47300 31956 47302
rect 32012 47300 32036 47302
rect 32092 47300 32116 47302
rect 32172 47300 32196 47302
rect 32252 47300 32258 47302
rect 31950 47291 32258 47300
rect 32610 46812 32918 46821
rect 32610 46810 32616 46812
rect 32672 46810 32696 46812
rect 32752 46810 32776 46812
rect 32832 46810 32856 46812
rect 32912 46810 32918 46812
rect 32672 46758 32674 46810
rect 32854 46758 32856 46810
rect 32610 46756 32616 46758
rect 32672 46756 32696 46758
rect 32752 46756 32776 46758
rect 32832 46756 32856 46758
rect 32912 46756 32918 46758
rect 32610 46747 32918 46756
rect 31950 46268 32258 46277
rect 31950 46266 31956 46268
rect 32012 46266 32036 46268
rect 32092 46266 32116 46268
rect 32172 46266 32196 46268
rect 32252 46266 32258 46268
rect 32012 46214 32014 46266
rect 32194 46214 32196 46266
rect 31950 46212 31956 46214
rect 32012 46212 32036 46214
rect 32092 46212 32116 46214
rect 32172 46212 32196 46214
rect 32252 46212 32258 46214
rect 31950 46203 32258 46212
rect 32610 45724 32918 45733
rect 32610 45722 32616 45724
rect 32672 45722 32696 45724
rect 32752 45722 32776 45724
rect 32832 45722 32856 45724
rect 32912 45722 32918 45724
rect 32672 45670 32674 45722
rect 32854 45670 32856 45722
rect 32610 45668 32616 45670
rect 32672 45668 32696 45670
rect 32752 45668 32776 45670
rect 32832 45668 32856 45670
rect 32912 45668 32918 45670
rect 32610 45659 32918 45668
rect 31950 45180 32258 45189
rect 31950 45178 31956 45180
rect 32012 45178 32036 45180
rect 32092 45178 32116 45180
rect 32172 45178 32196 45180
rect 32252 45178 32258 45180
rect 32012 45126 32014 45178
rect 32194 45126 32196 45178
rect 31950 45124 31956 45126
rect 32012 45124 32036 45126
rect 32092 45124 32116 45126
rect 32172 45124 32196 45126
rect 32252 45124 32258 45126
rect 31950 45115 32258 45124
rect 32404 44940 32456 44946
rect 32404 44882 32456 44888
rect 31852 44804 31904 44810
rect 31852 44746 31904 44752
rect 31864 40526 31892 44746
rect 32312 44736 32364 44742
rect 32312 44678 32364 44684
rect 31950 44092 32258 44101
rect 31950 44090 31956 44092
rect 32012 44090 32036 44092
rect 32092 44090 32116 44092
rect 32172 44090 32196 44092
rect 32252 44090 32258 44092
rect 32012 44038 32014 44090
rect 32194 44038 32196 44090
rect 31950 44036 31956 44038
rect 32012 44036 32036 44038
rect 32092 44036 32116 44038
rect 32172 44036 32196 44038
rect 32252 44036 32258 44038
rect 31950 44027 32258 44036
rect 31950 43004 32258 43013
rect 31950 43002 31956 43004
rect 32012 43002 32036 43004
rect 32092 43002 32116 43004
rect 32172 43002 32196 43004
rect 32252 43002 32258 43004
rect 32012 42950 32014 43002
rect 32194 42950 32196 43002
rect 31950 42948 31956 42950
rect 32012 42948 32036 42950
rect 32092 42948 32116 42950
rect 32172 42948 32196 42950
rect 32252 42948 32258 42950
rect 31950 42939 32258 42948
rect 31950 41916 32258 41925
rect 31950 41914 31956 41916
rect 32012 41914 32036 41916
rect 32092 41914 32116 41916
rect 32172 41914 32196 41916
rect 32252 41914 32258 41916
rect 32012 41862 32014 41914
rect 32194 41862 32196 41914
rect 31950 41860 31956 41862
rect 32012 41860 32036 41862
rect 32092 41860 32116 41862
rect 32172 41860 32196 41862
rect 32252 41860 32258 41862
rect 31950 41851 32258 41860
rect 32324 41546 32352 44678
rect 32312 41540 32364 41546
rect 32312 41482 32364 41488
rect 31950 40828 32258 40837
rect 31950 40826 31956 40828
rect 32012 40826 32036 40828
rect 32092 40826 32116 40828
rect 32172 40826 32196 40828
rect 32252 40826 32258 40828
rect 32012 40774 32014 40826
rect 32194 40774 32196 40826
rect 31950 40772 31956 40774
rect 32012 40772 32036 40774
rect 32092 40772 32116 40774
rect 32172 40772 32196 40774
rect 32252 40772 32258 40774
rect 31950 40763 32258 40772
rect 32416 40526 32444 44882
rect 32588 44872 32640 44878
rect 32508 44820 32588 44826
rect 32508 44814 32640 44820
rect 32508 44798 32628 44814
rect 32508 43994 32536 44798
rect 32610 44636 32918 44645
rect 32610 44634 32616 44636
rect 32672 44634 32696 44636
rect 32752 44634 32776 44636
rect 32832 44634 32856 44636
rect 32912 44634 32918 44636
rect 32672 44582 32674 44634
rect 32854 44582 32856 44634
rect 32610 44580 32616 44582
rect 32672 44580 32696 44582
rect 32752 44580 32776 44582
rect 32832 44580 32856 44582
rect 32912 44580 32918 44582
rect 32610 44571 32918 44580
rect 32496 43988 32548 43994
rect 32496 43930 32548 43936
rect 31852 40520 31904 40526
rect 31852 40462 31904 40468
rect 32404 40520 32456 40526
rect 32404 40462 32456 40468
rect 32312 40044 32364 40050
rect 32312 39986 32364 39992
rect 31950 39740 32258 39749
rect 31950 39738 31956 39740
rect 32012 39738 32036 39740
rect 32092 39738 32116 39740
rect 32172 39738 32196 39740
rect 32252 39738 32258 39740
rect 32012 39686 32014 39738
rect 32194 39686 32196 39738
rect 31950 39684 31956 39686
rect 32012 39684 32036 39686
rect 32092 39684 32116 39686
rect 32172 39684 32196 39686
rect 32252 39684 32258 39686
rect 31950 39675 32258 39684
rect 31852 39296 31904 39302
rect 31852 39238 31904 39244
rect 31760 35828 31812 35834
rect 31760 35770 31812 35776
rect 31864 35766 31892 39238
rect 32324 38758 32352 39986
rect 32312 38752 32364 38758
rect 32312 38694 32364 38700
rect 31950 38652 32258 38661
rect 31950 38650 31956 38652
rect 32012 38650 32036 38652
rect 32092 38650 32116 38652
rect 32172 38650 32196 38652
rect 32252 38650 32258 38652
rect 32012 38598 32014 38650
rect 32194 38598 32196 38650
rect 31950 38596 31956 38598
rect 32012 38596 32036 38598
rect 32092 38596 32116 38598
rect 32172 38596 32196 38598
rect 32252 38596 32258 38598
rect 31950 38587 32258 38596
rect 32312 38548 32364 38554
rect 32312 38490 32364 38496
rect 31950 37564 32258 37573
rect 31950 37562 31956 37564
rect 32012 37562 32036 37564
rect 32092 37562 32116 37564
rect 32172 37562 32196 37564
rect 32252 37562 32258 37564
rect 32012 37510 32014 37562
rect 32194 37510 32196 37562
rect 31950 37508 31956 37510
rect 32012 37508 32036 37510
rect 32092 37508 32116 37510
rect 32172 37508 32196 37510
rect 32252 37508 32258 37510
rect 31950 37499 32258 37508
rect 31950 36476 32258 36485
rect 31950 36474 31956 36476
rect 32012 36474 32036 36476
rect 32092 36474 32116 36476
rect 32172 36474 32196 36476
rect 32252 36474 32258 36476
rect 32012 36422 32014 36474
rect 32194 36422 32196 36474
rect 31950 36420 31956 36422
rect 32012 36420 32036 36422
rect 32092 36420 32116 36422
rect 32172 36420 32196 36422
rect 32252 36420 32258 36422
rect 31950 36411 32258 36420
rect 31852 35760 31904 35766
rect 31852 35702 31904 35708
rect 31950 35388 32258 35397
rect 31950 35386 31956 35388
rect 32012 35386 32036 35388
rect 32092 35386 32116 35388
rect 32172 35386 32196 35388
rect 32252 35386 32258 35388
rect 32012 35334 32014 35386
rect 32194 35334 32196 35386
rect 31950 35332 31956 35334
rect 32012 35332 32036 35334
rect 32092 35332 32116 35334
rect 32172 35332 32196 35334
rect 32252 35332 32258 35334
rect 31950 35323 32258 35332
rect 31950 34300 32258 34309
rect 31950 34298 31956 34300
rect 32012 34298 32036 34300
rect 32092 34298 32116 34300
rect 32172 34298 32196 34300
rect 32252 34298 32258 34300
rect 32012 34246 32014 34298
rect 32194 34246 32196 34298
rect 31950 34244 31956 34246
rect 32012 34244 32036 34246
rect 32092 34244 32116 34246
rect 32172 34244 32196 34246
rect 32252 34244 32258 34246
rect 31950 34235 32258 34244
rect 31950 33212 32258 33221
rect 31950 33210 31956 33212
rect 32012 33210 32036 33212
rect 32092 33210 32116 33212
rect 32172 33210 32196 33212
rect 32252 33210 32258 33212
rect 32012 33158 32014 33210
rect 32194 33158 32196 33210
rect 31950 33156 31956 33158
rect 32012 33156 32036 33158
rect 32092 33156 32116 33158
rect 32172 33156 32196 33158
rect 32252 33156 32258 33158
rect 31950 33147 32258 33156
rect 31950 32124 32258 32133
rect 31950 32122 31956 32124
rect 32012 32122 32036 32124
rect 32092 32122 32116 32124
rect 32172 32122 32196 32124
rect 32252 32122 32258 32124
rect 32012 32070 32014 32122
rect 32194 32070 32196 32122
rect 31950 32068 31956 32070
rect 32012 32068 32036 32070
rect 32092 32068 32116 32070
rect 32172 32068 32196 32070
rect 32252 32068 32258 32070
rect 31950 32059 32258 32068
rect 31950 31036 32258 31045
rect 31950 31034 31956 31036
rect 32012 31034 32036 31036
rect 32092 31034 32116 31036
rect 32172 31034 32196 31036
rect 32252 31034 32258 31036
rect 32012 30982 32014 31034
rect 32194 30982 32196 31034
rect 31950 30980 31956 30982
rect 32012 30980 32036 30982
rect 32092 30980 32116 30982
rect 32172 30980 32196 30982
rect 32252 30980 32258 30982
rect 31950 30971 32258 30980
rect 31950 29948 32258 29957
rect 31950 29946 31956 29948
rect 32012 29946 32036 29948
rect 32092 29946 32116 29948
rect 32172 29946 32196 29948
rect 32252 29946 32258 29948
rect 32012 29894 32014 29946
rect 32194 29894 32196 29946
rect 31950 29892 31956 29894
rect 32012 29892 32036 29894
rect 32092 29892 32116 29894
rect 32172 29892 32196 29894
rect 32252 29892 32258 29894
rect 31950 29883 32258 29892
rect 31944 29504 31996 29510
rect 31944 29446 31996 29452
rect 31668 29232 31720 29238
rect 31668 29174 31720 29180
rect 31484 25220 31536 25226
rect 31484 25162 31536 25168
rect 31392 15020 31444 15026
rect 31392 14962 31444 14968
rect 31496 14890 31524 25162
rect 31484 14884 31536 14890
rect 31484 14826 31536 14832
rect 31300 14408 31352 14414
rect 31300 14350 31352 14356
rect 31208 14340 31260 14346
rect 31208 14282 31260 14288
rect 31208 10464 31260 10470
rect 31208 10406 31260 10412
rect 30932 8016 30984 8022
rect 30932 7958 30984 7964
rect 30196 6656 30248 6662
rect 30196 6598 30248 6604
rect 31220 6322 31248 10406
rect 31680 6322 31708 29174
rect 31956 29050 31984 29446
rect 31864 29022 31984 29050
rect 31760 26376 31812 26382
rect 31760 26318 31812 26324
rect 31772 26246 31800 26318
rect 31760 26240 31812 26246
rect 31760 26182 31812 26188
rect 31760 21480 31812 21486
rect 31760 21422 31812 21428
rect 31772 14890 31800 21422
rect 31760 14884 31812 14890
rect 31760 14826 31812 14832
rect 31772 12170 31800 14826
rect 31760 12164 31812 12170
rect 31760 12106 31812 12112
rect 31864 6322 31892 29022
rect 31950 28860 32258 28869
rect 31950 28858 31956 28860
rect 32012 28858 32036 28860
rect 32092 28858 32116 28860
rect 32172 28858 32196 28860
rect 32252 28858 32258 28860
rect 32012 28806 32014 28858
rect 32194 28806 32196 28858
rect 31950 28804 31956 28806
rect 32012 28804 32036 28806
rect 32092 28804 32116 28806
rect 32172 28804 32196 28806
rect 32252 28804 32258 28806
rect 31950 28795 32258 28804
rect 31950 27772 32258 27781
rect 31950 27770 31956 27772
rect 32012 27770 32036 27772
rect 32092 27770 32116 27772
rect 32172 27770 32196 27772
rect 32252 27770 32258 27772
rect 32012 27718 32014 27770
rect 32194 27718 32196 27770
rect 31950 27716 31956 27718
rect 32012 27716 32036 27718
rect 32092 27716 32116 27718
rect 32172 27716 32196 27718
rect 32252 27716 32258 27718
rect 31950 27707 32258 27716
rect 31950 26684 32258 26693
rect 31950 26682 31956 26684
rect 32012 26682 32036 26684
rect 32092 26682 32116 26684
rect 32172 26682 32196 26684
rect 32252 26682 32258 26684
rect 32012 26630 32014 26682
rect 32194 26630 32196 26682
rect 31950 26628 31956 26630
rect 32012 26628 32036 26630
rect 32092 26628 32116 26630
rect 32172 26628 32196 26630
rect 32252 26628 32258 26630
rect 31950 26619 32258 26628
rect 31950 25596 32258 25605
rect 31950 25594 31956 25596
rect 32012 25594 32036 25596
rect 32092 25594 32116 25596
rect 32172 25594 32196 25596
rect 32252 25594 32258 25596
rect 32012 25542 32014 25594
rect 32194 25542 32196 25594
rect 31950 25540 31956 25542
rect 32012 25540 32036 25542
rect 32092 25540 32116 25542
rect 32172 25540 32196 25542
rect 32252 25540 32258 25542
rect 31950 25531 32258 25540
rect 31950 24508 32258 24517
rect 31950 24506 31956 24508
rect 32012 24506 32036 24508
rect 32092 24506 32116 24508
rect 32172 24506 32196 24508
rect 32252 24506 32258 24508
rect 32012 24454 32014 24506
rect 32194 24454 32196 24506
rect 31950 24452 31956 24454
rect 32012 24452 32036 24454
rect 32092 24452 32116 24454
rect 32172 24452 32196 24454
rect 32252 24452 32258 24454
rect 31950 24443 32258 24452
rect 31950 23420 32258 23429
rect 31950 23418 31956 23420
rect 32012 23418 32036 23420
rect 32092 23418 32116 23420
rect 32172 23418 32196 23420
rect 32252 23418 32258 23420
rect 32012 23366 32014 23418
rect 32194 23366 32196 23418
rect 31950 23364 31956 23366
rect 32012 23364 32036 23366
rect 32092 23364 32116 23366
rect 32172 23364 32196 23366
rect 32252 23364 32258 23366
rect 31950 23355 32258 23364
rect 31950 22332 32258 22341
rect 31950 22330 31956 22332
rect 32012 22330 32036 22332
rect 32092 22330 32116 22332
rect 32172 22330 32196 22332
rect 32252 22330 32258 22332
rect 32012 22278 32014 22330
rect 32194 22278 32196 22330
rect 31950 22276 31956 22278
rect 32012 22276 32036 22278
rect 32092 22276 32116 22278
rect 32172 22276 32196 22278
rect 32252 22276 32258 22278
rect 31950 22267 32258 22276
rect 31950 21244 32258 21253
rect 31950 21242 31956 21244
rect 32012 21242 32036 21244
rect 32092 21242 32116 21244
rect 32172 21242 32196 21244
rect 32252 21242 32258 21244
rect 32012 21190 32014 21242
rect 32194 21190 32196 21242
rect 31950 21188 31956 21190
rect 32012 21188 32036 21190
rect 32092 21188 32116 21190
rect 32172 21188 32196 21190
rect 32252 21188 32258 21190
rect 31950 21179 32258 21188
rect 31950 20156 32258 20165
rect 31950 20154 31956 20156
rect 32012 20154 32036 20156
rect 32092 20154 32116 20156
rect 32172 20154 32196 20156
rect 32252 20154 32258 20156
rect 32012 20102 32014 20154
rect 32194 20102 32196 20154
rect 31950 20100 31956 20102
rect 32012 20100 32036 20102
rect 32092 20100 32116 20102
rect 32172 20100 32196 20102
rect 32252 20100 32258 20102
rect 31950 20091 32258 20100
rect 31950 19068 32258 19077
rect 31950 19066 31956 19068
rect 32012 19066 32036 19068
rect 32092 19066 32116 19068
rect 32172 19066 32196 19068
rect 32252 19066 32258 19068
rect 32012 19014 32014 19066
rect 32194 19014 32196 19066
rect 31950 19012 31956 19014
rect 32012 19012 32036 19014
rect 32092 19012 32116 19014
rect 32172 19012 32196 19014
rect 32252 19012 32258 19014
rect 31950 19003 32258 19012
rect 31950 17980 32258 17989
rect 31950 17978 31956 17980
rect 32012 17978 32036 17980
rect 32092 17978 32116 17980
rect 32172 17978 32196 17980
rect 32252 17978 32258 17980
rect 32012 17926 32014 17978
rect 32194 17926 32196 17978
rect 31950 17924 31956 17926
rect 32012 17924 32036 17926
rect 32092 17924 32116 17926
rect 32172 17924 32196 17926
rect 32252 17924 32258 17926
rect 31950 17915 32258 17924
rect 31950 16892 32258 16901
rect 31950 16890 31956 16892
rect 32012 16890 32036 16892
rect 32092 16890 32116 16892
rect 32172 16890 32196 16892
rect 32252 16890 32258 16892
rect 32012 16838 32014 16890
rect 32194 16838 32196 16890
rect 31950 16836 31956 16838
rect 32012 16836 32036 16838
rect 32092 16836 32116 16838
rect 32172 16836 32196 16838
rect 32252 16836 32258 16838
rect 31950 16827 32258 16836
rect 31950 15804 32258 15813
rect 31950 15802 31956 15804
rect 32012 15802 32036 15804
rect 32092 15802 32116 15804
rect 32172 15802 32196 15804
rect 32252 15802 32258 15804
rect 32012 15750 32014 15802
rect 32194 15750 32196 15802
rect 31950 15748 31956 15750
rect 32012 15748 32036 15750
rect 32092 15748 32116 15750
rect 32172 15748 32196 15750
rect 32252 15748 32258 15750
rect 31950 15739 32258 15748
rect 31950 14716 32258 14725
rect 31950 14714 31956 14716
rect 32012 14714 32036 14716
rect 32092 14714 32116 14716
rect 32172 14714 32196 14716
rect 32252 14714 32258 14716
rect 32012 14662 32014 14714
rect 32194 14662 32196 14714
rect 31950 14660 31956 14662
rect 32012 14660 32036 14662
rect 32092 14660 32116 14662
rect 32172 14660 32196 14662
rect 32252 14660 32258 14662
rect 31950 14651 32258 14660
rect 32324 14550 32352 38490
rect 32416 38010 32444 40462
rect 32508 40066 32536 43930
rect 32610 43548 32918 43557
rect 32610 43546 32616 43548
rect 32672 43546 32696 43548
rect 32752 43546 32776 43548
rect 32832 43546 32856 43548
rect 32912 43546 32918 43548
rect 32672 43494 32674 43546
rect 32854 43494 32856 43546
rect 32610 43492 32616 43494
rect 32672 43492 32696 43494
rect 32752 43492 32776 43494
rect 32832 43492 32856 43494
rect 32912 43492 32918 43494
rect 32610 43483 32918 43492
rect 32610 42460 32918 42469
rect 32610 42458 32616 42460
rect 32672 42458 32696 42460
rect 32752 42458 32776 42460
rect 32832 42458 32856 42460
rect 32912 42458 32918 42460
rect 32672 42406 32674 42458
rect 32854 42406 32856 42458
rect 32610 42404 32616 42406
rect 32672 42404 32696 42406
rect 32752 42404 32776 42406
rect 32832 42404 32856 42406
rect 32912 42404 32918 42406
rect 32610 42395 32918 42404
rect 32968 42242 32996 48690
rect 33048 43444 33100 43450
rect 33048 43386 33100 43392
rect 32784 42214 32996 42242
rect 32784 41614 32812 42214
rect 32864 42152 32916 42158
rect 32864 42094 32916 42100
rect 32772 41608 32824 41614
rect 32772 41550 32824 41556
rect 32876 41562 32904 42094
rect 32876 41534 32996 41562
rect 32610 41372 32918 41381
rect 32610 41370 32616 41372
rect 32672 41370 32696 41372
rect 32752 41370 32776 41372
rect 32832 41370 32856 41372
rect 32912 41370 32918 41372
rect 32672 41318 32674 41370
rect 32854 41318 32856 41370
rect 32610 41316 32616 41318
rect 32672 41316 32696 41318
rect 32752 41316 32776 41318
rect 32832 41316 32856 41318
rect 32912 41316 32918 41318
rect 32610 41307 32918 41316
rect 32610 40284 32918 40293
rect 32610 40282 32616 40284
rect 32672 40282 32696 40284
rect 32752 40282 32776 40284
rect 32832 40282 32856 40284
rect 32912 40282 32918 40284
rect 32672 40230 32674 40282
rect 32854 40230 32856 40282
rect 32610 40228 32616 40230
rect 32672 40228 32696 40230
rect 32752 40228 32776 40230
rect 32832 40228 32856 40230
rect 32912 40228 32918 40230
rect 32610 40219 32918 40228
rect 32508 40038 32628 40066
rect 32600 39284 32628 40038
rect 32968 39370 32996 41534
rect 32956 39364 33008 39370
rect 32956 39306 33008 39312
rect 32508 39256 32628 39284
rect 32404 38004 32456 38010
rect 32404 37946 32456 37952
rect 32508 37856 32536 39256
rect 32610 39196 32918 39205
rect 32610 39194 32616 39196
rect 32672 39194 32696 39196
rect 32752 39194 32776 39196
rect 32832 39194 32856 39196
rect 32912 39194 32918 39196
rect 32672 39142 32674 39194
rect 32854 39142 32856 39194
rect 32610 39140 32616 39142
rect 32672 39140 32696 39142
rect 32752 39140 32776 39142
rect 32832 39140 32856 39142
rect 32912 39140 32918 39142
rect 32610 39131 32918 39140
rect 32968 38434 32996 39306
rect 33060 38554 33088 43386
rect 33152 39574 33180 60046
rect 33428 57594 33456 60046
rect 33416 57588 33468 57594
rect 33416 57530 33468 57536
rect 33508 57248 33560 57254
rect 33508 57190 33560 57196
rect 33232 42220 33284 42226
rect 33232 42162 33284 42168
rect 33244 41682 33272 42162
rect 33232 41676 33284 41682
rect 33232 41618 33284 41624
rect 33140 39568 33192 39574
rect 33140 39510 33192 39516
rect 33140 39432 33192 39438
rect 33140 39374 33192 39380
rect 33152 39098 33180 39374
rect 33140 39092 33192 39098
rect 33140 39034 33192 39040
rect 33048 38548 33100 38554
rect 33048 38490 33100 38496
rect 32968 38406 33088 38434
rect 32610 38108 32918 38117
rect 32610 38106 32616 38108
rect 32672 38106 32696 38108
rect 32752 38106 32776 38108
rect 32832 38106 32856 38108
rect 32912 38106 32918 38108
rect 32672 38054 32674 38106
rect 32854 38054 32856 38106
rect 32610 38052 32616 38054
rect 32672 38052 32696 38054
rect 32752 38052 32776 38054
rect 32832 38052 32856 38054
rect 32912 38052 32918 38054
rect 32610 38043 32918 38052
rect 32416 37828 32536 37856
rect 32312 14544 32364 14550
rect 32312 14486 32364 14492
rect 32416 14482 32444 37828
rect 32588 37800 32640 37806
rect 32588 37742 32640 37748
rect 32496 37392 32548 37398
rect 32600 37380 32628 37742
rect 32548 37352 32628 37380
rect 32496 37334 32548 37340
rect 32508 31822 32536 37334
rect 32610 37020 32918 37029
rect 32610 37018 32616 37020
rect 32672 37018 32696 37020
rect 32752 37018 32776 37020
rect 32832 37018 32856 37020
rect 32912 37018 32918 37020
rect 32672 36966 32674 37018
rect 32854 36966 32856 37018
rect 32610 36964 32616 36966
rect 32672 36964 32696 36966
rect 32752 36964 32776 36966
rect 32832 36964 32856 36966
rect 32912 36964 32918 36966
rect 32610 36955 32918 36964
rect 32610 35932 32918 35941
rect 32610 35930 32616 35932
rect 32672 35930 32696 35932
rect 32752 35930 32776 35932
rect 32832 35930 32856 35932
rect 32912 35930 32918 35932
rect 32672 35878 32674 35930
rect 32854 35878 32856 35930
rect 32610 35876 32616 35878
rect 32672 35876 32696 35878
rect 32752 35876 32776 35878
rect 32832 35876 32856 35878
rect 32912 35876 32918 35878
rect 32610 35867 32918 35876
rect 32610 34844 32918 34853
rect 32610 34842 32616 34844
rect 32672 34842 32696 34844
rect 32752 34842 32776 34844
rect 32832 34842 32856 34844
rect 32912 34842 32918 34844
rect 32672 34790 32674 34842
rect 32854 34790 32856 34842
rect 32610 34788 32616 34790
rect 32672 34788 32696 34790
rect 32752 34788 32776 34790
rect 32832 34788 32856 34790
rect 32912 34788 32918 34790
rect 32610 34779 32918 34788
rect 32610 33756 32918 33765
rect 32610 33754 32616 33756
rect 32672 33754 32696 33756
rect 32752 33754 32776 33756
rect 32832 33754 32856 33756
rect 32912 33754 32918 33756
rect 32672 33702 32674 33754
rect 32854 33702 32856 33754
rect 32610 33700 32616 33702
rect 32672 33700 32696 33702
rect 32752 33700 32776 33702
rect 32832 33700 32856 33702
rect 32912 33700 32918 33702
rect 32610 33691 32918 33700
rect 32610 32668 32918 32677
rect 32610 32666 32616 32668
rect 32672 32666 32696 32668
rect 32752 32666 32776 32668
rect 32832 32666 32856 32668
rect 32912 32666 32918 32668
rect 32672 32614 32674 32666
rect 32854 32614 32856 32666
rect 32610 32612 32616 32614
rect 32672 32612 32696 32614
rect 32752 32612 32776 32614
rect 32832 32612 32856 32614
rect 32912 32612 32918 32614
rect 32610 32603 32918 32612
rect 32496 31816 32548 31822
rect 32496 31758 32548 31764
rect 32610 31580 32918 31589
rect 32610 31578 32616 31580
rect 32672 31578 32696 31580
rect 32752 31578 32776 31580
rect 32832 31578 32856 31580
rect 32912 31578 32918 31580
rect 32672 31526 32674 31578
rect 32854 31526 32856 31578
rect 32610 31524 32616 31526
rect 32672 31524 32696 31526
rect 32752 31524 32776 31526
rect 32832 31524 32856 31526
rect 32912 31524 32918 31526
rect 32610 31515 32918 31524
rect 32610 30492 32918 30501
rect 32610 30490 32616 30492
rect 32672 30490 32696 30492
rect 32752 30490 32776 30492
rect 32832 30490 32856 30492
rect 32912 30490 32918 30492
rect 32672 30438 32674 30490
rect 32854 30438 32856 30490
rect 32610 30436 32616 30438
rect 32672 30436 32696 30438
rect 32752 30436 32776 30438
rect 32832 30436 32856 30438
rect 32912 30436 32918 30438
rect 32610 30427 32918 30436
rect 32496 29572 32548 29578
rect 32496 29514 32548 29520
rect 32508 27470 32536 29514
rect 32610 29404 32918 29413
rect 32610 29402 32616 29404
rect 32672 29402 32696 29404
rect 32752 29402 32776 29404
rect 32832 29402 32856 29404
rect 32912 29402 32918 29404
rect 32672 29350 32674 29402
rect 32854 29350 32856 29402
rect 32610 29348 32616 29350
rect 32672 29348 32696 29350
rect 32752 29348 32776 29350
rect 32832 29348 32856 29350
rect 32912 29348 32918 29350
rect 32610 29339 32918 29348
rect 32610 28316 32918 28325
rect 32610 28314 32616 28316
rect 32672 28314 32696 28316
rect 32752 28314 32776 28316
rect 32832 28314 32856 28316
rect 32912 28314 32918 28316
rect 32672 28262 32674 28314
rect 32854 28262 32856 28314
rect 32610 28260 32616 28262
rect 32672 28260 32696 28262
rect 32752 28260 32776 28262
rect 32832 28260 32856 28262
rect 32912 28260 32918 28262
rect 32610 28251 32918 28260
rect 32956 27872 33008 27878
rect 32956 27814 33008 27820
rect 32496 27464 32548 27470
rect 32496 27406 32548 27412
rect 32610 27228 32918 27237
rect 32610 27226 32616 27228
rect 32672 27226 32696 27228
rect 32752 27226 32776 27228
rect 32832 27226 32856 27228
rect 32912 27226 32918 27228
rect 32672 27174 32674 27226
rect 32854 27174 32856 27226
rect 32610 27172 32616 27174
rect 32672 27172 32696 27174
rect 32752 27172 32776 27174
rect 32832 27172 32856 27174
rect 32912 27172 32918 27174
rect 32610 27163 32918 27172
rect 32610 26140 32918 26149
rect 32610 26138 32616 26140
rect 32672 26138 32696 26140
rect 32752 26138 32776 26140
rect 32832 26138 32856 26140
rect 32912 26138 32918 26140
rect 32672 26086 32674 26138
rect 32854 26086 32856 26138
rect 32610 26084 32616 26086
rect 32672 26084 32696 26086
rect 32752 26084 32776 26086
rect 32832 26084 32856 26086
rect 32912 26084 32918 26086
rect 32610 26075 32918 26084
rect 32610 25052 32918 25061
rect 32610 25050 32616 25052
rect 32672 25050 32696 25052
rect 32752 25050 32776 25052
rect 32832 25050 32856 25052
rect 32912 25050 32918 25052
rect 32672 24998 32674 25050
rect 32854 24998 32856 25050
rect 32610 24996 32616 24998
rect 32672 24996 32696 24998
rect 32752 24996 32776 24998
rect 32832 24996 32856 24998
rect 32912 24996 32918 24998
rect 32610 24987 32918 24996
rect 32610 23964 32918 23973
rect 32610 23962 32616 23964
rect 32672 23962 32696 23964
rect 32752 23962 32776 23964
rect 32832 23962 32856 23964
rect 32912 23962 32918 23964
rect 32672 23910 32674 23962
rect 32854 23910 32856 23962
rect 32610 23908 32616 23910
rect 32672 23908 32696 23910
rect 32752 23908 32776 23910
rect 32832 23908 32856 23910
rect 32912 23908 32918 23910
rect 32610 23899 32918 23908
rect 32610 22876 32918 22885
rect 32610 22874 32616 22876
rect 32672 22874 32696 22876
rect 32752 22874 32776 22876
rect 32832 22874 32856 22876
rect 32912 22874 32918 22876
rect 32672 22822 32674 22874
rect 32854 22822 32856 22874
rect 32610 22820 32616 22822
rect 32672 22820 32696 22822
rect 32752 22820 32776 22822
rect 32832 22820 32856 22822
rect 32912 22820 32918 22822
rect 32610 22811 32918 22820
rect 32968 22574 32996 27814
rect 33060 24206 33088 38406
rect 33140 35216 33192 35222
rect 33140 35158 33192 35164
rect 33152 34542 33180 35158
rect 33140 34536 33192 34542
rect 33140 34478 33192 34484
rect 33244 32910 33272 41618
rect 33324 41472 33376 41478
rect 33324 41414 33376 41420
rect 33232 32904 33284 32910
rect 33232 32846 33284 32852
rect 33232 29028 33284 29034
rect 33232 28970 33284 28976
rect 33048 24200 33100 24206
rect 33048 24142 33100 24148
rect 33060 23662 33088 24142
rect 33048 23656 33100 23662
rect 33048 23598 33100 23604
rect 32956 22568 33008 22574
rect 32956 22510 33008 22516
rect 32610 21788 32918 21797
rect 32610 21786 32616 21788
rect 32672 21786 32696 21788
rect 32752 21786 32776 21788
rect 32832 21786 32856 21788
rect 32912 21786 32918 21788
rect 32672 21734 32674 21786
rect 32854 21734 32856 21786
rect 32610 21732 32616 21734
rect 32672 21732 32696 21734
rect 32752 21732 32776 21734
rect 32832 21732 32856 21734
rect 32912 21732 32918 21734
rect 32610 21723 32918 21732
rect 33244 21350 33272 28970
rect 33232 21344 33284 21350
rect 33232 21286 33284 21292
rect 32610 20700 32918 20709
rect 32610 20698 32616 20700
rect 32672 20698 32696 20700
rect 32752 20698 32776 20700
rect 32832 20698 32856 20700
rect 32912 20698 32918 20700
rect 32672 20646 32674 20698
rect 32854 20646 32856 20698
rect 32610 20644 32616 20646
rect 32672 20644 32696 20646
rect 32752 20644 32776 20646
rect 32832 20644 32856 20646
rect 32912 20644 32918 20646
rect 32610 20635 32918 20644
rect 33140 20256 33192 20262
rect 33140 20198 33192 20204
rect 32610 19612 32918 19621
rect 32610 19610 32616 19612
rect 32672 19610 32696 19612
rect 32752 19610 32776 19612
rect 32832 19610 32856 19612
rect 32912 19610 32918 19612
rect 32672 19558 32674 19610
rect 32854 19558 32856 19610
rect 32610 19556 32616 19558
rect 32672 19556 32696 19558
rect 32752 19556 32776 19558
rect 32832 19556 32856 19558
rect 32912 19556 32918 19558
rect 32610 19547 32918 19556
rect 33152 19514 33180 20198
rect 33232 20052 33284 20058
rect 33232 19994 33284 20000
rect 33244 19854 33272 19994
rect 33336 19854 33364 41414
rect 33416 30252 33468 30258
rect 33416 30194 33468 30200
rect 33428 27538 33456 30194
rect 33416 27532 33468 27538
rect 33416 27474 33468 27480
rect 33416 26920 33468 26926
rect 33416 26862 33468 26868
rect 33428 24206 33456 26862
rect 33416 24200 33468 24206
rect 33416 24142 33468 24148
rect 33232 19848 33284 19854
rect 33232 19790 33284 19796
rect 33324 19848 33376 19854
rect 33324 19790 33376 19796
rect 33232 19712 33284 19718
rect 33232 19654 33284 19660
rect 33140 19508 33192 19514
rect 33140 19450 33192 19456
rect 32610 18524 32918 18533
rect 32610 18522 32616 18524
rect 32672 18522 32696 18524
rect 32752 18522 32776 18524
rect 32832 18522 32856 18524
rect 32912 18522 32918 18524
rect 32672 18470 32674 18522
rect 32854 18470 32856 18522
rect 32610 18468 32616 18470
rect 32672 18468 32696 18470
rect 32752 18468 32776 18470
rect 32832 18468 32856 18470
rect 32912 18468 32918 18470
rect 32610 18459 32918 18468
rect 32610 17436 32918 17445
rect 32610 17434 32616 17436
rect 32672 17434 32696 17436
rect 32752 17434 32776 17436
rect 32832 17434 32856 17436
rect 32912 17434 32918 17436
rect 32672 17382 32674 17434
rect 32854 17382 32856 17434
rect 32610 17380 32616 17382
rect 32672 17380 32696 17382
rect 32752 17380 32776 17382
rect 32832 17380 32856 17382
rect 32912 17380 32918 17382
rect 32610 17371 32918 17380
rect 32610 16348 32918 16357
rect 32610 16346 32616 16348
rect 32672 16346 32696 16348
rect 32752 16346 32776 16348
rect 32832 16346 32856 16348
rect 32912 16346 32918 16348
rect 32672 16294 32674 16346
rect 32854 16294 32856 16346
rect 32610 16292 32616 16294
rect 32672 16292 32696 16294
rect 32752 16292 32776 16294
rect 32832 16292 32856 16294
rect 32912 16292 32918 16294
rect 32610 16283 32918 16292
rect 32610 15260 32918 15269
rect 32610 15258 32616 15260
rect 32672 15258 32696 15260
rect 32752 15258 32776 15260
rect 32832 15258 32856 15260
rect 32912 15258 32918 15260
rect 32672 15206 32674 15258
rect 32854 15206 32856 15258
rect 32610 15204 32616 15206
rect 32672 15204 32696 15206
rect 32752 15204 32776 15206
rect 32832 15204 32856 15206
rect 32912 15204 32918 15206
rect 32610 15195 32918 15204
rect 32404 14476 32456 14482
rect 32404 14418 32456 14424
rect 31950 13628 32258 13637
rect 31950 13626 31956 13628
rect 32012 13626 32036 13628
rect 32092 13626 32116 13628
rect 32172 13626 32196 13628
rect 32252 13626 32258 13628
rect 32012 13574 32014 13626
rect 32194 13574 32196 13626
rect 31950 13572 31956 13574
rect 32012 13572 32036 13574
rect 32092 13572 32116 13574
rect 32172 13572 32196 13574
rect 32252 13572 32258 13574
rect 31950 13563 32258 13572
rect 31950 12540 32258 12549
rect 31950 12538 31956 12540
rect 32012 12538 32036 12540
rect 32092 12538 32116 12540
rect 32172 12538 32196 12540
rect 32252 12538 32258 12540
rect 32012 12486 32014 12538
rect 32194 12486 32196 12538
rect 31950 12484 31956 12486
rect 32012 12484 32036 12486
rect 32092 12484 32116 12486
rect 32172 12484 32196 12486
rect 32252 12484 32258 12486
rect 31950 12475 32258 12484
rect 31950 11452 32258 11461
rect 31950 11450 31956 11452
rect 32012 11450 32036 11452
rect 32092 11450 32116 11452
rect 32172 11450 32196 11452
rect 32252 11450 32258 11452
rect 32012 11398 32014 11450
rect 32194 11398 32196 11450
rect 31950 11396 31956 11398
rect 32012 11396 32036 11398
rect 32092 11396 32116 11398
rect 32172 11396 32196 11398
rect 32252 11396 32258 11398
rect 31950 11387 32258 11396
rect 32416 11150 32444 14418
rect 32610 14172 32918 14181
rect 32610 14170 32616 14172
rect 32672 14170 32696 14172
rect 32752 14170 32776 14172
rect 32832 14170 32856 14172
rect 32912 14170 32918 14172
rect 32672 14118 32674 14170
rect 32854 14118 32856 14170
rect 32610 14116 32616 14118
rect 32672 14116 32696 14118
rect 32752 14116 32776 14118
rect 32832 14116 32856 14118
rect 32912 14116 32918 14118
rect 32610 14107 32918 14116
rect 32610 13084 32918 13093
rect 32610 13082 32616 13084
rect 32672 13082 32696 13084
rect 32752 13082 32776 13084
rect 32832 13082 32856 13084
rect 32912 13082 32918 13084
rect 32672 13030 32674 13082
rect 32854 13030 32856 13082
rect 32610 13028 32616 13030
rect 32672 13028 32696 13030
rect 32752 13028 32776 13030
rect 32832 13028 32856 13030
rect 32912 13028 32918 13030
rect 32610 13019 32918 13028
rect 32610 11996 32918 12005
rect 32610 11994 32616 11996
rect 32672 11994 32696 11996
rect 32752 11994 32776 11996
rect 32832 11994 32856 11996
rect 32912 11994 32918 11996
rect 32672 11942 32674 11994
rect 32854 11942 32856 11994
rect 32610 11940 32616 11942
rect 32672 11940 32696 11942
rect 32752 11940 32776 11942
rect 32832 11940 32856 11942
rect 32912 11940 32918 11942
rect 32610 11931 32918 11940
rect 32404 11144 32456 11150
rect 32404 11086 32456 11092
rect 31950 10364 32258 10373
rect 31950 10362 31956 10364
rect 32012 10362 32036 10364
rect 32092 10362 32116 10364
rect 32172 10362 32196 10364
rect 32252 10362 32258 10364
rect 32012 10310 32014 10362
rect 32194 10310 32196 10362
rect 31950 10308 31956 10310
rect 32012 10308 32036 10310
rect 32092 10308 32116 10310
rect 32172 10308 32196 10310
rect 32252 10308 32258 10310
rect 31950 10299 32258 10308
rect 32416 9654 32444 11086
rect 32610 10908 32918 10917
rect 32610 10906 32616 10908
rect 32672 10906 32696 10908
rect 32752 10906 32776 10908
rect 32832 10906 32856 10908
rect 32912 10906 32918 10908
rect 32672 10854 32674 10906
rect 32854 10854 32856 10906
rect 32610 10852 32616 10854
rect 32672 10852 32696 10854
rect 32752 10852 32776 10854
rect 32832 10852 32856 10854
rect 32912 10852 32918 10854
rect 32610 10843 32918 10852
rect 32610 9820 32918 9829
rect 32610 9818 32616 9820
rect 32672 9818 32696 9820
rect 32752 9818 32776 9820
rect 32832 9818 32856 9820
rect 32912 9818 32918 9820
rect 32672 9766 32674 9818
rect 32854 9766 32856 9818
rect 32610 9764 32616 9766
rect 32672 9764 32696 9766
rect 32752 9764 32776 9766
rect 32832 9764 32856 9766
rect 32912 9764 32918 9766
rect 32610 9755 32918 9764
rect 32404 9648 32456 9654
rect 32404 9590 32456 9596
rect 31950 9276 32258 9285
rect 31950 9274 31956 9276
rect 32012 9274 32036 9276
rect 32092 9274 32116 9276
rect 32172 9274 32196 9276
rect 32252 9274 32258 9276
rect 32012 9222 32014 9274
rect 32194 9222 32196 9274
rect 31950 9220 31956 9222
rect 32012 9220 32036 9222
rect 32092 9220 32116 9222
rect 32172 9220 32196 9222
rect 32252 9220 32258 9222
rect 31950 9211 32258 9220
rect 32610 8732 32918 8741
rect 32610 8730 32616 8732
rect 32672 8730 32696 8732
rect 32752 8730 32776 8732
rect 32832 8730 32856 8732
rect 32912 8730 32918 8732
rect 32672 8678 32674 8730
rect 32854 8678 32856 8730
rect 32610 8676 32616 8678
rect 32672 8676 32696 8678
rect 32752 8676 32776 8678
rect 32832 8676 32856 8678
rect 32912 8676 32918 8678
rect 32610 8667 32918 8676
rect 31950 8188 32258 8197
rect 31950 8186 31956 8188
rect 32012 8186 32036 8188
rect 32092 8186 32116 8188
rect 32172 8186 32196 8188
rect 32252 8186 32258 8188
rect 32012 8134 32014 8186
rect 32194 8134 32196 8186
rect 31950 8132 31956 8134
rect 32012 8132 32036 8134
rect 32092 8132 32116 8134
rect 32172 8132 32196 8134
rect 32252 8132 32258 8134
rect 31950 8123 32258 8132
rect 32610 7644 32918 7653
rect 32610 7642 32616 7644
rect 32672 7642 32696 7644
rect 32752 7642 32776 7644
rect 32832 7642 32856 7644
rect 32912 7642 32918 7644
rect 32672 7590 32674 7642
rect 32854 7590 32856 7642
rect 32610 7588 32616 7590
rect 32672 7588 32696 7590
rect 32752 7588 32776 7590
rect 32832 7588 32856 7590
rect 32912 7588 32918 7590
rect 32610 7579 32918 7588
rect 31950 7100 32258 7109
rect 31950 7098 31956 7100
rect 32012 7098 32036 7100
rect 32092 7098 32116 7100
rect 32172 7098 32196 7100
rect 32252 7098 32258 7100
rect 32012 7046 32014 7098
rect 32194 7046 32196 7098
rect 31950 7044 31956 7046
rect 32012 7044 32036 7046
rect 32092 7044 32116 7046
rect 32172 7044 32196 7046
rect 32252 7044 32258 7046
rect 31950 7035 32258 7044
rect 32610 6556 32918 6565
rect 32610 6554 32616 6556
rect 32672 6554 32696 6556
rect 32752 6554 32776 6556
rect 32832 6554 32856 6556
rect 32912 6554 32918 6556
rect 32672 6502 32674 6554
rect 32854 6502 32856 6554
rect 32610 6500 32616 6502
rect 32672 6500 32696 6502
rect 32752 6500 32776 6502
rect 32832 6500 32856 6502
rect 32912 6500 32918 6502
rect 32610 6491 32918 6500
rect 31208 6316 31260 6322
rect 31208 6258 31260 6264
rect 31668 6316 31720 6322
rect 31668 6258 31720 6264
rect 31852 6316 31904 6322
rect 31852 6258 31904 6264
rect 29552 6180 29604 6186
rect 29552 6122 29604 6128
rect 31950 6012 32258 6021
rect 31950 6010 31956 6012
rect 32012 6010 32036 6012
rect 32092 6010 32116 6012
rect 32172 6010 32196 6012
rect 32252 6010 32258 6012
rect 32012 5958 32014 6010
rect 32194 5958 32196 6010
rect 31950 5956 31956 5958
rect 32012 5956 32036 5958
rect 32092 5956 32116 5958
rect 32172 5956 32196 5958
rect 32252 5956 32258 5958
rect 31950 5947 32258 5956
rect 32610 5468 32918 5477
rect 32610 5466 32616 5468
rect 32672 5466 32696 5468
rect 32752 5466 32776 5468
rect 32832 5466 32856 5468
rect 32912 5466 32918 5468
rect 32672 5414 32674 5466
rect 32854 5414 32856 5466
rect 32610 5412 32616 5414
rect 32672 5412 32696 5414
rect 32752 5412 32776 5414
rect 32832 5412 32856 5414
rect 32912 5412 32918 5414
rect 32610 5403 32918 5412
rect 31024 5024 31076 5030
rect 31024 4966 31076 4972
rect 31036 4826 31064 4966
rect 31950 4924 32258 4933
rect 31950 4922 31956 4924
rect 32012 4922 32036 4924
rect 32092 4922 32116 4924
rect 32172 4922 32196 4924
rect 32252 4922 32258 4924
rect 32012 4870 32014 4922
rect 32194 4870 32196 4922
rect 31950 4868 31956 4870
rect 32012 4868 32036 4870
rect 32092 4868 32116 4870
rect 32172 4868 32196 4870
rect 32252 4868 32258 4870
rect 31950 4859 32258 4868
rect 31024 4820 31076 4826
rect 31024 4762 31076 4768
rect 32610 4380 32918 4389
rect 32610 4378 32616 4380
rect 32672 4378 32696 4380
rect 32752 4378 32776 4380
rect 32832 4378 32856 4380
rect 32912 4378 32918 4380
rect 32672 4326 32674 4378
rect 32854 4326 32856 4378
rect 32610 4324 32616 4326
rect 32672 4324 32696 4326
rect 32752 4324 32776 4326
rect 32832 4324 32856 4326
rect 32912 4324 32918 4326
rect 32610 4315 32918 4324
rect 31950 3836 32258 3845
rect 31950 3834 31956 3836
rect 32012 3834 32036 3836
rect 32092 3834 32116 3836
rect 32172 3834 32196 3836
rect 32252 3834 32258 3836
rect 32012 3782 32014 3834
rect 32194 3782 32196 3834
rect 31950 3780 31956 3782
rect 32012 3780 32036 3782
rect 32092 3780 32116 3782
rect 32172 3780 32196 3782
rect 32252 3780 32258 3782
rect 31950 3771 32258 3780
rect 29644 3392 29696 3398
rect 29644 3334 29696 3340
rect 29656 3126 29684 3334
rect 32610 3292 32918 3301
rect 32610 3290 32616 3292
rect 32672 3290 32696 3292
rect 32752 3290 32776 3292
rect 32832 3290 32856 3292
rect 32912 3290 32918 3292
rect 32672 3238 32674 3290
rect 32854 3238 32856 3290
rect 32610 3236 32616 3238
rect 32672 3236 32696 3238
rect 32752 3236 32776 3238
rect 32832 3236 32856 3238
rect 32912 3236 32918 3238
rect 32610 3227 32918 3236
rect 29644 3120 29696 3126
rect 29644 3062 29696 3068
rect 33244 3058 33272 19654
rect 33428 14414 33456 24142
rect 33520 20058 33548 57190
rect 33704 53106 33732 64398
rect 33876 61192 33928 61198
rect 33876 61134 33928 61140
rect 33784 60104 33836 60110
rect 33784 60046 33836 60052
rect 33692 53100 33744 53106
rect 33692 53042 33744 53048
rect 33796 49842 33824 60046
rect 33784 49836 33836 49842
rect 33784 49778 33836 49784
rect 33784 49700 33836 49706
rect 33784 49642 33836 49648
rect 33600 44464 33652 44470
rect 33600 44406 33652 44412
rect 33508 20052 33560 20058
rect 33508 19994 33560 20000
rect 33416 14408 33468 14414
rect 33416 14350 33468 14356
rect 33428 13870 33456 14350
rect 33416 13864 33468 13870
rect 33416 13806 33468 13812
rect 33612 11150 33640 44406
rect 33692 44192 33744 44198
rect 33692 44134 33744 44140
rect 33704 38350 33732 44134
rect 33692 38344 33744 38350
rect 33692 38286 33744 38292
rect 33704 15026 33732 38286
rect 33796 31278 33824 49642
rect 33784 31272 33836 31278
rect 33784 31214 33836 31220
rect 33784 23588 33836 23594
rect 33784 23530 33836 23536
rect 33796 19718 33824 23530
rect 33784 19712 33836 19718
rect 33784 19654 33836 19660
rect 33888 18086 33916 61134
rect 34716 60314 34744 66506
rect 35268 64054 35296 67662
rect 35256 64048 35308 64054
rect 35256 63990 35308 63996
rect 35268 63578 35296 63990
rect 34796 63572 34848 63578
rect 34796 63514 34848 63520
rect 35256 63572 35308 63578
rect 35256 63514 35308 63520
rect 34704 60308 34756 60314
rect 34704 60250 34756 60256
rect 34152 60104 34204 60110
rect 34152 60046 34204 60052
rect 33968 56160 34020 56166
rect 33968 56102 34020 56108
rect 33980 54534 34008 56102
rect 33968 54528 34020 54534
rect 33968 54470 34020 54476
rect 33980 29034 34008 54470
rect 34060 53100 34112 53106
rect 34060 53042 34112 53048
rect 34072 41206 34100 53042
rect 34164 49706 34192 60046
rect 34704 60036 34756 60042
rect 34704 59978 34756 59984
rect 34716 55894 34744 59978
rect 34704 55888 34756 55894
rect 34704 55830 34756 55836
rect 34704 52420 34756 52426
rect 34704 52362 34756 52368
rect 34716 51105 34744 52362
rect 34702 51096 34758 51105
rect 34702 51031 34758 51040
rect 34152 49700 34204 49706
rect 34152 49642 34204 49648
rect 34060 41200 34112 41206
rect 34060 41142 34112 41148
rect 34704 37256 34756 37262
rect 34704 37198 34756 37204
rect 34152 35216 34204 35222
rect 34152 35158 34204 35164
rect 34060 31816 34112 31822
rect 34060 31758 34112 31764
rect 33968 29028 34020 29034
rect 33968 28970 34020 28976
rect 34072 25430 34100 31758
rect 34060 25424 34112 25430
rect 34060 25366 34112 25372
rect 33876 18080 33928 18086
rect 33876 18022 33928 18028
rect 34072 16574 34100 25366
rect 34164 23662 34192 35158
rect 34244 34672 34296 34678
rect 34244 34614 34296 34620
rect 34256 24206 34284 34614
rect 34520 27668 34572 27674
rect 34520 27610 34572 27616
rect 34244 24200 34296 24206
rect 34244 24142 34296 24148
rect 34256 23730 34284 24142
rect 34244 23724 34296 23730
rect 34244 23666 34296 23672
rect 34152 23656 34204 23662
rect 34152 23598 34204 23604
rect 34336 17876 34388 17882
rect 34336 17818 34388 17824
rect 34072 16546 34284 16574
rect 34256 15026 34284 16546
rect 33692 15020 33744 15026
rect 33692 14962 33744 14968
rect 34244 15020 34296 15026
rect 34244 14962 34296 14968
rect 33600 11144 33652 11150
rect 33600 11086 33652 11092
rect 33704 3670 33732 14962
rect 34256 13394 34284 14962
rect 34348 14958 34376 17818
rect 34336 14952 34388 14958
rect 34336 14894 34388 14900
rect 34244 13388 34296 13394
rect 34244 13330 34296 13336
rect 34532 6866 34560 27610
rect 34612 16652 34664 16658
rect 34612 16594 34664 16600
rect 34624 11150 34652 16594
rect 34716 15502 34744 37198
rect 34704 15496 34756 15502
rect 34704 15438 34756 15444
rect 34612 11144 34664 11150
rect 34612 11086 34664 11092
rect 34612 8356 34664 8362
rect 34612 8298 34664 8304
rect 34520 6860 34572 6866
rect 34520 6802 34572 6808
rect 34152 6248 34204 6254
rect 34152 6190 34204 6196
rect 34164 4146 34192 6190
rect 34152 4140 34204 4146
rect 34152 4082 34204 4088
rect 34164 3738 34192 4082
rect 34152 3732 34204 3738
rect 34152 3674 34204 3680
rect 33692 3664 33744 3670
rect 33692 3606 33744 3612
rect 34164 3194 34192 3674
rect 34152 3188 34204 3194
rect 34152 3130 34204 3136
rect 28172 3052 28224 3058
rect 28172 2994 28224 3000
rect 28632 3052 28684 3058
rect 28632 2994 28684 3000
rect 33232 3052 33284 3058
rect 33232 2994 33284 3000
rect 27988 2984 28040 2990
rect 28644 2938 28672 2994
rect 28040 2932 28672 2938
rect 27988 2926 28672 2932
rect 26332 2916 26384 2922
rect 28000 2910 28672 2926
rect 26332 2858 26384 2864
rect 26950 2748 27258 2757
rect 26950 2746 26956 2748
rect 27012 2746 27036 2748
rect 27092 2746 27116 2748
rect 27172 2746 27196 2748
rect 27252 2746 27258 2748
rect 27012 2694 27014 2746
rect 27194 2694 27196 2746
rect 26950 2692 26956 2694
rect 27012 2692 27036 2694
rect 27092 2692 27116 2694
rect 27172 2692 27196 2694
rect 27252 2692 27258 2694
rect 26950 2683 27258 2692
rect 31950 2748 32258 2757
rect 31950 2746 31956 2748
rect 32012 2746 32036 2748
rect 32092 2746 32116 2748
rect 32172 2746 32196 2748
rect 32252 2746 32258 2748
rect 32012 2694 32014 2746
rect 32194 2694 32196 2746
rect 31950 2692 31956 2694
rect 32012 2692 32036 2694
rect 32092 2692 32116 2694
rect 32172 2692 32196 2694
rect 32252 2692 32258 2694
rect 31950 2683 32258 2692
rect 24584 2644 24636 2650
rect 24584 2586 24636 2592
rect 14372 2576 14424 2582
rect 14372 2518 14424 2524
rect 11704 2508 11756 2514
rect 11704 2450 11756 2456
rect 34164 2446 34192 3130
rect 34624 2514 34652 8298
rect 34808 6914 34836 63514
rect 35256 62280 35308 62286
rect 35256 62222 35308 62228
rect 35268 61713 35296 62222
rect 35254 61704 35310 61713
rect 35254 61639 35310 61648
rect 34888 59968 34940 59974
rect 34888 59910 34940 59916
rect 34900 59702 34928 59910
rect 34888 59696 34940 59702
rect 34888 59638 34940 59644
rect 35164 58948 35216 58954
rect 35164 58890 35216 58896
rect 35176 57050 35204 58890
rect 35164 57044 35216 57050
rect 35164 56986 35216 56992
rect 35176 55214 35204 56986
rect 34992 55186 35204 55214
rect 34888 54732 34940 54738
rect 34888 54674 34940 54680
rect 34900 52358 34928 54674
rect 34992 52358 35020 55186
rect 35072 54800 35124 54806
rect 35072 54742 35124 54748
rect 34888 52352 34940 52358
rect 34888 52294 34940 52300
rect 34980 52352 35032 52358
rect 34980 52294 35032 52300
rect 34900 37262 34928 52294
rect 34980 44328 35032 44334
rect 34980 44270 35032 44276
rect 34992 41614 35020 44270
rect 34980 41608 35032 41614
rect 34980 41550 35032 41556
rect 34888 37256 34940 37262
rect 34888 37198 34940 37204
rect 35084 36174 35112 54742
rect 35256 50448 35308 50454
rect 35256 50390 35308 50396
rect 35268 36174 35296 50390
rect 35072 36168 35124 36174
rect 35072 36110 35124 36116
rect 35256 36168 35308 36174
rect 35256 36110 35308 36116
rect 34980 20460 35032 20466
rect 34980 20402 35032 20408
rect 34992 14958 35020 20402
rect 35072 20392 35124 20398
rect 35072 20334 35124 20340
rect 35084 17610 35112 20334
rect 35164 20256 35216 20262
rect 35164 20198 35216 20204
rect 35072 17604 35124 17610
rect 35072 17546 35124 17552
rect 34980 14952 35032 14958
rect 34980 14894 35032 14900
rect 35084 8974 35112 17546
rect 35176 9178 35204 20198
rect 35360 17882 35388 67866
rect 35452 63306 35480 69294
rect 36950 69116 37258 69125
rect 36950 69114 36956 69116
rect 37012 69114 37036 69116
rect 37092 69114 37116 69116
rect 37172 69114 37196 69116
rect 37252 69114 37258 69116
rect 37012 69062 37014 69114
rect 37194 69062 37196 69114
rect 36950 69060 36956 69062
rect 37012 69060 37036 69062
rect 37092 69060 37116 69062
rect 37172 69060 37196 69062
rect 37252 69060 37258 69062
rect 36950 69051 37258 69060
rect 37610 68572 37918 68581
rect 37610 68570 37616 68572
rect 37672 68570 37696 68572
rect 37752 68570 37776 68572
rect 37832 68570 37856 68572
rect 37912 68570 37918 68572
rect 37672 68518 37674 68570
rect 37854 68518 37856 68570
rect 37610 68516 37616 68518
rect 37672 68516 37696 68518
rect 37752 68516 37776 68518
rect 37832 68516 37856 68518
rect 37912 68516 37918 68518
rect 37610 68507 37918 68516
rect 36950 68028 37258 68037
rect 36950 68026 36956 68028
rect 37012 68026 37036 68028
rect 37092 68026 37116 68028
rect 37172 68026 37196 68028
rect 37252 68026 37258 68028
rect 37012 67974 37014 68026
rect 37194 67974 37196 68026
rect 36950 67972 36956 67974
rect 37012 67972 37036 67974
rect 37092 67972 37116 67974
rect 37172 67972 37196 67974
rect 37252 67972 37258 67974
rect 36950 67963 37258 67972
rect 38016 67856 38068 67862
rect 38014 67824 38016 67833
rect 38068 67824 38070 67833
rect 38014 67759 38070 67768
rect 38108 67788 38160 67794
rect 38108 67730 38160 67736
rect 37096 67720 37148 67726
rect 37094 67688 37096 67697
rect 37148 67688 37150 67697
rect 36360 67652 36412 67658
rect 37094 67623 37150 67632
rect 36360 67594 36412 67600
rect 35992 66088 36044 66094
rect 35992 66030 36044 66036
rect 35440 63300 35492 63306
rect 35440 63242 35492 63248
rect 35452 44334 35480 63242
rect 35624 62280 35676 62286
rect 35624 62222 35676 62228
rect 35440 44328 35492 44334
rect 35440 44270 35492 44276
rect 35532 37936 35584 37942
rect 35532 37878 35584 37884
rect 35544 35894 35572 37878
rect 35452 35866 35572 35894
rect 35452 35018 35480 35866
rect 35440 35012 35492 35018
rect 35440 34954 35492 34960
rect 35452 31754 35480 34954
rect 35452 31726 35572 31754
rect 35440 30320 35492 30326
rect 35440 30262 35492 30268
rect 35452 29850 35480 30262
rect 35440 29844 35492 29850
rect 35440 29786 35492 29792
rect 35452 29646 35480 29786
rect 35440 29640 35492 29646
rect 35440 29582 35492 29588
rect 35452 23798 35480 29582
rect 35440 23792 35492 23798
rect 35440 23734 35492 23740
rect 35348 17876 35400 17882
rect 35348 17818 35400 17824
rect 35256 16516 35308 16522
rect 35256 16458 35308 16464
rect 35268 14958 35296 16458
rect 35544 15434 35572 31726
rect 35636 18426 35664 62222
rect 35808 52488 35860 52494
rect 35808 52430 35860 52436
rect 35820 52154 35848 52430
rect 35808 52148 35860 52154
rect 35808 52090 35860 52096
rect 35808 49836 35860 49842
rect 35808 49778 35860 49784
rect 35820 47734 35848 49778
rect 35808 47728 35860 47734
rect 35808 47670 35860 47676
rect 35900 44260 35952 44266
rect 35900 44202 35952 44208
rect 35716 20528 35768 20534
rect 35716 20470 35768 20476
rect 35624 18420 35676 18426
rect 35624 18362 35676 18368
rect 35532 15428 35584 15434
rect 35532 15370 35584 15376
rect 35346 15056 35402 15065
rect 35346 14991 35348 15000
rect 35400 14991 35402 15000
rect 35348 14962 35400 14968
rect 35256 14952 35308 14958
rect 35256 14894 35308 14900
rect 35544 13258 35572 15370
rect 35728 14278 35756 20470
rect 35716 14272 35768 14278
rect 35716 14214 35768 14220
rect 35532 13252 35584 13258
rect 35532 13194 35584 13200
rect 35164 9172 35216 9178
rect 35164 9114 35216 9120
rect 35072 8968 35124 8974
rect 35072 8910 35124 8916
rect 34716 6886 34836 6914
rect 34716 6730 34744 6886
rect 35532 6792 35584 6798
rect 35532 6734 35584 6740
rect 35624 6792 35676 6798
rect 35624 6734 35676 6740
rect 34704 6724 34756 6730
rect 34704 6666 34756 6672
rect 34716 4622 34744 6666
rect 34704 4616 34756 4622
rect 34704 4558 34756 4564
rect 35544 4486 35572 6734
rect 35636 6662 35664 6734
rect 35624 6656 35676 6662
rect 35624 6598 35676 6604
rect 35636 4826 35664 6598
rect 35624 4820 35676 4826
rect 35624 4762 35676 4768
rect 35532 4480 35584 4486
rect 35532 4422 35584 4428
rect 35912 3602 35940 44202
rect 36004 42090 36032 66030
rect 36372 63986 36400 67594
rect 37610 67484 37918 67493
rect 37610 67482 37616 67484
rect 37672 67482 37696 67484
rect 37752 67482 37776 67484
rect 37832 67482 37856 67484
rect 37912 67482 37918 67484
rect 37672 67430 37674 67482
rect 37854 67430 37856 67482
rect 37610 67428 37616 67430
rect 37672 67428 37696 67430
rect 37752 67428 37776 67430
rect 37832 67428 37856 67430
rect 37912 67428 37918 67430
rect 37610 67419 37918 67428
rect 37280 67312 37332 67318
rect 37280 67254 37332 67260
rect 36950 66940 37258 66949
rect 36950 66938 36956 66940
rect 37012 66938 37036 66940
rect 37092 66938 37116 66940
rect 37172 66938 37196 66940
rect 37252 66938 37258 66940
rect 37012 66886 37014 66938
rect 37194 66886 37196 66938
rect 36950 66884 36956 66886
rect 37012 66884 37036 66886
rect 37092 66884 37116 66886
rect 37172 66884 37196 66886
rect 37252 66884 37258 66886
rect 36950 66875 37258 66884
rect 36950 65852 37258 65861
rect 36950 65850 36956 65852
rect 37012 65850 37036 65852
rect 37092 65850 37116 65852
rect 37172 65850 37196 65852
rect 37252 65850 37258 65852
rect 37012 65798 37014 65850
rect 37194 65798 37196 65850
rect 36950 65796 36956 65798
rect 37012 65796 37036 65798
rect 37092 65796 37116 65798
rect 37172 65796 37196 65798
rect 37252 65796 37258 65798
rect 36950 65787 37258 65796
rect 37292 65618 37320 67254
rect 38016 67244 38068 67250
rect 38016 67186 38068 67192
rect 37610 66396 37918 66405
rect 37610 66394 37616 66396
rect 37672 66394 37696 66396
rect 37752 66394 37776 66396
rect 37832 66394 37856 66396
rect 37912 66394 37918 66396
rect 37672 66342 37674 66394
rect 37854 66342 37856 66394
rect 37610 66340 37616 66342
rect 37672 66340 37696 66342
rect 37752 66340 37776 66342
rect 37832 66340 37856 66342
rect 37912 66340 37918 66342
rect 37610 66331 37918 66340
rect 37280 65612 37332 65618
rect 37280 65554 37332 65560
rect 37610 65308 37918 65317
rect 37610 65306 37616 65308
rect 37672 65306 37696 65308
rect 37752 65306 37776 65308
rect 37832 65306 37856 65308
rect 37912 65306 37918 65308
rect 37672 65254 37674 65306
rect 37854 65254 37856 65306
rect 37610 65252 37616 65254
rect 37672 65252 37696 65254
rect 37752 65252 37776 65254
rect 37832 65252 37856 65254
rect 37912 65252 37918 65254
rect 37610 65243 37918 65252
rect 36950 64764 37258 64773
rect 36950 64762 36956 64764
rect 37012 64762 37036 64764
rect 37092 64762 37116 64764
rect 37172 64762 37196 64764
rect 37252 64762 37258 64764
rect 37012 64710 37014 64762
rect 37194 64710 37196 64762
rect 36950 64708 36956 64710
rect 37012 64708 37036 64710
rect 37092 64708 37116 64710
rect 37172 64708 37196 64710
rect 37252 64708 37258 64710
rect 36950 64699 37258 64708
rect 36728 64456 36780 64462
rect 36728 64398 36780 64404
rect 36360 63980 36412 63986
rect 36360 63922 36412 63928
rect 36268 51944 36320 51950
rect 36268 51886 36320 51892
rect 36084 42152 36136 42158
rect 36084 42094 36136 42100
rect 35992 42084 36044 42090
rect 35992 42026 36044 42032
rect 35992 33108 36044 33114
rect 35992 33050 36044 33056
rect 36004 32842 36032 33050
rect 35992 32836 36044 32842
rect 35992 32778 36044 32784
rect 35992 30932 36044 30938
rect 35992 30874 36044 30880
rect 36004 27878 36032 30874
rect 36096 30682 36124 42094
rect 36280 40594 36308 51886
rect 36268 40588 36320 40594
rect 36268 40530 36320 40536
rect 36176 34536 36228 34542
rect 36176 34478 36228 34484
rect 36188 30818 36216 34478
rect 36372 30938 36400 63922
rect 36544 61396 36596 61402
rect 36544 61338 36596 61344
rect 36452 53168 36504 53174
rect 36452 53110 36504 53116
rect 36464 44266 36492 53110
rect 36556 52494 36584 61338
rect 36740 53174 36768 64398
rect 37610 64220 37918 64229
rect 37610 64218 37616 64220
rect 37672 64218 37696 64220
rect 37752 64218 37776 64220
rect 37832 64218 37856 64220
rect 37912 64218 37918 64220
rect 37672 64166 37674 64218
rect 37854 64166 37856 64218
rect 37610 64164 37616 64166
rect 37672 64164 37696 64166
rect 37752 64164 37776 64166
rect 37832 64164 37856 64166
rect 37912 64164 37918 64166
rect 37610 64155 37918 64164
rect 37372 63912 37424 63918
rect 37372 63854 37424 63860
rect 36950 63676 37258 63685
rect 36950 63674 36956 63676
rect 37012 63674 37036 63676
rect 37092 63674 37116 63676
rect 37172 63674 37196 63676
rect 37252 63674 37258 63676
rect 37012 63622 37014 63674
rect 37194 63622 37196 63674
rect 36950 63620 36956 63622
rect 37012 63620 37036 63622
rect 37092 63620 37116 63622
rect 37172 63620 37196 63622
rect 37252 63620 37258 63622
rect 36950 63611 37258 63620
rect 36950 62588 37258 62597
rect 36950 62586 36956 62588
rect 37012 62586 37036 62588
rect 37092 62586 37116 62588
rect 37172 62586 37196 62588
rect 37252 62586 37258 62588
rect 37012 62534 37014 62586
rect 37194 62534 37196 62586
rect 36950 62532 36956 62534
rect 37012 62532 37036 62534
rect 37092 62532 37116 62534
rect 37172 62532 37196 62534
rect 37252 62532 37258 62534
rect 36950 62523 37258 62532
rect 36950 61500 37258 61509
rect 36950 61498 36956 61500
rect 37012 61498 37036 61500
rect 37092 61498 37116 61500
rect 37172 61498 37196 61500
rect 37252 61498 37258 61500
rect 37012 61446 37014 61498
rect 37194 61446 37196 61498
rect 36950 61444 36956 61446
rect 37012 61444 37036 61446
rect 37092 61444 37116 61446
rect 37172 61444 37196 61446
rect 37252 61444 37258 61446
rect 36950 61435 37258 61444
rect 36950 60412 37258 60421
rect 36950 60410 36956 60412
rect 37012 60410 37036 60412
rect 37092 60410 37116 60412
rect 37172 60410 37196 60412
rect 37252 60410 37258 60412
rect 37012 60358 37014 60410
rect 37194 60358 37196 60410
rect 36950 60356 36956 60358
rect 37012 60356 37036 60358
rect 37092 60356 37116 60358
rect 37172 60356 37196 60358
rect 37252 60356 37258 60358
rect 36950 60347 37258 60356
rect 36950 59324 37258 59333
rect 36950 59322 36956 59324
rect 37012 59322 37036 59324
rect 37092 59322 37116 59324
rect 37172 59322 37196 59324
rect 37252 59322 37258 59324
rect 37012 59270 37014 59322
rect 37194 59270 37196 59322
rect 36950 59268 36956 59270
rect 37012 59268 37036 59270
rect 37092 59268 37116 59270
rect 37172 59268 37196 59270
rect 37252 59268 37258 59270
rect 36950 59259 37258 59268
rect 36950 58236 37258 58245
rect 36950 58234 36956 58236
rect 37012 58234 37036 58236
rect 37092 58234 37116 58236
rect 37172 58234 37196 58236
rect 37252 58234 37258 58236
rect 37012 58182 37014 58234
rect 37194 58182 37196 58234
rect 36950 58180 36956 58182
rect 37012 58180 37036 58182
rect 37092 58180 37116 58182
rect 37172 58180 37196 58182
rect 37252 58180 37258 58182
rect 36950 58171 37258 58180
rect 36950 57148 37258 57157
rect 36950 57146 36956 57148
rect 37012 57146 37036 57148
rect 37092 57146 37116 57148
rect 37172 57146 37196 57148
rect 37252 57146 37258 57148
rect 37012 57094 37014 57146
rect 37194 57094 37196 57146
rect 36950 57092 36956 57094
rect 37012 57092 37036 57094
rect 37092 57092 37116 57094
rect 37172 57092 37196 57094
rect 37252 57092 37258 57094
rect 36950 57083 37258 57092
rect 36950 56060 37258 56069
rect 36950 56058 36956 56060
rect 37012 56058 37036 56060
rect 37092 56058 37116 56060
rect 37172 56058 37196 56060
rect 37252 56058 37258 56060
rect 37012 56006 37014 56058
rect 37194 56006 37196 56058
rect 36950 56004 36956 56006
rect 37012 56004 37036 56006
rect 37092 56004 37116 56006
rect 37172 56004 37196 56006
rect 37252 56004 37258 56006
rect 36950 55995 37258 56004
rect 37384 55214 37412 63854
rect 37610 63132 37918 63141
rect 37610 63130 37616 63132
rect 37672 63130 37696 63132
rect 37752 63130 37776 63132
rect 37832 63130 37856 63132
rect 37912 63130 37918 63132
rect 37672 63078 37674 63130
rect 37854 63078 37856 63130
rect 37610 63076 37616 63078
rect 37672 63076 37696 63078
rect 37752 63076 37776 63078
rect 37832 63076 37856 63078
rect 37912 63076 37918 63078
rect 37610 63067 37918 63076
rect 37610 62044 37918 62053
rect 37610 62042 37616 62044
rect 37672 62042 37696 62044
rect 37752 62042 37776 62044
rect 37832 62042 37856 62044
rect 37912 62042 37918 62044
rect 37672 61990 37674 62042
rect 37854 61990 37856 62042
rect 37610 61988 37616 61990
rect 37672 61988 37696 61990
rect 37752 61988 37776 61990
rect 37832 61988 37856 61990
rect 37912 61988 37918 61990
rect 37610 61979 37918 61988
rect 37610 60956 37918 60965
rect 37610 60954 37616 60956
rect 37672 60954 37696 60956
rect 37752 60954 37776 60956
rect 37832 60954 37856 60956
rect 37912 60954 37918 60956
rect 37672 60902 37674 60954
rect 37854 60902 37856 60954
rect 37610 60900 37616 60902
rect 37672 60900 37696 60902
rect 37752 60900 37776 60902
rect 37832 60900 37856 60902
rect 37912 60900 37918 60902
rect 37610 60891 37918 60900
rect 37610 59868 37918 59877
rect 37610 59866 37616 59868
rect 37672 59866 37696 59868
rect 37752 59866 37776 59868
rect 37832 59866 37856 59868
rect 37912 59866 37918 59868
rect 37672 59814 37674 59866
rect 37854 59814 37856 59866
rect 37610 59812 37616 59814
rect 37672 59812 37696 59814
rect 37752 59812 37776 59814
rect 37832 59812 37856 59814
rect 37912 59812 37918 59814
rect 37610 59803 37918 59812
rect 38028 59090 38056 67186
rect 38120 63986 38148 67730
rect 38384 67652 38436 67658
rect 38384 67594 38436 67600
rect 38292 67244 38344 67250
rect 38292 67186 38344 67192
rect 38304 67114 38332 67186
rect 38292 67108 38344 67114
rect 38292 67050 38344 67056
rect 38108 63980 38160 63986
rect 38108 63922 38160 63928
rect 38016 59084 38068 59090
rect 38016 59026 38068 59032
rect 37610 58780 37918 58789
rect 37610 58778 37616 58780
rect 37672 58778 37696 58780
rect 37752 58778 37776 58780
rect 37832 58778 37856 58780
rect 37912 58778 37918 58780
rect 37672 58726 37674 58778
rect 37854 58726 37856 58778
rect 37610 58724 37616 58726
rect 37672 58724 37696 58726
rect 37752 58724 37776 58726
rect 37832 58724 37856 58726
rect 37912 58724 37918 58726
rect 37610 58715 37918 58724
rect 38016 58472 38068 58478
rect 38016 58414 38068 58420
rect 37610 57692 37918 57701
rect 37610 57690 37616 57692
rect 37672 57690 37696 57692
rect 37752 57690 37776 57692
rect 37832 57690 37856 57692
rect 37912 57690 37918 57692
rect 37672 57638 37674 57690
rect 37854 57638 37856 57690
rect 37610 57636 37616 57638
rect 37672 57636 37696 57638
rect 37752 57636 37776 57638
rect 37832 57636 37856 57638
rect 37912 57636 37918 57638
rect 37610 57627 37918 57636
rect 37610 56604 37918 56613
rect 37610 56602 37616 56604
rect 37672 56602 37696 56604
rect 37752 56602 37776 56604
rect 37832 56602 37856 56604
rect 37912 56602 37918 56604
rect 37672 56550 37674 56602
rect 37854 56550 37856 56602
rect 37610 56548 37616 56550
rect 37672 56548 37696 56550
rect 37752 56548 37776 56550
rect 37832 56548 37856 56550
rect 37912 56548 37918 56550
rect 37610 56539 37918 56548
rect 37610 55516 37918 55525
rect 37610 55514 37616 55516
rect 37672 55514 37696 55516
rect 37752 55514 37776 55516
rect 37832 55514 37856 55516
rect 37912 55514 37918 55516
rect 37672 55462 37674 55514
rect 37854 55462 37856 55514
rect 37610 55460 37616 55462
rect 37672 55460 37696 55462
rect 37752 55460 37776 55462
rect 37832 55460 37856 55462
rect 37912 55460 37918 55462
rect 37610 55451 37918 55460
rect 37292 55186 37412 55214
rect 38028 55214 38056 58414
rect 38028 55186 38148 55214
rect 36950 54972 37258 54981
rect 36950 54970 36956 54972
rect 37012 54970 37036 54972
rect 37092 54970 37116 54972
rect 37172 54970 37196 54972
rect 37252 54970 37258 54972
rect 37012 54918 37014 54970
rect 37194 54918 37196 54970
rect 36950 54916 36956 54918
rect 37012 54916 37036 54918
rect 37092 54916 37116 54918
rect 37172 54916 37196 54918
rect 37252 54916 37258 54918
rect 36950 54907 37258 54916
rect 36950 53884 37258 53893
rect 36950 53882 36956 53884
rect 37012 53882 37036 53884
rect 37092 53882 37116 53884
rect 37172 53882 37196 53884
rect 37252 53882 37258 53884
rect 37012 53830 37014 53882
rect 37194 53830 37196 53882
rect 36950 53828 36956 53830
rect 37012 53828 37036 53830
rect 37092 53828 37116 53830
rect 37172 53828 37196 53830
rect 37252 53828 37258 53830
rect 36950 53819 37258 53828
rect 36728 53168 36780 53174
rect 36728 53110 36780 53116
rect 36728 52896 36780 52902
rect 36728 52838 36780 52844
rect 36544 52488 36596 52494
rect 36544 52430 36596 52436
rect 36452 44260 36504 44266
rect 36452 44202 36504 44208
rect 36556 35630 36584 52430
rect 36636 49836 36688 49842
rect 36636 49778 36688 49784
rect 36648 43654 36676 49778
rect 36740 46374 36768 52838
rect 36950 52796 37258 52805
rect 36950 52794 36956 52796
rect 37012 52794 37036 52796
rect 37092 52794 37116 52796
rect 37172 52794 37196 52796
rect 37252 52794 37258 52796
rect 37012 52742 37014 52794
rect 37194 52742 37196 52794
rect 36950 52740 36956 52742
rect 37012 52740 37036 52742
rect 37092 52740 37116 52742
rect 37172 52740 37196 52742
rect 37252 52740 37258 52742
rect 36950 52731 37258 52740
rect 36820 52692 36872 52698
rect 36820 52634 36872 52640
rect 36832 51406 36860 52634
rect 36950 51708 37258 51717
rect 36950 51706 36956 51708
rect 37012 51706 37036 51708
rect 37092 51706 37116 51708
rect 37172 51706 37196 51708
rect 37252 51706 37258 51708
rect 37012 51654 37014 51706
rect 37194 51654 37196 51706
rect 36950 51652 36956 51654
rect 37012 51652 37036 51654
rect 37092 51652 37116 51654
rect 37172 51652 37196 51654
rect 37252 51652 37258 51654
rect 36950 51643 37258 51652
rect 36820 51400 36872 51406
rect 36820 51342 36872 51348
rect 36950 50620 37258 50629
rect 36950 50618 36956 50620
rect 37012 50618 37036 50620
rect 37092 50618 37116 50620
rect 37172 50618 37196 50620
rect 37252 50618 37258 50620
rect 37012 50566 37014 50618
rect 37194 50566 37196 50618
rect 36950 50564 36956 50566
rect 37012 50564 37036 50566
rect 37092 50564 37116 50566
rect 37172 50564 37196 50566
rect 37252 50564 37258 50566
rect 36950 50555 37258 50564
rect 36950 49532 37258 49541
rect 36950 49530 36956 49532
rect 37012 49530 37036 49532
rect 37092 49530 37116 49532
rect 37172 49530 37196 49532
rect 37252 49530 37258 49532
rect 37012 49478 37014 49530
rect 37194 49478 37196 49530
rect 36950 49476 36956 49478
rect 37012 49476 37036 49478
rect 37092 49476 37116 49478
rect 37172 49476 37196 49478
rect 37252 49476 37258 49478
rect 36950 49467 37258 49476
rect 36950 48444 37258 48453
rect 36950 48442 36956 48444
rect 37012 48442 37036 48444
rect 37092 48442 37116 48444
rect 37172 48442 37196 48444
rect 37252 48442 37258 48444
rect 37012 48390 37014 48442
rect 37194 48390 37196 48442
rect 36950 48388 36956 48390
rect 37012 48388 37036 48390
rect 37092 48388 37116 48390
rect 37172 48388 37196 48390
rect 37252 48388 37258 48390
rect 36950 48379 37258 48388
rect 36950 47356 37258 47365
rect 36950 47354 36956 47356
rect 37012 47354 37036 47356
rect 37092 47354 37116 47356
rect 37172 47354 37196 47356
rect 37252 47354 37258 47356
rect 37012 47302 37014 47354
rect 37194 47302 37196 47354
rect 36950 47300 36956 47302
rect 37012 47300 37036 47302
rect 37092 47300 37116 47302
rect 37172 47300 37196 47302
rect 37252 47300 37258 47302
rect 36950 47291 37258 47300
rect 36728 46368 36780 46374
rect 36728 46310 36780 46316
rect 36950 46268 37258 46277
rect 36950 46266 36956 46268
rect 37012 46266 37036 46268
rect 37092 46266 37116 46268
rect 37172 46266 37196 46268
rect 37252 46266 37258 46268
rect 37012 46214 37014 46266
rect 37194 46214 37196 46266
rect 36950 46212 36956 46214
rect 37012 46212 37036 46214
rect 37092 46212 37116 46214
rect 37172 46212 37196 46214
rect 37252 46212 37258 46214
rect 36950 46203 37258 46212
rect 36950 45180 37258 45189
rect 36950 45178 36956 45180
rect 37012 45178 37036 45180
rect 37092 45178 37116 45180
rect 37172 45178 37196 45180
rect 37252 45178 37258 45180
rect 37012 45126 37014 45178
rect 37194 45126 37196 45178
rect 36950 45124 36956 45126
rect 37012 45124 37036 45126
rect 37092 45124 37116 45126
rect 37172 45124 37196 45126
rect 37252 45124 37258 45126
rect 36950 45115 37258 45124
rect 36950 44092 37258 44101
rect 36950 44090 36956 44092
rect 37012 44090 37036 44092
rect 37092 44090 37116 44092
rect 37172 44090 37196 44092
rect 37252 44090 37258 44092
rect 37012 44038 37014 44090
rect 37194 44038 37196 44090
rect 36950 44036 36956 44038
rect 37012 44036 37036 44038
rect 37092 44036 37116 44038
rect 37172 44036 37196 44038
rect 37252 44036 37258 44038
rect 36950 44027 37258 44036
rect 36636 43648 36688 43654
rect 36636 43590 36688 43596
rect 36950 43004 37258 43013
rect 36950 43002 36956 43004
rect 37012 43002 37036 43004
rect 37092 43002 37116 43004
rect 37172 43002 37196 43004
rect 37252 43002 37258 43004
rect 37012 42950 37014 43002
rect 37194 42950 37196 43002
rect 36950 42948 36956 42950
rect 37012 42948 37036 42950
rect 37092 42948 37116 42950
rect 37172 42948 37196 42950
rect 37252 42948 37258 42950
rect 36950 42939 37258 42948
rect 36950 41916 37258 41925
rect 36950 41914 36956 41916
rect 37012 41914 37036 41916
rect 37092 41914 37116 41916
rect 37172 41914 37196 41916
rect 37252 41914 37258 41916
rect 37012 41862 37014 41914
rect 37194 41862 37196 41914
rect 36950 41860 36956 41862
rect 37012 41860 37036 41862
rect 37092 41860 37116 41862
rect 37172 41860 37196 41862
rect 37252 41860 37258 41862
rect 36950 41851 37258 41860
rect 36636 41472 36688 41478
rect 36636 41414 36688 41420
rect 36544 35624 36596 35630
rect 36544 35566 36596 35572
rect 36452 33924 36504 33930
rect 36452 33866 36504 33872
rect 36360 30932 36412 30938
rect 36360 30874 36412 30880
rect 36188 30790 36400 30818
rect 36096 30654 36216 30682
rect 36084 30048 36136 30054
rect 36084 29990 36136 29996
rect 36096 29646 36124 29990
rect 36188 29850 36216 30654
rect 36268 30592 36320 30598
rect 36268 30534 36320 30540
rect 36176 29844 36228 29850
rect 36176 29786 36228 29792
rect 36084 29640 36136 29646
rect 36084 29582 36136 29588
rect 36176 29640 36228 29646
rect 36176 29582 36228 29588
rect 36188 29306 36216 29582
rect 36176 29300 36228 29306
rect 36176 29242 36228 29248
rect 35992 27872 36044 27878
rect 35992 27814 36044 27820
rect 36280 8362 36308 30534
rect 36372 24410 36400 30790
rect 36464 30598 36492 33866
rect 36556 32910 36584 35566
rect 36544 32904 36596 32910
rect 36544 32846 36596 32852
rect 36452 30592 36504 30598
rect 36452 30534 36504 30540
rect 36648 26586 36676 41414
rect 36950 40828 37258 40837
rect 36950 40826 36956 40828
rect 37012 40826 37036 40828
rect 37092 40826 37116 40828
rect 37172 40826 37196 40828
rect 37252 40826 37258 40828
rect 37012 40774 37014 40826
rect 37194 40774 37196 40826
rect 36950 40772 36956 40774
rect 37012 40772 37036 40774
rect 37092 40772 37116 40774
rect 37172 40772 37196 40774
rect 37252 40772 37258 40774
rect 36950 40763 37258 40772
rect 36728 39840 36780 39846
rect 36728 39782 36780 39788
rect 36740 34746 36768 39782
rect 36950 39740 37258 39749
rect 36950 39738 36956 39740
rect 37012 39738 37036 39740
rect 37092 39738 37116 39740
rect 37172 39738 37196 39740
rect 37252 39738 37258 39740
rect 37012 39686 37014 39738
rect 37194 39686 37196 39738
rect 36950 39684 36956 39686
rect 37012 39684 37036 39686
rect 37092 39684 37116 39686
rect 37172 39684 37196 39686
rect 37252 39684 37258 39686
rect 36950 39675 37258 39684
rect 36950 38652 37258 38661
rect 36950 38650 36956 38652
rect 37012 38650 37036 38652
rect 37092 38650 37116 38652
rect 37172 38650 37196 38652
rect 37252 38650 37258 38652
rect 37012 38598 37014 38650
rect 37194 38598 37196 38650
rect 36950 38596 36956 38598
rect 37012 38596 37036 38598
rect 37092 38596 37116 38598
rect 37172 38596 37196 38598
rect 37252 38596 37258 38598
rect 36950 38587 37258 38596
rect 36950 37564 37258 37573
rect 36950 37562 36956 37564
rect 37012 37562 37036 37564
rect 37092 37562 37116 37564
rect 37172 37562 37196 37564
rect 37252 37562 37258 37564
rect 37012 37510 37014 37562
rect 37194 37510 37196 37562
rect 36950 37508 36956 37510
rect 37012 37508 37036 37510
rect 37092 37508 37116 37510
rect 37172 37508 37196 37510
rect 37252 37508 37258 37510
rect 36950 37499 37258 37508
rect 36950 36476 37258 36485
rect 36950 36474 36956 36476
rect 37012 36474 37036 36476
rect 37092 36474 37116 36476
rect 37172 36474 37196 36476
rect 37252 36474 37258 36476
rect 37012 36422 37014 36474
rect 37194 36422 37196 36474
rect 36950 36420 36956 36422
rect 37012 36420 37036 36422
rect 37092 36420 37116 36422
rect 37172 36420 37196 36422
rect 37252 36420 37258 36422
rect 36950 36411 37258 36420
rect 36950 35388 37258 35397
rect 36950 35386 36956 35388
rect 37012 35386 37036 35388
rect 37092 35386 37116 35388
rect 37172 35386 37196 35388
rect 37252 35386 37258 35388
rect 37012 35334 37014 35386
rect 37194 35334 37196 35386
rect 36950 35332 36956 35334
rect 37012 35332 37036 35334
rect 37092 35332 37116 35334
rect 37172 35332 37196 35334
rect 37252 35332 37258 35334
rect 36950 35323 37258 35332
rect 36728 34740 36780 34746
rect 36728 34682 36780 34688
rect 36950 34300 37258 34309
rect 36950 34298 36956 34300
rect 37012 34298 37036 34300
rect 37092 34298 37116 34300
rect 37172 34298 37196 34300
rect 37252 34298 37258 34300
rect 37012 34246 37014 34298
rect 37194 34246 37196 34298
rect 36950 34244 36956 34246
rect 37012 34244 37036 34246
rect 37092 34244 37116 34246
rect 37172 34244 37196 34246
rect 37252 34244 37258 34246
rect 36950 34235 37258 34244
rect 36950 33212 37258 33221
rect 36950 33210 36956 33212
rect 37012 33210 37036 33212
rect 37092 33210 37116 33212
rect 37172 33210 37196 33212
rect 37252 33210 37258 33212
rect 37012 33158 37014 33210
rect 37194 33158 37196 33210
rect 36950 33156 36956 33158
rect 37012 33156 37036 33158
rect 37092 33156 37116 33158
rect 37172 33156 37196 33158
rect 37252 33156 37258 33158
rect 36950 33147 37258 33156
rect 36950 32124 37258 32133
rect 36950 32122 36956 32124
rect 37012 32122 37036 32124
rect 37092 32122 37116 32124
rect 37172 32122 37196 32124
rect 37252 32122 37258 32124
rect 37012 32070 37014 32122
rect 37194 32070 37196 32122
rect 36950 32068 36956 32070
rect 37012 32068 37036 32070
rect 37092 32068 37116 32070
rect 37172 32068 37196 32070
rect 37252 32068 37258 32070
rect 36950 32059 37258 32068
rect 36950 31036 37258 31045
rect 36950 31034 36956 31036
rect 37012 31034 37036 31036
rect 37092 31034 37116 31036
rect 37172 31034 37196 31036
rect 37252 31034 37258 31036
rect 37012 30982 37014 31034
rect 37194 30982 37196 31034
rect 36950 30980 36956 30982
rect 37012 30980 37036 30982
rect 37092 30980 37116 30982
rect 37172 30980 37196 30982
rect 37252 30980 37258 30982
rect 36950 30971 37258 30980
rect 36728 30864 36780 30870
rect 36728 30806 36780 30812
rect 36636 26580 36688 26586
rect 36636 26522 36688 26528
rect 36360 24404 36412 24410
rect 36360 24346 36412 24352
rect 36544 24132 36596 24138
rect 36544 24074 36596 24080
rect 36268 8356 36320 8362
rect 36268 8298 36320 8304
rect 36556 7954 36584 24074
rect 36740 17882 36768 30806
rect 36820 30728 36872 30734
rect 36820 30670 36872 30676
rect 36728 17876 36780 17882
rect 36728 17818 36780 17824
rect 36832 10538 36860 30670
rect 36950 29948 37258 29957
rect 36950 29946 36956 29948
rect 37012 29946 37036 29948
rect 37092 29946 37116 29948
rect 37172 29946 37196 29948
rect 37252 29946 37258 29948
rect 37012 29894 37014 29946
rect 37194 29894 37196 29946
rect 36950 29892 36956 29894
rect 37012 29892 37036 29894
rect 37092 29892 37116 29894
rect 37172 29892 37196 29894
rect 37252 29892 37258 29894
rect 36950 29883 37258 29892
rect 36950 28860 37258 28869
rect 36950 28858 36956 28860
rect 37012 28858 37036 28860
rect 37092 28858 37116 28860
rect 37172 28858 37196 28860
rect 37252 28858 37258 28860
rect 37012 28806 37014 28858
rect 37194 28806 37196 28858
rect 36950 28804 36956 28806
rect 37012 28804 37036 28806
rect 37092 28804 37116 28806
rect 37172 28804 37196 28806
rect 37252 28804 37258 28806
rect 36950 28795 37258 28804
rect 36950 27772 37258 27781
rect 36950 27770 36956 27772
rect 37012 27770 37036 27772
rect 37092 27770 37116 27772
rect 37172 27770 37196 27772
rect 37252 27770 37258 27772
rect 37012 27718 37014 27770
rect 37194 27718 37196 27770
rect 36950 27716 36956 27718
rect 37012 27716 37036 27718
rect 37092 27716 37116 27718
rect 37172 27716 37196 27718
rect 37252 27716 37258 27718
rect 36950 27707 37258 27716
rect 36950 26684 37258 26693
rect 36950 26682 36956 26684
rect 37012 26682 37036 26684
rect 37092 26682 37116 26684
rect 37172 26682 37196 26684
rect 37252 26682 37258 26684
rect 37012 26630 37014 26682
rect 37194 26630 37196 26682
rect 36950 26628 36956 26630
rect 37012 26628 37036 26630
rect 37092 26628 37116 26630
rect 37172 26628 37196 26630
rect 37252 26628 37258 26630
rect 36950 26619 37258 26628
rect 36950 25596 37258 25605
rect 36950 25594 36956 25596
rect 37012 25594 37036 25596
rect 37092 25594 37116 25596
rect 37172 25594 37196 25596
rect 37252 25594 37258 25596
rect 37012 25542 37014 25594
rect 37194 25542 37196 25594
rect 36950 25540 36956 25542
rect 37012 25540 37036 25542
rect 37092 25540 37116 25542
rect 37172 25540 37196 25542
rect 37252 25540 37258 25542
rect 36950 25531 37258 25540
rect 36950 24508 37258 24517
rect 36950 24506 36956 24508
rect 37012 24506 37036 24508
rect 37092 24506 37116 24508
rect 37172 24506 37196 24508
rect 37252 24506 37258 24508
rect 37012 24454 37014 24506
rect 37194 24454 37196 24506
rect 36950 24452 36956 24454
rect 37012 24452 37036 24454
rect 37092 24452 37116 24454
rect 37172 24452 37196 24454
rect 37252 24452 37258 24454
rect 36950 24443 37258 24452
rect 36950 23420 37258 23429
rect 36950 23418 36956 23420
rect 37012 23418 37036 23420
rect 37092 23418 37116 23420
rect 37172 23418 37196 23420
rect 37252 23418 37258 23420
rect 37012 23366 37014 23418
rect 37194 23366 37196 23418
rect 36950 23364 36956 23366
rect 37012 23364 37036 23366
rect 37092 23364 37116 23366
rect 37172 23364 37196 23366
rect 37252 23364 37258 23366
rect 36950 23355 37258 23364
rect 36950 22332 37258 22341
rect 36950 22330 36956 22332
rect 37012 22330 37036 22332
rect 37092 22330 37116 22332
rect 37172 22330 37196 22332
rect 37252 22330 37258 22332
rect 37012 22278 37014 22330
rect 37194 22278 37196 22330
rect 36950 22276 36956 22278
rect 37012 22276 37036 22278
rect 37092 22276 37116 22278
rect 37172 22276 37196 22278
rect 37252 22276 37258 22278
rect 36950 22267 37258 22276
rect 36950 21244 37258 21253
rect 36950 21242 36956 21244
rect 37012 21242 37036 21244
rect 37092 21242 37116 21244
rect 37172 21242 37196 21244
rect 37252 21242 37258 21244
rect 37012 21190 37014 21242
rect 37194 21190 37196 21242
rect 36950 21188 36956 21190
rect 37012 21188 37036 21190
rect 37092 21188 37116 21190
rect 37172 21188 37196 21190
rect 37252 21188 37258 21190
rect 36950 21179 37258 21188
rect 36950 20156 37258 20165
rect 36950 20154 36956 20156
rect 37012 20154 37036 20156
rect 37092 20154 37116 20156
rect 37172 20154 37196 20156
rect 37252 20154 37258 20156
rect 37012 20102 37014 20154
rect 37194 20102 37196 20154
rect 36950 20100 36956 20102
rect 37012 20100 37036 20102
rect 37092 20100 37116 20102
rect 37172 20100 37196 20102
rect 37252 20100 37258 20102
rect 36950 20091 37258 20100
rect 36950 19068 37258 19077
rect 36950 19066 36956 19068
rect 37012 19066 37036 19068
rect 37092 19066 37116 19068
rect 37172 19066 37196 19068
rect 37252 19066 37258 19068
rect 37012 19014 37014 19066
rect 37194 19014 37196 19066
rect 36950 19012 36956 19014
rect 37012 19012 37036 19014
rect 37092 19012 37116 19014
rect 37172 19012 37196 19014
rect 37252 19012 37258 19014
rect 36950 19003 37258 19012
rect 36950 17980 37258 17989
rect 36950 17978 36956 17980
rect 37012 17978 37036 17980
rect 37092 17978 37116 17980
rect 37172 17978 37196 17980
rect 37252 17978 37258 17980
rect 37012 17926 37014 17978
rect 37194 17926 37196 17978
rect 36950 17924 36956 17926
rect 37012 17924 37036 17926
rect 37092 17924 37116 17926
rect 37172 17924 37196 17926
rect 37252 17924 37258 17926
rect 36950 17915 37258 17924
rect 36950 16892 37258 16901
rect 36950 16890 36956 16892
rect 37012 16890 37036 16892
rect 37092 16890 37116 16892
rect 37172 16890 37196 16892
rect 37252 16890 37258 16892
rect 37012 16838 37014 16890
rect 37194 16838 37196 16890
rect 36950 16836 36956 16838
rect 37012 16836 37036 16838
rect 37092 16836 37116 16838
rect 37172 16836 37196 16838
rect 37252 16836 37258 16838
rect 36950 16827 37258 16836
rect 36950 15804 37258 15813
rect 36950 15802 36956 15804
rect 37012 15802 37036 15804
rect 37092 15802 37116 15804
rect 37172 15802 37196 15804
rect 37252 15802 37258 15804
rect 37012 15750 37014 15802
rect 37194 15750 37196 15802
rect 36950 15748 36956 15750
rect 37012 15748 37036 15750
rect 37092 15748 37116 15750
rect 37172 15748 37196 15750
rect 37252 15748 37258 15750
rect 36950 15739 37258 15748
rect 36950 14716 37258 14725
rect 36950 14714 36956 14716
rect 37012 14714 37036 14716
rect 37092 14714 37116 14716
rect 37172 14714 37196 14716
rect 37252 14714 37258 14716
rect 37012 14662 37014 14714
rect 37194 14662 37196 14714
rect 36950 14660 36956 14662
rect 37012 14660 37036 14662
rect 37092 14660 37116 14662
rect 37172 14660 37196 14662
rect 37252 14660 37258 14662
rect 36950 14651 37258 14660
rect 36950 13628 37258 13637
rect 36950 13626 36956 13628
rect 37012 13626 37036 13628
rect 37092 13626 37116 13628
rect 37172 13626 37196 13628
rect 37252 13626 37258 13628
rect 37012 13574 37014 13626
rect 37194 13574 37196 13626
rect 36950 13572 36956 13574
rect 37012 13572 37036 13574
rect 37092 13572 37116 13574
rect 37172 13572 37196 13574
rect 37252 13572 37258 13574
rect 36950 13563 37258 13572
rect 36950 12540 37258 12549
rect 36950 12538 36956 12540
rect 37012 12538 37036 12540
rect 37092 12538 37116 12540
rect 37172 12538 37196 12540
rect 37252 12538 37258 12540
rect 37012 12486 37014 12538
rect 37194 12486 37196 12538
rect 36950 12484 36956 12486
rect 37012 12484 37036 12486
rect 37092 12484 37116 12486
rect 37172 12484 37196 12486
rect 37252 12484 37258 12486
rect 36950 12475 37258 12484
rect 36950 11452 37258 11461
rect 36950 11450 36956 11452
rect 37012 11450 37036 11452
rect 37092 11450 37116 11452
rect 37172 11450 37196 11452
rect 37252 11450 37258 11452
rect 37012 11398 37014 11450
rect 37194 11398 37196 11450
rect 36950 11396 36956 11398
rect 37012 11396 37036 11398
rect 37092 11396 37116 11398
rect 37172 11396 37196 11398
rect 37252 11396 37258 11398
rect 36950 11387 37258 11396
rect 36820 10532 36872 10538
rect 36820 10474 36872 10480
rect 36950 10364 37258 10373
rect 36950 10362 36956 10364
rect 37012 10362 37036 10364
rect 37092 10362 37116 10364
rect 37172 10362 37196 10364
rect 37252 10362 37258 10364
rect 37012 10310 37014 10362
rect 37194 10310 37196 10362
rect 36950 10308 36956 10310
rect 37012 10308 37036 10310
rect 37092 10308 37116 10310
rect 37172 10308 37196 10310
rect 37252 10308 37258 10310
rect 36950 10299 37258 10308
rect 36950 9276 37258 9285
rect 36950 9274 36956 9276
rect 37012 9274 37036 9276
rect 37092 9274 37116 9276
rect 37172 9274 37196 9276
rect 37252 9274 37258 9276
rect 37012 9222 37014 9274
rect 37194 9222 37196 9274
rect 36950 9220 36956 9222
rect 37012 9220 37036 9222
rect 37092 9220 37116 9222
rect 37172 9220 37196 9222
rect 37252 9220 37258 9222
rect 36950 9211 37258 9220
rect 36950 8188 37258 8197
rect 36950 8186 36956 8188
rect 37012 8186 37036 8188
rect 37092 8186 37116 8188
rect 37172 8186 37196 8188
rect 37252 8186 37258 8188
rect 37012 8134 37014 8186
rect 37194 8134 37196 8186
rect 36950 8132 36956 8134
rect 37012 8132 37036 8134
rect 37092 8132 37116 8134
rect 37172 8132 37196 8134
rect 37252 8132 37258 8134
rect 36950 8123 37258 8132
rect 36544 7948 36596 7954
rect 36544 7890 36596 7896
rect 36950 7100 37258 7109
rect 36950 7098 36956 7100
rect 37012 7098 37036 7100
rect 37092 7098 37116 7100
rect 37172 7098 37196 7100
rect 37252 7098 37258 7100
rect 37012 7046 37014 7098
rect 37194 7046 37196 7098
rect 36950 7044 36956 7046
rect 37012 7044 37036 7046
rect 37092 7044 37116 7046
rect 37172 7044 37196 7046
rect 37252 7044 37258 7046
rect 36950 7035 37258 7044
rect 37292 6914 37320 55186
rect 37610 54428 37918 54437
rect 37610 54426 37616 54428
rect 37672 54426 37696 54428
rect 37752 54426 37776 54428
rect 37832 54426 37856 54428
rect 37912 54426 37918 54428
rect 37672 54374 37674 54426
rect 37854 54374 37856 54426
rect 37610 54372 37616 54374
rect 37672 54372 37696 54374
rect 37752 54372 37776 54374
rect 37832 54372 37856 54374
rect 37912 54372 37918 54374
rect 37610 54363 37918 54372
rect 37610 53340 37918 53349
rect 37610 53338 37616 53340
rect 37672 53338 37696 53340
rect 37752 53338 37776 53340
rect 37832 53338 37856 53340
rect 37912 53338 37918 53340
rect 37672 53286 37674 53338
rect 37854 53286 37856 53338
rect 37610 53284 37616 53286
rect 37672 53284 37696 53286
rect 37752 53284 37776 53286
rect 37832 53284 37856 53286
rect 37912 53284 37918 53286
rect 37610 53275 37918 53284
rect 37610 52252 37918 52261
rect 37610 52250 37616 52252
rect 37672 52250 37696 52252
rect 37752 52250 37776 52252
rect 37832 52250 37856 52252
rect 37912 52250 37918 52252
rect 37672 52198 37674 52250
rect 37854 52198 37856 52250
rect 37610 52196 37616 52198
rect 37672 52196 37696 52198
rect 37752 52196 37776 52198
rect 37832 52196 37856 52198
rect 37912 52196 37918 52198
rect 37610 52187 37918 52196
rect 37610 51164 37918 51173
rect 37610 51162 37616 51164
rect 37672 51162 37696 51164
rect 37752 51162 37776 51164
rect 37832 51162 37856 51164
rect 37912 51162 37918 51164
rect 37672 51110 37674 51162
rect 37854 51110 37856 51162
rect 37610 51108 37616 51110
rect 37672 51108 37696 51110
rect 37752 51108 37776 51110
rect 37832 51108 37856 51110
rect 37912 51108 37918 51110
rect 37610 51099 37918 51108
rect 37464 51060 37516 51066
rect 37464 51002 37516 51008
rect 37372 49156 37424 49162
rect 37372 49098 37424 49104
rect 37384 48890 37412 49098
rect 37372 48884 37424 48890
rect 37372 48826 37424 48832
rect 37476 48770 37504 51002
rect 37610 50076 37918 50085
rect 37610 50074 37616 50076
rect 37672 50074 37696 50076
rect 37752 50074 37776 50076
rect 37832 50074 37856 50076
rect 37912 50074 37918 50076
rect 37672 50022 37674 50074
rect 37854 50022 37856 50074
rect 37610 50020 37616 50022
rect 37672 50020 37696 50022
rect 37752 50020 37776 50022
rect 37832 50020 37856 50022
rect 37912 50020 37918 50022
rect 37610 50011 37918 50020
rect 37610 48988 37918 48997
rect 37610 48986 37616 48988
rect 37672 48986 37696 48988
rect 37752 48986 37776 48988
rect 37832 48986 37856 48988
rect 37912 48986 37918 48988
rect 37672 48934 37674 48986
rect 37854 48934 37856 48986
rect 37610 48932 37616 48934
rect 37672 48932 37696 48934
rect 37752 48932 37776 48934
rect 37832 48932 37856 48934
rect 37912 48932 37918 48934
rect 37610 48923 37918 48932
rect 37384 48742 37504 48770
rect 37384 26874 37412 48742
rect 37464 48680 37516 48686
rect 37464 48622 37516 48628
rect 37476 27010 37504 48622
rect 37610 47900 37918 47909
rect 37610 47898 37616 47900
rect 37672 47898 37696 47900
rect 37752 47898 37776 47900
rect 37832 47898 37856 47900
rect 37912 47898 37918 47900
rect 37672 47846 37674 47898
rect 37854 47846 37856 47898
rect 37610 47844 37616 47846
rect 37672 47844 37696 47846
rect 37752 47844 37776 47846
rect 37832 47844 37856 47846
rect 37912 47844 37918 47846
rect 37610 47835 37918 47844
rect 37610 46812 37918 46821
rect 37610 46810 37616 46812
rect 37672 46810 37696 46812
rect 37752 46810 37776 46812
rect 37832 46810 37856 46812
rect 37912 46810 37918 46812
rect 37672 46758 37674 46810
rect 37854 46758 37856 46810
rect 37610 46756 37616 46758
rect 37672 46756 37696 46758
rect 37752 46756 37776 46758
rect 37832 46756 37856 46758
rect 37912 46756 37918 46758
rect 37610 46747 37918 46756
rect 37610 45724 37918 45733
rect 37610 45722 37616 45724
rect 37672 45722 37696 45724
rect 37752 45722 37776 45724
rect 37832 45722 37856 45724
rect 37912 45722 37918 45724
rect 37672 45670 37674 45722
rect 37854 45670 37856 45722
rect 37610 45668 37616 45670
rect 37672 45668 37696 45670
rect 37752 45668 37776 45670
rect 37832 45668 37856 45670
rect 37912 45668 37918 45670
rect 37610 45659 37918 45668
rect 37610 44636 37918 44645
rect 37610 44634 37616 44636
rect 37672 44634 37696 44636
rect 37752 44634 37776 44636
rect 37832 44634 37856 44636
rect 37912 44634 37918 44636
rect 37672 44582 37674 44634
rect 37854 44582 37856 44634
rect 37610 44580 37616 44582
rect 37672 44580 37696 44582
rect 37752 44580 37776 44582
rect 37832 44580 37856 44582
rect 37912 44580 37918 44582
rect 37610 44571 37918 44580
rect 37610 43548 37918 43557
rect 37610 43546 37616 43548
rect 37672 43546 37696 43548
rect 37752 43546 37776 43548
rect 37832 43546 37856 43548
rect 37912 43546 37918 43548
rect 37672 43494 37674 43546
rect 37854 43494 37856 43546
rect 37610 43492 37616 43494
rect 37672 43492 37696 43494
rect 37752 43492 37776 43494
rect 37832 43492 37856 43494
rect 37912 43492 37918 43494
rect 37610 43483 37918 43492
rect 37610 42460 37918 42469
rect 37610 42458 37616 42460
rect 37672 42458 37696 42460
rect 37752 42458 37776 42460
rect 37832 42458 37856 42460
rect 37912 42458 37918 42460
rect 37672 42406 37674 42458
rect 37854 42406 37856 42458
rect 37610 42404 37616 42406
rect 37672 42404 37696 42406
rect 37752 42404 37776 42406
rect 37832 42404 37856 42406
rect 37912 42404 37918 42406
rect 37610 42395 37918 42404
rect 37610 41372 37918 41381
rect 37610 41370 37616 41372
rect 37672 41370 37696 41372
rect 37752 41370 37776 41372
rect 37832 41370 37856 41372
rect 37912 41370 37918 41372
rect 37672 41318 37674 41370
rect 37854 41318 37856 41370
rect 37610 41316 37616 41318
rect 37672 41316 37696 41318
rect 37752 41316 37776 41318
rect 37832 41316 37856 41318
rect 37912 41316 37918 41318
rect 37610 41307 37918 41316
rect 37610 40284 37918 40293
rect 37610 40282 37616 40284
rect 37672 40282 37696 40284
rect 37752 40282 37776 40284
rect 37832 40282 37856 40284
rect 37912 40282 37918 40284
rect 37672 40230 37674 40282
rect 37854 40230 37856 40282
rect 37610 40228 37616 40230
rect 37672 40228 37696 40230
rect 37752 40228 37776 40230
rect 37832 40228 37856 40230
rect 37912 40228 37918 40230
rect 37610 40219 37918 40228
rect 37610 39196 37918 39205
rect 37610 39194 37616 39196
rect 37672 39194 37696 39196
rect 37752 39194 37776 39196
rect 37832 39194 37856 39196
rect 37912 39194 37918 39196
rect 37672 39142 37674 39194
rect 37854 39142 37856 39194
rect 37610 39140 37616 39142
rect 37672 39140 37696 39142
rect 37752 39140 37776 39142
rect 37832 39140 37856 39142
rect 37912 39140 37918 39142
rect 37610 39131 37918 39140
rect 37610 38108 37918 38117
rect 37610 38106 37616 38108
rect 37672 38106 37696 38108
rect 37752 38106 37776 38108
rect 37832 38106 37856 38108
rect 37912 38106 37918 38108
rect 37672 38054 37674 38106
rect 37854 38054 37856 38106
rect 37610 38052 37616 38054
rect 37672 38052 37696 38054
rect 37752 38052 37776 38054
rect 37832 38052 37856 38054
rect 37912 38052 37918 38054
rect 37610 38043 37918 38052
rect 38016 37120 38068 37126
rect 38016 37062 38068 37068
rect 37610 37020 37918 37029
rect 37610 37018 37616 37020
rect 37672 37018 37696 37020
rect 37752 37018 37776 37020
rect 37832 37018 37856 37020
rect 37912 37018 37918 37020
rect 37672 36966 37674 37018
rect 37854 36966 37856 37018
rect 37610 36964 37616 36966
rect 37672 36964 37696 36966
rect 37752 36964 37776 36966
rect 37832 36964 37856 36966
rect 37912 36964 37918 36966
rect 37610 36955 37918 36964
rect 38028 36786 38056 37062
rect 38120 36854 38148 55186
rect 38292 53576 38344 53582
rect 38292 53518 38344 53524
rect 38200 52488 38252 52494
rect 38200 52430 38252 52436
rect 38212 39438 38240 52430
rect 38304 52018 38332 53518
rect 38292 52012 38344 52018
rect 38292 51954 38344 51960
rect 38396 48754 38424 67594
rect 38844 67312 38896 67318
rect 38844 67254 38896 67260
rect 40498 67280 40554 67289
rect 38660 60716 38712 60722
rect 38660 60658 38712 60664
rect 38752 60716 38804 60722
rect 38752 60658 38804 60664
rect 38384 48748 38436 48754
rect 38384 48690 38436 48696
rect 38672 41478 38700 60658
rect 38764 52970 38792 60658
rect 38856 60654 38884 67254
rect 40498 67215 40500 67224
rect 40552 67215 40554 67224
rect 40500 67186 40552 67192
rect 39580 66224 39632 66230
rect 39580 66166 39632 66172
rect 38844 60648 38896 60654
rect 38844 60590 38896 60596
rect 39120 60512 39172 60518
rect 39120 60454 39172 60460
rect 39132 60314 39160 60454
rect 39120 60308 39172 60314
rect 39120 60250 39172 60256
rect 39304 58608 39356 58614
rect 39304 58550 39356 58556
rect 39120 58540 39172 58546
rect 39120 58482 39172 58488
rect 39132 57610 39160 58482
rect 38856 57582 39160 57610
rect 38752 52964 38804 52970
rect 38752 52906 38804 52912
rect 38856 48006 38884 57582
rect 38936 57452 38988 57458
rect 38936 57394 38988 57400
rect 39212 57452 39264 57458
rect 39212 57394 39264 57400
rect 38844 48000 38896 48006
rect 38844 47942 38896 47948
rect 38844 47796 38896 47802
rect 38844 47738 38896 47744
rect 38752 45008 38804 45014
rect 38752 44950 38804 44956
rect 38660 41472 38712 41478
rect 38660 41414 38712 41420
rect 38660 40384 38712 40390
rect 38660 40326 38712 40332
rect 38200 39432 38252 39438
rect 38200 39374 38252 39380
rect 38384 38004 38436 38010
rect 38384 37946 38436 37952
rect 38108 36848 38160 36854
rect 38108 36790 38160 36796
rect 38016 36780 38068 36786
rect 38016 36722 38068 36728
rect 37610 35932 37918 35941
rect 37610 35930 37616 35932
rect 37672 35930 37696 35932
rect 37752 35930 37776 35932
rect 37832 35930 37856 35932
rect 37912 35930 37918 35932
rect 37672 35878 37674 35930
rect 37854 35878 37856 35930
rect 37610 35876 37616 35878
rect 37672 35876 37696 35878
rect 37752 35876 37776 35878
rect 37832 35876 37856 35878
rect 37912 35876 37918 35878
rect 37610 35867 37918 35876
rect 38396 34950 38424 37946
rect 38568 36712 38620 36718
rect 38568 36654 38620 36660
rect 38384 34944 38436 34950
rect 38384 34886 38436 34892
rect 37610 34844 37918 34853
rect 37610 34842 37616 34844
rect 37672 34842 37696 34844
rect 37752 34842 37776 34844
rect 37832 34842 37856 34844
rect 37912 34842 37918 34844
rect 37672 34790 37674 34842
rect 37854 34790 37856 34842
rect 37610 34788 37616 34790
rect 37672 34788 37696 34790
rect 37752 34788 37776 34790
rect 37832 34788 37856 34790
rect 37912 34788 37918 34790
rect 37610 34779 37918 34788
rect 37610 33756 37918 33765
rect 37610 33754 37616 33756
rect 37672 33754 37696 33756
rect 37752 33754 37776 33756
rect 37832 33754 37856 33756
rect 37912 33754 37918 33756
rect 37672 33702 37674 33754
rect 37854 33702 37856 33754
rect 37610 33700 37616 33702
rect 37672 33700 37696 33702
rect 37752 33700 37776 33702
rect 37832 33700 37856 33702
rect 37912 33700 37918 33702
rect 37610 33691 37918 33700
rect 38200 32904 38252 32910
rect 38200 32846 38252 32852
rect 38212 32774 38240 32846
rect 38200 32768 38252 32774
rect 38200 32710 38252 32716
rect 37610 32668 37918 32677
rect 37610 32666 37616 32668
rect 37672 32666 37696 32668
rect 37752 32666 37776 32668
rect 37832 32666 37856 32668
rect 37912 32666 37918 32668
rect 37672 32614 37674 32666
rect 37854 32614 37856 32666
rect 37610 32612 37616 32614
rect 37672 32612 37696 32614
rect 37752 32612 37776 32614
rect 37832 32612 37856 32614
rect 37912 32612 37918 32614
rect 37610 32603 37918 32612
rect 37610 31580 37918 31589
rect 37610 31578 37616 31580
rect 37672 31578 37696 31580
rect 37752 31578 37776 31580
rect 37832 31578 37856 31580
rect 37912 31578 37918 31580
rect 37672 31526 37674 31578
rect 37854 31526 37856 31578
rect 37610 31524 37616 31526
rect 37672 31524 37696 31526
rect 37752 31524 37776 31526
rect 37832 31524 37856 31526
rect 37912 31524 37918 31526
rect 37610 31515 37918 31524
rect 37610 30492 37918 30501
rect 37610 30490 37616 30492
rect 37672 30490 37696 30492
rect 37752 30490 37776 30492
rect 37832 30490 37856 30492
rect 37912 30490 37918 30492
rect 37672 30438 37674 30490
rect 37854 30438 37856 30490
rect 37610 30436 37616 30438
rect 37672 30436 37696 30438
rect 37752 30436 37776 30438
rect 37832 30436 37856 30438
rect 37912 30436 37918 30438
rect 37610 30427 37918 30436
rect 37610 29404 37918 29413
rect 37610 29402 37616 29404
rect 37672 29402 37696 29404
rect 37752 29402 37776 29404
rect 37832 29402 37856 29404
rect 37912 29402 37918 29404
rect 37672 29350 37674 29402
rect 37854 29350 37856 29402
rect 37610 29348 37616 29350
rect 37672 29348 37696 29350
rect 37752 29348 37776 29350
rect 37832 29348 37856 29350
rect 37912 29348 37918 29350
rect 37610 29339 37918 29348
rect 37610 28316 37918 28325
rect 37610 28314 37616 28316
rect 37672 28314 37696 28316
rect 37752 28314 37776 28316
rect 37832 28314 37856 28316
rect 37912 28314 37918 28316
rect 37672 28262 37674 28314
rect 37854 28262 37856 28314
rect 37610 28260 37616 28262
rect 37672 28260 37696 28262
rect 37752 28260 37776 28262
rect 37832 28260 37856 28262
rect 37912 28260 37918 28262
rect 37610 28251 37918 28260
rect 37610 27228 37918 27237
rect 37610 27226 37616 27228
rect 37672 27226 37696 27228
rect 37752 27226 37776 27228
rect 37832 27226 37856 27228
rect 37912 27226 37918 27228
rect 37672 27174 37674 27226
rect 37854 27174 37856 27226
rect 37610 27172 37616 27174
rect 37672 27172 37696 27174
rect 37752 27172 37776 27174
rect 37832 27172 37856 27174
rect 37912 27172 37918 27174
rect 37610 27163 37918 27172
rect 37476 26982 37596 27010
rect 37384 26846 37504 26874
rect 37372 26240 37424 26246
rect 37372 26182 37424 26188
rect 37384 22982 37412 26182
rect 37372 22976 37424 22982
rect 37372 22918 37424 22924
rect 37372 22772 37424 22778
rect 37372 22714 37424 22720
rect 37384 19854 37412 22714
rect 37476 22094 37504 26846
rect 37568 26246 37596 26982
rect 37556 26240 37608 26246
rect 37556 26182 37608 26188
rect 37610 26140 37918 26149
rect 37610 26138 37616 26140
rect 37672 26138 37696 26140
rect 37752 26138 37776 26140
rect 37832 26138 37856 26140
rect 37912 26138 37918 26140
rect 37672 26086 37674 26138
rect 37854 26086 37856 26138
rect 37610 26084 37616 26086
rect 37672 26084 37696 26086
rect 37752 26084 37776 26086
rect 37832 26084 37856 26086
rect 37912 26084 37918 26086
rect 37610 26075 37918 26084
rect 38212 25362 38240 32710
rect 38292 31272 38344 31278
rect 38292 31214 38344 31220
rect 38200 25356 38252 25362
rect 38200 25298 38252 25304
rect 37610 25052 37918 25061
rect 37610 25050 37616 25052
rect 37672 25050 37696 25052
rect 37752 25050 37776 25052
rect 37832 25050 37856 25052
rect 37912 25050 37918 25052
rect 37672 24998 37674 25050
rect 37854 24998 37856 25050
rect 37610 24996 37616 24998
rect 37672 24996 37696 24998
rect 37752 24996 37776 24998
rect 37832 24996 37856 24998
rect 37912 24996 37918 24998
rect 37610 24987 37918 24996
rect 38304 24750 38332 31214
rect 38396 25294 38424 34886
rect 38580 34542 38608 36654
rect 38568 34536 38620 34542
rect 38568 34478 38620 34484
rect 38580 26926 38608 34478
rect 38568 26920 38620 26926
rect 38568 26862 38620 26868
rect 38384 25288 38436 25294
rect 38384 25230 38436 25236
rect 38292 24744 38344 24750
rect 38292 24686 38344 24692
rect 37610 23964 37918 23973
rect 37610 23962 37616 23964
rect 37672 23962 37696 23964
rect 37752 23962 37776 23964
rect 37832 23962 37856 23964
rect 37912 23962 37918 23964
rect 37672 23910 37674 23962
rect 37854 23910 37856 23962
rect 37610 23908 37616 23910
rect 37672 23908 37696 23910
rect 37752 23908 37776 23910
rect 37832 23908 37856 23910
rect 37912 23908 37918 23910
rect 37610 23899 37918 23908
rect 37610 22876 37918 22885
rect 37610 22874 37616 22876
rect 37672 22874 37696 22876
rect 37752 22874 37776 22876
rect 37832 22874 37856 22876
rect 37912 22874 37918 22876
rect 37672 22822 37674 22874
rect 37854 22822 37856 22874
rect 37610 22820 37616 22822
rect 37672 22820 37696 22822
rect 37752 22820 37776 22822
rect 37832 22820 37856 22822
rect 37912 22820 37918 22822
rect 37610 22811 37918 22820
rect 37476 22066 38056 22094
rect 37610 21788 37918 21797
rect 37610 21786 37616 21788
rect 37672 21786 37696 21788
rect 37752 21786 37776 21788
rect 37832 21786 37856 21788
rect 37912 21786 37918 21788
rect 37672 21734 37674 21786
rect 37854 21734 37856 21786
rect 37610 21732 37616 21734
rect 37672 21732 37696 21734
rect 37752 21732 37776 21734
rect 37832 21732 37856 21734
rect 37912 21732 37918 21734
rect 37610 21723 37918 21732
rect 37610 20700 37918 20709
rect 37610 20698 37616 20700
rect 37672 20698 37696 20700
rect 37752 20698 37776 20700
rect 37832 20698 37856 20700
rect 37912 20698 37918 20700
rect 37672 20646 37674 20698
rect 37854 20646 37856 20698
rect 37610 20644 37616 20646
rect 37672 20644 37696 20646
rect 37752 20644 37776 20646
rect 37832 20644 37856 20646
rect 37912 20644 37918 20646
rect 37610 20635 37918 20644
rect 37464 20596 37516 20602
rect 37464 20538 37516 20544
rect 37476 19922 37504 20538
rect 38028 19990 38056 22066
rect 38016 19984 38068 19990
rect 38016 19926 38068 19932
rect 37464 19916 37516 19922
rect 37464 19858 37516 19864
rect 37372 19848 37424 19854
rect 37372 19790 37424 19796
rect 37610 19612 37918 19621
rect 37610 19610 37616 19612
rect 37672 19610 37696 19612
rect 37752 19610 37776 19612
rect 37832 19610 37856 19612
rect 37912 19610 37918 19612
rect 37672 19558 37674 19610
rect 37854 19558 37856 19610
rect 37610 19556 37616 19558
rect 37672 19556 37696 19558
rect 37752 19556 37776 19558
rect 37832 19556 37856 19558
rect 37912 19556 37918 19558
rect 37610 19547 37918 19556
rect 37610 18524 37918 18533
rect 37610 18522 37616 18524
rect 37672 18522 37696 18524
rect 37752 18522 37776 18524
rect 37832 18522 37856 18524
rect 37912 18522 37918 18524
rect 37672 18470 37674 18522
rect 37854 18470 37856 18522
rect 37610 18468 37616 18470
rect 37672 18468 37696 18470
rect 37752 18468 37776 18470
rect 37832 18468 37856 18470
rect 37912 18468 37918 18470
rect 37610 18459 37918 18468
rect 37372 18080 37424 18086
rect 37372 18022 37424 18028
rect 37384 15094 37412 18022
rect 37610 17436 37918 17445
rect 37610 17434 37616 17436
rect 37672 17434 37696 17436
rect 37752 17434 37776 17436
rect 37832 17434 37856 17436
rect 37912 17434 37918 17436
rect 37672 17382 37674 17434
rect 37854 17382 37856 17434
rect 37610 17380 37616 17382
rect 37672 17380 37696 17382
rect 37752 17380 37776 17382
rect 37832 17380 37856 17382
rect 37912 17380 37918 17382
rect 37610 17371 37918 17380
rect 38028 16574 38056 19926
rect 38028 16546 38148 16574
rect 37610 16348 37918 16357
rect 37610 16346 37616 16348
rect 37672 16346 37696 16348
rect 37752 16346 37776 16348
rect 37832 16346 37856 16348
rect 37912 16346 37918 16348
rect 37672 16294 37674 16346
rect 37854 16294 37856 16346
rect 37610 16292 37616 16294
rect 37672 16292 37696 16294
rect 37752 16292 37776 16294
rect 37832 16292 37856 16294
rect 37912 16292 37918 16294
rect 37610 16283 37918 16292
rect 37610 15260 37918 15269
rect 37610 15258 37616 15260
rect 37672 15258 37696 15260
rect 37752 15258 37776 15260
rect 37832 15258 37856 15260
rect 37912 15258 37918 15260
rect 37672 15206 37674 15258
rect 37854 15206 37856 15258
rect 37610 15204 37616 15206
rect 37672 15204 37696 15206
rect 37752 15204 37776 15206
rect 37832 15204 37856 15206
rect 37912 15204 37918 15206
rect 37610 15195 37918 15204
rect 37372 15088 37424 15094
rect 37372 15030 37424 15036
rect 37610 14172 37918 14181
rect 37610 14170 37616 14172
rect 37672 14170 37696 14172
rect 37752 14170 37776 14172
rect 37832 14170 37856 14172
rect 37912 14170 37918 14172
rect 37672 14118 37674 14170
rect 37854 14118 37856 14170
rect 37610 14116 37616 14118
rect 37672 14116 37696 14118
rect 37752 14116 37776 14118
rect 37832 14116 37856 14118
rect 37912 14116 37918 14118
rect 37610 14107 37918 14116
rect 37610 13084 37918 13093
rect 37610 13082 37616 13084
rect 37672 13082 37696 13084
rect 37752 13082 37776 13084
rect 37832 13082 37856 13084
rect 37912 13082 37918 13084
rect 37672 13030 37674 13082
rect 37854 13030 37856 13082
rect 37610 13028 37616 13030
rect 37672 13028 37696 13030
rect 37752 13028 37776 13030
rect 37832 13028 37856 13030
rect 37912 13028 37918 13030
rect 37610 13019 37918 13028
rect 37610 11996 37918 12005
rect 37610 11994 37616 11996
rect 37672 11994 37696 11996
rect 37752 11994 37776 11996
rect 37832 11994 37856 11996
rect 37912 11994 37918 11996
rect 37672 11942 37674 11994
rect 37854 11942 37856 11994
rect 37610 11940 37616 11942
rect 37672 11940 37696 11942
rect 37752 11940 37776 11942
rect 37832 11940 37856 11942
rect 37912 11940 37918 11942
rect 37610 11931 37918 11940
rect 37610 10908 37918 10917
rect 37610 10906 37616 10908
rect 37672 10906 37696 10908
rect 37752 10906 37776 10908
rect 37832 10906 37856 10908
rect 37912 10906 37918 10908
rect 37672 10854 37674 10906
rect 37854 10854 37856 10906
rect 37610 10852 37616 10854
rect 37672 10852 37696 10854
rect 37752 10852 37776 10854
rect 37832 10852 37856 10854
rect 37912 10852 37918 10854
rect 37610 10843 37918 10852
rect 37610 9820 37918 9829
rect 37610 9818 37616 9820
rect 37672 9818 37696 9820
rect 37752 9818 37776 9820
rect 37832 9818 37856 9820
rect 37912 9818 37918 9820
rect 37672 9766 37674 9818
rect 37854 9766 37856 9818
rect 37610 9764 37616 9766
rect 37672 9764 37696 9766
rect 37752 9764 37776 9766
rect 37832 9764 37856 9766
rect 37912 9764 37918 9766
rect 37610 9755 37918 9764
rect 37610 8732 37918 8741
rect 37610 8730 37616 8732
rect 37672 8730 37696 8732
rect 37752 8730 37776 8732
rect 37832 8730 37856 8732
rect 37912 8730 37918 8732
rect 37672 8678 37674 8730
rect 37854 8678 37856 8730
rect 37610 8676 37616 8678
rect 37672 8676 37696 8678
rect 37752 8676 37776 8678
rect 37832 8676 37856 8678
rect 37912 8676 37918 8678
rect 37610 8667 37918 8676
rect 37610 7644 37918 7653
rect 37610 7642 37616 7644
rect 37672 7642 37696 7644
rect 37752 7642 37776 7644
rect 37832 7642 37856 7644
rect 37912 7642 37918 7644
rect 37672 7590 37674 7642
rect 37854 7590 37856 7642
rect 37610 7588 37616 7590
rect 37672 7588 37696 7590
rect 37752 7588 37776 7590
rect 37832 7588 37856 7590
rect 37912 7588 37918 7590
rect 37610 7579 37918 7588
rect 37292 6886 37504 6914
rect 37280 6724 37332 6730
rect 37280 6666 37332 6672
rect 36950 6012 37258 6021
rect 36950 6010 36956 6012
rect 37012 6010 37036 6012
rect 37092 6010 37116 6012
rect 37172 6010 37196 6012
rect 37252 6010 37258 6012
rect 37012 5958 37014 6010
rect 37194 5958 37196 6010
rect 36950 5956 36956 5958
rect 37012 5956 37036 5958
rect 37092 5956 37116 5958
rect 37172 5956 37196 5958
rect 37252 5956 37258 5958
rect 36950 5947 37258 5956
rect 36950 4924 37258 4933
rect 36950 4922 36956 4924
rect 37012 4922 37036 4924
rect 37092 4922 37116 4924
rect 37172 4922 37196 4924
rect 37252 4922 37258 4924
rect 37012 4870 37014 4922
rect 37194 4870 37196 4922
rect 36950 4868 36956 4870
rect 37012 4868 37036 4870
rect 37092 4868 37116 4870
rect 37172 4868 37196 4870
rect 37252 4868 37258 4870
rect 36950 4859 37258 4868
rect 37292 4554 37320 6666
rect 37372 6452 37424 6458
rect 37372 6394 37424 6400
rect 37384 4690 37412 6394
rect 37476 5030 37504 6886
rect 37610 6556 37918 6565
rect 37610 6554 37616 6556
rect 37672 6554 37696 6556
rect 37752 6554 37776 6556
rect 37832 6554 37856 6556
rect 37912 6554 37918 6556
rect 37672 6502 37674 6554
rect 37854 6502 37856 6554
rect 37610 6500 37616 6502
rect 37672 6500 37696 6502
rect 37752 6500 37776 6502
rect 37832 6500 37856 6502
rect 37912 6500 37918 6502
rect 37610 6491 37918 6500
rect 37610 5468 37918 5477
rect 37610 5466 37616 5468
rect 37672 5466 37696 5468
rect 37752 5466 37776 5468
rect 37832 5466 37856 5468
rect 37912 5466 37918 5468
rect 37672 5414 37674 5466
rect 37854 5414 37856 5466
rect 37610 5412 37616 5414
rect 37672 5412 37696 5414
rect 37752 5412 37776 5414
rect 37832 5412 37856 5414
rect 37912 5412 37918 5414
rect 37610 5403 37918 5412
rect 37464 5024 37516 5030
rect 37464 4966 37516 4972
rect 38120 4690 38148 16546
rect 38200 15496 38252 15502
rect 38200 15438 38252 15444
rect 38212 14822 38240 15438
rect 38304 15026 38332 24686
rect 38396 15366 38424 25230
rect 38568 24812 38620 24818
rect 38568 24754 38620 24760
rect 38476 21412 38528 21418
rect 38476 21354 38528 21360
rect 38384 15360 38436 15366
rect 38384 15302 38436 15308
rect 38488 15178 38516 21354
rect 38580 15502 38608 24754
rect 38568 15496 38620 15502
rect 38568 15438 38620 15444
rect 38568 15360 38620 15366
rect 38568 15302 38620 15308
rect 38396 15150 38516 15178
rect 38292 15020 38344 15026
rect 38292 14962 38344 14968
rect 38200 14816 38252 14822
rect 38200 14758 38252 14764
rect 38396 13938 38424 15150
rect 38384 13932 38436 13938
rect 38384 13874 38436 13880
rect 38580 13190 38608 15302
rect 38672 15094 38700 40326
rect 38660 15088 38712 15094
rect 38660 15030 38712 15036
rect 38764 14074 38792 44950
rect 38856 37262 38884 47738
rect 38844 37256 38896 37262
rect 38844 37198 38896 37204
rect 38948 35222 38976 57394
rect 39224 53514 39252 57394
rect 39316 55962 39344 58550
rect 39592 57458 39620 66166
rect 39948 59628 40000 59634
rect 39948 59570 40000 59576
rect 39672 59560 39724 59566
rect 39672 59502 39724 59508
rect 39580 57452 39632 57458
rect 39580 57394 39632 57400
rect 39304 55956 39356 55962
rect 39304 55898 39356 55904
rect 39212 53508 39264 53514
rect 39212 53450 39264 53456
rect 39028 37256 39080 37262
rect 39028 37198 39080 37204
rect 38936 35216 38988 35222
rect 38936 35158 38988 35164
rect 38936 29708 38988 29714
rect 38936 29650 38988 29656
rect 38948 29306 38976 29650
rect 38936 29300 38988 29306
rect 38936 29242 38988 29248
rect 38936 25764 38988 25770
rect 38936 25706 38988 25712
rect 38844 22568 38896 22574
rect 38844 22510 38896 22516
rect 38856 22098 38884 22510
rect 38844 22092 38896 22098
rect 38844 22034 38896 22040
rect 38752 14068 38804 14074
rect 38752 14010 38804 14016
rect 38764 13530 38792 14010
rect 38856 13938 38884 22034
rect 38948 17678 38976 25706
rect 39040 21486 39068 37198
rect 39224 24818 39252 53450
rect 39684 50386 39712 59502
rect 39960 58313 39988 59570
rect 39946 58304 40002 58313
rect 39946 58239 40002 58248
rect 39856 57452 39908 57458
rect 39856 57394 39908 57400
rect 39868 56982 39896 57394
rect 39856 56976 39908 56982
rect 39856 56918 39908 56924
rect 39672 50380 39724 50386
rect 39672 50322 39724 50328
rect 40500 49836 40552 49842
rect 40500 49778 40552 49784
rect 40512 49337 40540 49778
rect 40498 49328 40554 49337
rect 40498 49263 40554 49272
rect 39488 46436 39540 46442
rect 39488 46378 39540 46384
rect 39304 40588 39356 40594
rect 39304 40530 39356 40536
rect 39316 40118 39344 40530
rect 39304 40112 39356 40118
rect 39304 40054 39356 40060
rect 39212 24812 39264 24818
rect 39212 24754 39264 24760
rect 39028 21480 39080 21486
rect 39028 21422 39080 21428
rect 38936 17672 38988 17678
rect 38936 17614 38988 17620
rect 39304 15904 39356 15910
rect 39304 15846 39356 15852
rect 39028 14884 39080 14890
rect 39028 14826 39080 14832
rect 38844 13932 38896 13938
rect 38844 13874 38896 13880
rect 38752 13524 38804 13530
rect 38752 13466 38804 13472
rect 38568 13184 38620 13190
rect 38568 13126 38620 13132
rect 38764 12986 38792 13466
rect 39040 13326 39068 14826
rect 39316 14414 39344 15846
rect 39500 14482 39528 46378
rect 40866 40352 40922 40361
rect 40866 40287 40922 40296
rect 40880 40118 40908 40287
rect 40868 40112 40920 40118
rect 40868 40054 40920 40060
rect 40498 31376 40554 31385
rect 40498 31311 40500 31320
rect 40552 31311 40554 31320
rect 40500 31282 40552 31288
rect 40500 22636 40552 22642
rect 40500 22578 40552 22584
rect 40512 22409 40540 22578
rect 40498 22400 40554 22409
rect 40498 22335 40554 22344
rect 39488 14476 39540 14482
rect 39488 14418 39540 14424
rect 39304 14408 39356 14414
rect 39304 14350 39356 14356
rect 39948 13932 40000 13938
rect 39948 13874 40000 13880
rect 39960 13433 39988 13874
rect 39946 13424 40002 13433
rect 39946 13359 40002 13368
rect 39028 13320 39080 13326
rect 39028 13262 39080 13268
rect 38752 12980 38804 12986
rect 38752 12922 38804 12928
rect 38568 5024 38620 5030
rect 38568 4966 38620 4972
rect 38580 4758 38608 4966
rect 38568 4752 38620 4758
rect 38568 4694 38620 4700
rect 37372 4684 37424 4690
rect 37372 4626 37424 4632
rect 38108 4684 38160 4690
rect 38108 4626 38160 4632
rect 37280 4548 37332 4554
rect 37280 4490 37332 4496
rect 40498 4448 40554 4457
rect 37610 4380 37918 4389
rect 40498 4383 40554 4392
rect 37610 4378 37616 4380
rect 37672 4378 37696 4380
rect 37752 4378 37776 4380
rect 37832 4378 37856 4380
rect 37912 4378 37918 4380
rect 37672 4326 37674 4378
rect 37854 4326 37856 4378
rect 37610 4324 37616 4326
rect 37672 4324 37696 4326
rect 37752 4324 37776 4326
rect 37832 4324 37856 4326
rect 37912 4324 37918 4326
rect 37610 4315 37918 4324
rect 40512 4214 40540 4383
rect 40500 4208 40552 4214
rect 40500 4150 40552 4156
rect 36820 4072 36872 4078
rect 36820 4014 36872 4020
rect 36832 3602 36860 4014
rect 36950 3836 37258 3845
rect 36950 3834 36956 3836
rect 37012 3834 37036 3836
rect 37092 3834 37116 3836
rect 37172 3834 37196 3836
rect 37252 3834 37258 3836
rect 37012 3782 37014 3834
rect 37194 3782 37196 3834
rect 36950 3780 36956 3782
rect 37012 3780 37036 3782
rect 37092 3780 37116 3782
rect 37172 3780 37196 3782
rect 37252 3780 37258 3782
rect 36950 3771 37258 3780
rect 35900 3596 35952 3602
rect 35900 3538 35952 3544
rect 36820 3596 36872 3602
rect 36820 3538 36872 3544
rect 37610 3292 37918 3301
rect 37610 3290 37616 3292
rect 37672 3290 37696 3292
rect 37752 3290 37776 3292
rect 37832 3290 37856 3292
rect 37912 3290 37918 3292
rect 37672 3238 37674 3290
rect 37854 3238 37856 3290
rect 37610 3236 37616 3238
rect 37672 3236 37696 3238
rect 37752 3236 37776 3238
rect 37832 3236 37856 3238
rect 37912 3236 37918 3238
rect 37610 3227 37918 3236
rect 36950 2748 37258 2757
rect 36950 2746 36956 2748
rect 37012 2746 37036 2748
rect 37092 2746 37116 2748
rect 37172 2746 37196 2748
rect 37252 2746 37258 2748
rect 37012 2694 37014 2746
rect 37194 2694 37196 2746
rect 36950 2692 36956 2694
rect 37012 2692 37036 2694
rect 37092 2692 37116 2694
rect 37172 2692 37196 2694
rect 37252 2692 37258 2694
rect 36950 2683 37258 2692
rect 34612 2508 34664 2514
rect 34612 2450 34664 2456
rect 10140 2440 10192 2446
rect 34152 2440 34204 2446
rect 10140 2382 10192 2388
rect 28630 2408 28686 2417
rect 8024 2372 8076 2378
rect 34152 2382 34204 2388
rect 28630 2343 28632 2352
rect 8024 2314 8076 2320
rect 28684 2343 28686 2352
rect 28632 2314 28684 2320
rect 2610 2204 2918 2213
rect 2610 2202 2616 2204
rect 2672 2202 2696 2204
rect 2752 2202 2776 2204
rect 2832 2202 2856 2204
rect 2912 2202 2918 2204
rect 2672 2150 2674 2202
rect 2854 2150 2856 2202
rect 2610 2148 2616 2150
rect 2672 2148 2696 2150
rect 2752 2148 2776 2150
rect 2832 2148 2856 2150
rect 2912 2148 2918 2150
rect 2610 2139 2918 2148
rect 7610 2204 7918 2213
rect 7610 2202 7616 2204
rect 7672 2202 7696 2204
rect 7752 2202 7776 2204
rect 7832 2202 7856 2204
rect 7912 2202 7918 2204
rect 7672 2150 7674 2202
rect 7854 2150 7856 2202
rect 7610 2148 7616 2150
rect 7672 2148 7696 2150
rect 7752 2148 7776 2150
rect 7832 2148 7856 2150
rect 7912 2148 7918 2150
rect 7610 2139 7918 2148
rect 8036 1170 8064 2314
rect 13084 2304 13136 2310
rect 13084 2246 13136 2252
rect 18328 2304 18380 2310
rect 18328 2246 18380 2252
rect 23572 2304 23624 2310
rect 23572 2246 23624 2252
rect 28816 2304 28868 2310
rect 28816 2246 28868 2252
rect 34060 2304 34112 2310
rect 34060 2246 34112 2252
rect 39304 2304 39356 2310
rect 39304 2246 39356 2252
rect 12610 2204 12918 2213
rect 12610 2202 12616 2204
rect 12672 2202 12696 2204
rect 12752 2202 12776 2204
rect 12832 2202 12856 2204
rect 12912 2202 12918 2204
rect 12672 2150 12674 2202
rect 12854 2150 12856 2202
rect 12610 2148 12616 2150
rect 12672 2148 12696 2150
rect 12752 2148 12776 2150
rect 12832 2148 12856 2150
rect 12912 2148 12918 2150
rect 12610 2139 12918 2148
rect 2516 1142 2636 1170
rect 2608 800 2636 1142
rect 7852 1142 8064 1170
rect 7852 800 7880 1142
rect 13096 800 13124 2246
rect 17610 2204 17918 2213
rect 17610 2202 17616 2204
rect 17672 2202 17696 2204
rect 17752 2202 17776 2204
rect 17832 2202 17856 2204
rect 17912 2202 17918 2204
rect 17672 2150 17674 2202
rect 17854 2150 17856 2202
rect 17610 2148 17616 2150
rect 17672 2148 17696 2150
rect 17752 2148 17776 2150
rect 17832 2148 17856 2150
rect 17912 2148 17918 2150
rect 17610 2139 17918 2148
rect 18340 800 18368 2246
rect 22610 2204 22918 2213
rect 22610 2202 22616 2204
rect 22672 2202 22696 2204
rect 22752 2202 22776 2204
rect 22832 2202 22856 2204
rect 22912 2202 22918 2204
rect 22672 2150 22674 2202
rect 22854 2150 22856 2202
rect 22610 2148 22616 2150
rect 22672 2148 22696 2150
rect 22752 2148 22776 2150
rect 22832 2148 22856 2150
rect 22912 2148 22918 2150
rect 22610 2139 22918 2148
rect 23584 800 23612 2246
rect 27610 2204 27918 2213
rect 27610 2202 27616 2204
rect 27672 2202 27696 2204
rect 27752 2202 27776 2204
rect 27832 2202 27856 2204
rect 27912 2202 27918 2204
rect 27672 2150 27674 2202
rect 27854 2150 27856 2202
rect 27610 2148 27616 2150
rect 27672 2148 27696 2150
rect 27752 2148 27776 2150
rect 27832 2148 27856 2150
rect 27912 2148 27918 2150
rect 27610 2139 27918 2148
rect 28828 800 28856 2246
rect 32610 2204 32918 2213
rect 32610 2202 32616 2204
rect 32672 2202 32696 2204
rect 32752 2202 32776 2204
rect 32832 2202 32856 2204
rect 32912 2202 32918 2204
rect 32672 2150 32674 2202
rect 32854 2150 32856 2202
rect 32610 2148 32616 2150
rect 32672 2148 32696 2150
rect 32752 2148 32776 2150
rect 32832 2148 32856 2150
rect 32912 2148 32918 2150
rect 32610 2139 32918 2148
rect 34072 800 34100 2246
rect 37610 2204 37918 2213
rect 37610 2202 37616 2204
rect 37672 2202 37696 2204
rect 37752 2202 37776 2204
rect 37832 2202 37856 2204
rect 37912 2202 37918 2204
rect 37672 2150 37674 2202
rect 37854 2150 37856 2202
rect 37610 2148 37616 2150
rect 37672 2148 37696 2150
rect 37752 2148 37776 2150
rect 37832 2148 37856 2150
rect 37912 2148 37918 2150
rect 37610 2139 37918 2148
rect 39316 800 39344 2246
rect 2594 0 2650 800
rect 7838 0 7894 800
rect 13082 0 13138 800
rect 18326 0 18382 800
rect 23570 0 23626 800
rect 28814 0 28870 800
rect 34058 0 34114 800
rect 39302 0 39358 800
<< via2 >>
rect 2616 69658 2672 69660
rect 2696 69658 2752 69660
rect 2776 69658 2832 69660
rect 2856 69658 2912 69660
rect 2616 69606 2662 69658
rect 2662 69606 2672 69658
rect 2696 69606 2726 69658
rect 2726 69606 2738 69658
rect 2738 69606 2752 69658
rect 2776 69606 2790 69658
rect 2790 69606 2802 69658
rect 2802 69606 2832 69658
rect 2856 69606 2866 69658
rect 2866 69606 2912 69658
rect 2616 69604 2672 69606
rect 2696 69604 2752 69606
rect 2776 69604 2832 69606
rect 2856 69604 2912 69606
rect 7616 69658 7672 69660
rect 7696 69658 7752 69660
rect 7776 69658 7832 69660
rect 7856 69658 7912 69660
rect 7616 69606 7662 69658
rect 7662 69606 7672 69658
rect 7696 69606 7726 69658
rect 7726 69606 7738 69658
rect 7738 69606 7752 69658
rect 7776 69606 7790 69658
rect 7790 69606 7802 69658
rect 7802 69606 7832 69658
rect 7856 69606 7866 69658
rect 7866 69606 7912 69658
rect 7616 69604 7672 69606
rect 7696 69604 7752 69606
rect 7776 69604 7832 69606
rect 7856 69604 7912 69606
rect 12616 69658 12672 69660
rect 12696 69658 12752 69660
rect 12776 69658 12832 69660
rect 12856 69658 12912 69660
rect 12616 69606 12662 69658
rect 12662 69606 12672 69658
rect 12696 69606 12726 69658
rect 12726 69606 12738 69658
rect 12738 69606 12752 69658
rect 12776 69606 12790 69658
rect 12790 69606 12802 69658
rect 12802 69606 12832 69658
rect 12856 69606 12866 69658
rect 12866 69606 12912 69658
rect 12616 69604 12672 69606
rect 12696 69604 12752 69606
rect 12776 69604 12832 69606
rect 12856 69604 12912 69606
rect 17616 69658 17672 69660
rect 17696 69658 17752 69660
rect 17776 69658 17832 69660
rect 17856 69658 17912 69660
rect 17616 69606 17662 69658
rect 17662 69606 17672 69658
rect 17696 69606 17726 69658
rect 17726 69606 17738 69658
rect 17738 69606 17752 69658
rect 17776 69606 17790 69658
rect 17790 69606 17802 69658
rect 17802 69606 17832 69658
rect 17856 69606 17866 69658
rect 17866 69606 17912 69658
rect 17616 69604 17672 69606
rect 17696 69604 17752 69606
rect 17776 69604 17832 69606
rect 17856 69604 17912 69606
rect 22616 69658 22672 69660
rect 22696 69658 22752 69660
rect 22776 69658 22832 69660
rect 22856 69658 22912 69660
rect 22616 69606 22662 69658
rect 22662 69606 22672 69658
rect 22696 69606 22726 69658
rect 22726 69606 22738 69658
rect 22738 69606 22752 69658
rect 22776 69606 22790 69658
rect 22790 69606 22802 69658
rect 22802 69606 22832 69658
rect 22856 69606 22866 69658
rect 22866 69606 22912 69658
rect 22616 69604 22672 69606
rect 22696 69604 22752 69606
rect 22776 69604 22832 69606
rect 22856 69604 22912 69606
rect 27616 69658 27672 69660
rect 27696 69658 27752 69660
rect 27776 69658 27832 69660
rect 27856 69658 27912 69660
rect 27616 69606 27662 69658
rect 27662 69606 27672 69658
rect 27696 69606 27726 69658
rect 27726 69606 27738 69658
rect 27738 69606 27752 69658
rect 27776 69606 27790 69658
rect 27790 69606 27802 69658
rect 27802 69606 27832 69658
rect 27856 69606 27866 69658
rect 27866 69606 27912 69658
rect 27616 69604 27672 69606
rect 27696 69604 27752 69606
rect 27776 69604 27832 69606
rect 27856 69604 27912 69606
rect 32616 69658 32672 69660
rect 32696 69658 32752 69660
rect 32776 69658 32832 69660
rect 32856 69658 32912 69660
rect 32616 69606 32662 69658
rect 32662 69606 32672 69658
rect 32696 69606 32726 69658
rect 32726 69606 32738 69658
rect 32738 69606 32752 69658
rect 32776 69606 32790 69658
rect 32790 69606 32802 69658
rect 32802 69606 32832 69658
rect 32856 69606 32866 69658
rect 32866 69606 32912 69658
rect 32616 69604 32672 69606
rect 32696 69604 32752 69606
rect 32776 69604 32832 69606
rect 32856 69604 32912 69606
rect 37616 69658 37672 69660
rect 37696 69658 37752 69660
rect 37776 69658 37832 69660
rect 37856 69658 37912 69660
rect 37616 69606 37662 69658
rect 37662 69606 37672 69658
rect 37696 69606 37726 69658
rect 37726 69606 37738 69658
rect 37738 69606 37752 69658
rect 37776 69606 37790 69658
rect 37790 69606 37802 69658
rect 37802 69606 37832 69658
rect 37856 69606 37866 69658
rect 37866 69606 37912 69658
rect 37616 69604 37672 69606
rect 37696 69604 37752 69606
rect 37776 69604 37832 69606
rect 37856 69604 37912 69606
rect 1956 69114 2012 69116
rect 2036 69114 2092 69116
rect 2116 69114 2172 69116
rect 2196 69114 2252 69116
rect 1956 69062 2002 69114
rect 2002 69062 2012 69114
rect 2036 69062 2066 69114
rect 2066 69062 2078 69114
rect 2078 69062 2092 69114
rect 2116 69062 2130 69114
rect 2130 69062 2142 69114
rect 2142 69062 2172 69114
rect 2196 69062 2206 69114
rect 2206 69062 2252 69114
rect 1956 69060 2012 69062
rect 2036 69060 2092 69062
rect 2116 69060 2172 69062
rect 2196 69060 2252 69062
rect 6956 69114 7012 69116
rect 7036 69114 7092 69116
rect 7116 69114 7172 69116
rect 7196 69114 7252 69116
rect 6956 69062 7002 69114
rect 7002 69062 7012 69114
rect 7036 69062 7066 69114
rect 7066 69062 7078 69114
rect 7078 69062 7092 69114
rect 7116 69062 7130 69114
rect 7130 69062 7142 69114
rect 7142 69062 7172 69114
rect 7196 69062 7206 69114
rect 7206 69062 7252 69114
rect 6956 69060 7012 69062
rect 7036 69060 7092 69062
rect 7116 69060 7172 69062
rect 7196 69060 7252 69062
rect 2616 68570 2672 68572
rect 2696 68570 2752 68572
rect 2776 68570 2832 68572
rect 2856 68570 2912 68572
rect 2616 68518 2662 68570
rect 2662 68518 2672 68570
rect 2696 68518 2726 68570
rect 2726 68518 2738 68570
rect 2738 68518 2752 68570
rect 2776 68518 2790 68570
rect 2790 68518 2802 68570
rect 2802 68518 2832 68570
rect 2856 68518 2866 68570
rect 2866 68518 2912 68570
rect 2616 68516 2672 68518
rect 2696 68516 2752 68518
rect 2776 68516 2832 68518
rect 2856 68516 2912 68518
rect 7616 68570 7672 68572
rect 7696 68570 7752 68572
rect 7776 68570 7832 68572
rect 7856 68570 7912 68572
rect 7616 68518 7662 68570
rect 7662 68518 7672 68570
rect 7696 68518 7726 68570
rect 7726 68518 7738 68570
rect 7738 68518 7752 68570
rect 7776 68518 7790 68570
rect 7790 68518 7802 68570
rect 7802 68518 7832 68570
rect 7856 68518 7866 68570
rect 7866 68518 7912 68570
rect 7616 68516 7672 68518
rect 7696 68516 7752 68518
rect 7776 68516 7832 68518
rect 7856 68516 7912 68518
rect 1956 68026 2012 68028
rect 2036 68026 2092 68028
rect 2116 68026 2172 68028
rect 2196 68026 2252 68028
rect 1956 67974 2002 68026
rect 2002 67974 2012 68026
rect 2036 67974 2066 68026
rect 2066 67974 2078 68026
rect 2078 67974 2092 68026
rect 2116 67974 2130 68026
rect 2130 67974 2142 68026
rect 2142 67974 2172 68026
rect 2196 67974 2206 68026
rect 2206 67974 2252 68026
rect 1956 67972 2012 67974
rect 2036 67972 2092 67974
rect 2116 67972 2172 67974
rect 2196 67972 2252 67974
rect 6956 68026 7012 68028
rect 7036 68026 7092 68028
rect 7116 68026 7172 68028
rect 7196 68026 7252 68028
rect 6956 67974 7002 68026
rect 7002 67974 7012 68026
rect 7036 67974 7066 68026
rect 7066 67974 7078 68026
rect 7078 67974 7092 68026
rect 7116 67974 7130 68026
rect 7130 67974 7142 68026
rect 7142 67974 7172 68026
rect 7196 67974 7206 68026
rect 7206 67974 7252 68026
rect 6956 67972 7012 67974
rect 7036 67972 7092 67974
rect 7116 67972 7172 67974
rect 7196 67972 7252 67974
rect 2616 67482 2672 67484
rect 2696 67482 2752 67484
rect 2776 67482 2832 67484
rect 2856 67482 2912 67484
rect 2616 67430 2662 67482
rect 2662 67430 2672 67482
rect 2696 67430 2726 67482
rect 2726 67430 2738 67482
rect 2738 67430 2752 67482
rect 2776 67430 2790 67482
rect 2790 67430 2802 67482
rect 2802 67430 2832 67482
rect 2856 67430 2866 67482
rect 2866 67430 2912 67482
rect 2616 67428 2672 67430
rect 2696 67428 2752 67430
rect 2776 67428 2832 67430
rect 2856 67428 2912 67430
rect 1398 67224 1454 67280
rect 1956 66938 2012 66940
rect 2036 66938 2092 66940
rect 2116 66938 2172 66940
rect 2196 66938 2252 66940
rect 1956 66886 2002 66938
rect 2002 66886 2012 66938
rect 2036 66886 2066 66938
rect 2066 66886 2078 66938
rect 2078 66886 2092 66938
rect 2116 66886 2130 66938
rect 2130 66886 2142 66938
rect 2142 66886 2172 66938
rect 2196 66886 2206 66938
rect 2206 66886 2252 66938
rect 1956 66884 2012 66886
rect 2036 66884 2092 66886
rect 2116 66884 2172 66886
rect 2196 66884 2252 66886
rect 2616 66394 2672 66396
rect 2696 66394 2752 66396
rect 2776 66394 2832 66396
rect 2856 66394 2912 66396
rect 2616 66342 2662 66394
rect 2662 66342 2672 66394
rect 2696 66342 2726 66394
rect 2726 66342 2738 66394
rect 2738 66342 2752 66394
rect 2776 66342 2790 66394
rect 2790 66342 2802 66394
rect 2802 66342 2832 66394
rect 2856 66342 2866 66394
rect 2866 66342 2912 66394
rect 2616 66340 2672 66342
rect 2696 66340 2752 66342
rect 2776 66340 2832 66342
rect 2856 66340 2912 66342
rect 1956 65850 2012 65852
rect 2036 65850 2092 65852
rect 2116 65850 2172 65852
rect 2196 65850 2252 65852
rect 1956 65798 2002 65850
rect 2002 65798 2012 65850
rect 2036 65798 2066 65850
rect 2066 65798 2078 65850
rect 2078 65798 2092 65850
rect 2116 65798 2130 65850
rect 2130 65798 2142 65850
rect 2142 65798 2172 65850
rect 2196 65798 2206 65850
rect 2206 65798 2252 65850
rect 1956 65796 2012 65798
rect 2036 65796 2092 65798
rect 2116 65796 2172 65798
rect 2196 65796 2252 65798
rect 846 58384 902 58440
rect 1398 49272 1454 49328
rect 846 40160 902 40216
rect 1398 31320 1454 31376
rect 846 22480 902 22536
rect 1398 13368 1454 13424
rect 2616 65306 2672 65308
rect 2696 65306 2752 65308
rect 2776 65306 2832 65308
rect 2856 65306 2912 65308
rect 2616 65254 2662 65306
rect 2662 65254 2672 65306
rect 2696 65254 2726 65306
rect 2726 65254 2738 65306
rect 2738 65254 2752 65306
rect 2776 65254 2790 65306
rect 2790 65254 2802 65306
rect 2802 65254 2832 65306
rect 2856 65254 2866 65306
rect 2866 65254 2912 65306
rect 2616 65252 2672 65254
rect 2696 65252 2752 65254
rect 2776 65252 2832 65254
rect 2856 65252 2912 65254
rect 1956 64762 2012 64764
rect 2036 64762 2092 64764
rect 2116 64762 2172 64764
rect 2196 64762 2252 64764
rect 1956 64710 2002 64762
rect 2002 64710 2012 64762
rect 2036 64710 2066 64762
rect 2066 64710 2078 64762
rect 2078 64710 2092 64762
rect 2116 64710 2130 64762
rect 2130 64710 2142 64762
rect 2142 64710 2172 64762
rect 2196 64710 2206 64762
rect 2206 64710 2252 64762
rect 1956 64708 2012 64710
rect 2036 64708 2092 64710
rect 2116 64708 2172 64710
rect 2196 64708 2252 64710
rect 2616 64218 2672 64220
rect 2696 64218 2752 64220
rect 2776 64218 2832 64220
rect 2856 64218 2912 64220
rect 2616 64166 2662 64218
rect 2662 64166 2672 64218
rect 2696 64166 2726 64218
rect 2726 64166 2738 64218
rect 2738 64166 2752 64218
rect 2776 64166 2790 64218
rect 2790 64166 2802 64218
rect 2802 64166 2832 64218
rect 2856 64166 2866 64218
rect 2866 64166 2912 64218
rect 2616 64164 2672 64166
rect 2696 64164 2752 64166
rect 2776 64164 2832 64166
rect 2856 64164 2912 64166
rect 1956 63674 2012 63676
rect 2036 63674 2092 63676
rect 2116 63674 2172 63676
rect 2196 63674 2252 63676
rect 1956 63622 2002 63674
rect 2002 63622 2012 63674
rect 2036 63622 2066 63674
rect 2066 63622 2078 63674
rect 2078 63622 2092 63674
rect 2116 63622 2130 63674
rect 2130 63622 2142 63674
rect 2142 63622 2172 63674
rect 2196 63622 2206 63674
rect 2206 63622 2252 63674
rect 1956 63620 2012 63622
rect 2036 63620 2092 63622
rect 2116 63620 2172 63622
rect 2196 63620 2252 63622
rect 2616 63130 2672 63132
rect 2696 63130 2752 63132
rect 2776 63130 2832 63132
rect 2856 63130 2912 63132
rect 2616 63078 2662 63130
rect 2662 63078 2672 63130
rect 2696 63078 2726 63130
rect 2726 63078 2738 63130
rect 2738 63078 2752 63130
rect 2776 63078 2790 63130
rect 2790 63078 2802 63130
rect 2802 63078 2832 63130
rect 2856 63078 2866 63130
rect 2866 63078 2912 63130
rect 2616 63076 2672 63078
rect 2696 63076 2752 63078
rect 2776 63076 2832 63078
rect 2856 63076 2912 63078
rect 1956 62586 2012 62588
rect 2036 62586 2092 62588
rect 2116 62586 2172 62588
rect 2196 62586 2252 62588
rect 1956 62534 2002 62586
rect 2002 62534 2012 62586
rect 2036 62534 2066 62586
rect 2066 62534 2078 62586
rect 2078 62534 2092 62586
rect 2116 62534 2130 62586
rect 2130 62534 2142 62586
rect 2142 62534 2172 62586
rect 2196 62534 2206 62586
rect 2206 62534 2252 62586
rect 1956 62532 2012 62534
rect 2036 62532 2092 62534
rect 2116 62532 2172 62534
rect 2196 62532 2252 62534
rect 2616 62042 2672 62044
rect 2696 62042 2752 62044
rect 2776 62042 2832 62044
rect 2856 62042 2912 62044
rect 2616 61990 2662 62042
rect 2662 61990 2672 62042
rect 2696 61990 2726 62042
rect 2726 61990 2738 62042
rect 2738 61990 2752 62042
rect 2776 61990 2790 62042
rect 2790 61990 2802 62042
rect 2802 61990 2832 62042
rect 2856 61990 2866 62042
rect 2866 61990 2912 62042
rect 2616 61988 2672 61990
rect 2696 61988 2752 61990
rect 2776 61988 2832 61990
rect 2856 61988 2912 61990
rect 1956 61498 2012 61500
rect 2036 61498 2092 61500
rect 2116 61498 2172 61500
rect 2196 61498 2252 61500
rect 1956 61446 2002 61498
rect 2002 61446 2012 61498
rect 2036 61446 2066 61498
rect 2066 61446 2078 61498
rect 2078 61446 2092 61498
rect 2116 61446 2130 61498
rect 2130 61446 2142 61498
rect 2142 61446 2172 61498
rect 2196 61446 2206 61498
rect 2206 61446 2252 61498
rect 1956 61444 2012 61446
rect 2036 61444 2092 61446
rect 2116 61444 2172 61446
rect 2196 61444 2252 61446
rect 1956 60410 2012 60412
rect 2036 60410 2092 60412
rect 2116 60410 2172 60412
rect 2196 60410 2252 60412
rect 1956 60358 2002 60410
rect 2002 60358 2012 60410
rect 2036 60358 2066 60410
rect 2066 60358 2078 60410
rect 2078 60358 2092 60410
rect 2116 60358 2130 60410
rect 2130 60358 2142 60410
rect 2142 60358 2172 60410
rect 2196 60358 2206 60410
rect 2206 60358 2252 60410
rect 1956 60356 2012 60358
rect 2036 60356 2092 60358
rect 2116 60356 2172 60358
rect 2196 60356 2252 60358
rect 1956 59322 2012 59324
rect 2036 59322 2092 59324
rect 2116 59322 2172 59324
rect 2196 59322 2252 59324
rect 1956 59270 2002 59322
rect 2002 59270 2012 59322
rect 2036 59270 2066 59322
rect 2066 59270 2078 59322
rect 2078 59270 2092 59322
rect 2116 59270 2130 59322
rect 2130 59270 2142 59322
rect 2142 59270 2172 59322
rect 2196 59270 2206 59322
rect 2206 59270 2252 59322
rect 1956 59268 2012 59270
rect 2036 59268 2092 59270
rect 2116 59268 2172 59270
rect 2196 59268 2252 59270
rect 1956 58234 2012 58236
rect 2036 58234 2092 58236
rect 2116 58234 2172 58236
rect 2196 58234 2252 58236
rect 1956 58182 2002 58234
rect 2002 58182 2012 58234
rect 2036 58182 2066 58234
rect 2066 58182 2078 58234
rect 2078 58182 2092 58234
rect 2116 58182 2130 58234
rect 2130 58182 2142 58234
rect 2142 58182 2172 58234
rect 2196 58182 2206 58234
rect 2206 58182 2252 58234
rect 1956 58180 2012 58182
rect 2036 58180 2092 58182
rect 2116 58180 2172 58182
rect 2196 58180 2252 58182
rect 1956 57146 2012 57148
rect 2036 57146 2092 57148
rect 2116 57146 2172 57148
rect 2196 57146 2252 57148
rect 1956 57094 2002 57146
rect 2002 57094 2012 57146
rect 2036 57094 2066 57146
rect 2066 57094 2078 57146
rect 2078 57094 2092 57146
rect 2116 57094 2130 57146
rect 2130 57094 2142 57146
rect 2142 57094 2172 57146
rect 2196 57094 2206 57146
rect 2206 57094 2252 57146
rect 1956 57092 2012 57094
rect 2036 57092 2092 57094
rect 2116 57092 2172 57094
rect 2196 57092 2252 57094
rect 1956 56058 2012 56060
rect 2036 56058 2092 56060
rect 2116 56058 2172 56060
rect 2196 56058 2252 56060
rect 1956 56006 2002 56058
rect 2002 56006 2012 56058
rect 2036 56006 2066 56058
rect 2066 56006 2078 56058
rect 2078 56006 2092 56058
rect 2116 56006 2130 56058
rect 2130 56006 2142 56058
rect 2142 56006 2172 56058
rect 2196 56006 2206 56058
rect 2206 56006 2252 56058
rect 1956 56004 2012 56006
rect 2036 56004 2092 56006
rect 2116 56004 2172 56006
rect 2196 56004 2252 56006
rect 1956 54970 2012 54972
rect 2036 54970 2092 54972
rect 2116 54970 2172 54972
rect 2196 54970 2252 54972
rect 1956 54918 2002 54970
rect 2002 54918 2012 54970
rect 2036 54918 2066 54970
rect 2066 54918 2078 54970
rect 2078 54918 2092 54970
rect 2116 54918 2130 54970
rect 2130 54918 2142 54970
rect 2142 54918 2172 54970
rect 2196 54918 2206 54970
rect 2206 54918 2252 54970
rect 1956 54916 2012 54918
rect 2036 54916 2092 54918
rect 2116 54916 2172 54918
rect 2196 54916 2252 54918
rect 1956 53882 2012 53884
rect 2036 53882 2092 53884
rect 2116 53882 2172 53884
rect 2196 53882 2252 53884
rect 1956 53830 2002 53882
rect 2002 53830 2012 53882
rect 2036 53830 2066 53882
rect 2066 53830 2078 53882
rect 2078 53830 2092 53882
rect 2116 53830 2130 53882
rect 2130 53830 2142 53882
rect 2142 53830 2172 53882
rect 2196 53830 2206 53882
rect 2206 53830 2252 53882
rect 1956 53828 2012 53830
rect 2036 53828 2092 53830
rect 2116 53828 2172 53830
rect 2196 53828 2252 53830
rect 2616 60954 2672 60956
rect 2696 60954 2752 60956
rect 2776 60954 2832 60956
rect 2856 60954 2912 60956
rect 2616 60902 2662 60954
rect 2662 60902 2672 60954
rect 2696 60902 2726 60954
rect 2726 60902 2738 60954
rect 2738 60902 2752 60954
rect 2776 60902 2790 60954
rect 2790 60902 2802 60954
rect 2802 60902 2832 60954
rect 2856 60902 2866 60954
rect 2866 60902 2912 60954
rect 2616 60900 2672 60902
rect 2696 60900 2752 60902
rect 2776 60900 2832 60902
rect 2856 60900 2912 60902
rect 2616 59866 2672 59868
rect 2696 59866 2752 59868
rect 2776 59866 2832 59868
rect 2856 59866 2912 59868
rect 2616 59814 2662 59866
rect 2662 59814 2672 59866
rect 2696 59814 2726 59866
rect 2726 59814 2738 59866
rect 2738 59814 2752 59866
rect 2776 59814 2790 59866
rect 2790 59814 2802 59866
rect 2802 59814 2832 59866
rect 2856 59814 2866 59866
rect 2866 59814 2912 59866
rect 2616 59812 2672 59814
rect 2696 59812 2752 59814
rect 2776 59812 2832 59814
rect 2856 59812 2912 59814
rect 2616 58778 2672 58780
rect 2696 58778 2752 58780
rect 2776 58778 2832 58780
rect 2856 58778 2912 58780
rect 2616 58726 2662 58778
rect 2662 58726 2672 58778
rect 2696 58726 2726 58778
rect 2726 58726 2738 58778
rect 2738 58726 2752 58778
rect 2776 58726 2790 58778
rect 2790 58726 2802 58778
rect 2802 58726 2832 58778
rect 2856 58726 2866 58778
rect 2866 58726 2912 58778
rect 2616 58724 2672 58726
rect 2696 58724 2752 58726
rect 2776 58724 2832 58726
rect 2856 58724 2912 58726
rect 2616 57690 2672 57692
rect 2696 57690 2752 57692
rect 2776 57690 2832 57692
rect 2856 57690 2912 57692
rect 2616 57638 2662 57690
rect 2662 57638 2672 57690
rect 2696 57638 2726 57690
rect 2726 57638 2738 57690
rect 2738 57638 2752 57690
rect 2776 57638 2790 57690
rect 2790 57638 2802 57690
rect 2802 57638 2832 57690
rect 2856 57638 2866 57690
rect 2866 57638 2912 57690
rect 2616 57636 2672 57638
rect 2696 57636 2752 57638
rect 2776 57636 2832 57638
rect 2856 57636 2912 57638
rect 2616 56602 2672 56604
rect 2696 56602 2752 56604
rect 2776 56602 2832 56604
rect 2856 56602 2912 56604
rect 2616 56550 2662 56602
rect 2662 56550 2672 56602
rect 2696 56550 2726 56602
rect 2726 56550 2738 56602
rect 2738 56550 2752 56602
rect 2776 56550 2790 56602
rect 2790 56550 2802 56602
rect 2802 56550 2832 56602
rect 2856 56550 2866 56602
rect 2866 56550 2912 56602
rect 2616 56548 2672 56550
rect 2696 56548 2752 56550
rect 2776 56548 2832 56550
rect 2856 56548 2912 56550
rect 2616 55514 2672 55516
rect 2696 55514 2752 55516
rect 2776 55514 2832 55516
rect 2856 55514 2912 55516
rect 2616 55462 2662 55514
rect 2662 55462 2672 55514
rect 2696 55462 2726 55514
rect 2726 55462 2738 55514
rect 2738 55462 2752 55514
rect 2776 55462 2790 55514
rect 2790 55462 2802 55514
rect 2802 55462 2832 55514
rect 2856 55462 2866 55514
rect 2866 55462 2912 55514
rect 2616 55460 2672 55462
rect 2696 55460 2752 55462
rect 2776 55460 2832 55462
rect 2856 55460 2912 55462
rect 2616 54426 2672 54428
rect 2696 54426 2752 54428
rect 2776 54426 2832 54428
rect 2856 54426 2912 54428
rect 2616 54374 2662 54426
rect 2662 54374 2672 54426
rect 2696 54374 2726 54426
rect 2726 54374 2738 54426
rect 2738 54374 2752 54426
rect 2776 54374 2790 54426
rect 2790 54374 2802 54426
rect 2802 54374 2832 54426
rect 2856 54374 2866 54426
rect 2866 54374 2912 54426
rect 2616 54372 2672 54374
rect 2696 54372 2752 54374
rect 2776 54372 2832 54374
rect 2856 54372 2912 54374
rect 2616 53338 2672 53340
rect 2696 53338 2752 53340
rect 2776 53338 2832 53340
rect 2856 53338 2912 53340
rect 2616 53286 2662 53338
rect 2662 53286 2672 53338
rect 2696 53286 2726 53338
rect 2726 53286 2738 53338
rect 2738 53286 2752 53338
rect 2776 53286 2790 53338
rect 2790 53286 2802 53338
rect 2802 53286 2832 53338
rect 2856 53286 2866 53338
rect 2866 53286 2912 53338
rect 2616 53284 2672 53286
rect 2696 53284 2752 53286
rect 2776 53284 2832 53286
rect 2856 53284 2912 53286
rect 1956 52794 2012 52796
rect 2036 52794 2092 52796
rect 2116 52794 2172 52796
rect 2196 52794 2252 52796
rect 1956 52742 2002 52794
rect 2002 52742 2012 52794
rect 2036 52742 2066 52794
rect 2066 52742 2078 52794
rect 2078 52742 2092 52794
rect 2116 52742 2130 52794
rect 2130 52742 2142 52794
rect 2142 52742 2172 52794
rect 2196 52742 2206 52794
rect 2206 52742 2252 52794
rect 1956 52740 2012 52742
rect 2036 52740 2092 52742
rect 2116 52740 2172 52742
rect 2196 52740 2252 52742
rect 2616 52250 2672 52252
rect 2696 52250 2752 52252
rect 2776 52250 2832 52252
rect 2856 52250 2912 52252
rect 2616 52198 2662 52250
rect 2662 52198 2672 52250
rect 2696 52198 2726 52250
rect 2726 52198 2738 52250
rect 2738 52198 2752 52250
rect 2776 52198 2790 52250
rect 2790 52198 2802 52250
rect 2802 52198 2832 52250
rect 2856 52198 2866 52250
rect 2866 52198 2912 52250
rect 2616 52196 2672 52198
rect 2696 52196 2752 52198
rect 2776 52196 2832 52198
rect 2856 52196 2912 52198
rect 1956 51706 2012 51708
rect 2036 51706 2092 51708
rect 2116 51706 2172 51708
rect 2196 51706 2252 51708
rect 1956 51654 2002 51706
rect 2002 51654 2012 51706
rect 2036 51654 2066 51706
rect 2066 51654 2078 51706
rect 2078 51654 2092 51706
rect 2116 51654 2130 51706
rect 2130 51654 2142 51706
rect 2142 51654 2172 51706
rect 2196 51654 2206 51706
rect 2206 51654 2252 51706
rect 1956 51652 2012 51654
rect 2036 51652 2092 51654
rect 2116 51652 2172 51654
rect 2196 51652 2252 51654
rect 2616 51162 2672 51164
rect 2696 51162 2752 51164
rect 2776 51162 2832 51164
rect 2856 51162 2912 51164
rect 2616 51110 2662 51162
rect 2662 51110 2672 51162
rect 2696 51110 2726 51162
rect 2726 51110 2738 51162
rect 2738 51110 2752 51162
rect 2776 51110 2790 51162
rect 2790 51110 2802 51162
rect 2802 51110 2832 51162
rect 2856 51110 2866 51162
rect 2866 51110 2912 51162
rect 2616 51108 2672 51110
rect 2696 51108 2752 51110
rect 2776 51108 2832 51110
rect 2856 51108 2912 51110
rect 1956 50618 2012 50620
rect 2036 50618 2092 50620
rect 2116 50618 2172 50620
rect 2196 50618 2252 50620
rect 1956 50566 2002 50618
rect 2002 50566 2012 50618
rect 2036 50566 2066 50618
rect 2066 50566 2078 50618
rect 2078 50566 2092 50618
rect 2116 50566 2130 50618
rect 2130 50566 2142 50618
rect 2142 50566 2172 50618
rect 2196 50566 2206 50618
rect 2206 50566 2252 50618
rect 1956 50564 2012 50566
rect 2036 50564 2092 50566
rect 2116 50564 2172 50566
rect 2196 50564 2252 50566
rect 2616 50074 2672 50076
rect 2696 50074 2752 50076
rect 2776 50074 2832 50076
rect 2856 50074 2912 50076
rect 2616 50022 2662 50074
rect 2662 50022 2672 50074
rect 2696 50022 2726 50074
rect 2726 50022 2738 50074
rect 2738 50022 2752 50074
rect 2776 50022 2790 50074
rect 2790 50022 2802 50074
rect 2802 50022 2832 50074
rect 2856 50022 2866 50074
rect 2866 50022 2912 50074
rect 2616 50020 2672 50022
rect 2696 50020 2752 50022
rect 2776 50020 2832 50022
rect 2856 50020 2912 50022
rect 1956 49530 2012 49532
rect 2036 49530 2092 49532
rect 2116 49530 2172 49532
rect 2196 49530 2252 49532
rect 1956 49478 2002 49530
rect 2002 49478 2012 49530
rect 2036 49478 2066 49530
rect 2066 49478 2078 49530
rect 2078 49478 2092 49530
rect 2116 49478 2130 49530
rect 2130 49478 2142 49530
rect 2142 49478 2172 49530
rect 2196 49478 2206 49530
rect 2206 49478 2252 49530
rect 1956 49476 2012 49478
rect 2036 49476 2092 49478
rect 2116 49476 2172 49478
rect 2196 49476 2252 49478
rect 2616 48986 2672 48988
rect 2696 48986 2752 48988
rect 2776 48986 2832 48988
rect 2856 48986 2912 48988
rect 2616 48934 2662 48986
rect 2662 48934 2672 48986
rect 2696 48934 2726 48986
rect 2726 48934 2738 48986
rect 2738 48934 2752 48986
rect 2776 48934 2790 48986
rect 2790 48934 2802 48986
rect 2802 48934 2832 48986
rect 2856 48934 2866 48986
rect 2866 48934 2912 48986
rect 2616 48932 2672 48934
rect 2696 48932 2752 48934
rect 2776 48932 2832 48934
rect 2856 48932 2912 48934
rect 1956 48442 2012 48444
rect 2036 48442 2092 48444
rect 2116 48442 2172 48444
rect 2196 48442 2252 48444
rect 1956 48390 2002 48442
rect 2002 48390 2012 48442
rect 2036 48390 2066 48442
rect 2066 48390 2078 48442
rect 2078 48390 2092 48442
rect 2116 48390 2130 48442
rect 2130 48390 2142 48442
rect 2142 48390 2172 48442
rect 2196 48390 2206 48442
rect 2206 48390 2252 48442
rect 1956 48388 2012 48390
rect 2036 48388 2092 48390
rect 2116 48388 2172 48390
rect 2196 48388 2252 48390
rect 2616 47898 2672 47900
rect 2696 47898 2752 47900
rect 2776 47898 2832 47900
rect 2856 47898 2912 47900
rect 2616 47846 2662 47898
rect 2662 47846 2672 47898
rect 2696 47846 2726 47898
rect 2726 47846 2738 47898
rect 2738 47846 2752 47898
rect 2776 47846 2790 47898
rect 2790 47846 2802 47898
rect 2802 47846 2832 47898
rect 2856 47846 2866 47898
rect 2866 47846 2912 47898
rect 2616 47844 2672 47846
rect 2696 47844 2752 47846
rect 2776 47844 2832 47846
rect 2856 47844 2912 47846
rect 1956 47354 2012 47356
rect 2036 47354 2092 47356
rect 2116 47354 2172 47356
rect 2196 47354 2252 47356
rect 1956 47302 2002 47354
rect 2002 47302 2012 47354
rect 2036 47302 2066 47354
rect 2066 47302 2078 47354
rect 2078 47302 2092 47354
rect 2116 47302 2130 47354
rect 2130 47302 2142 47354
rect 2142 47302 2172 47354
rect 2196 47302 2206 47354
rect 2206 47302 2252 47354
rect 1956 47300 2012 47302
rect 2036 47300 2092 47302
rect 2116 47300 2172 47302
rect 2196 47300 2252 47302
rect 1956 46266 2012 46268
rect 2036 46266 2092 46268
rect 2116 46266 2172 46268
rect 2196 46266 2252 46268
rect 1956 46214 2002 46266
rect 2002 46214 2012 46266
rect 2036 46214 2066 46266
rect 2066 46214 2078 46266
rect 2078 46214 2092 46266
rect 2116 46214 2130 46266
rect 2130 46214 2142 46266
rect 2142 46214 2172 46266
rect 2196 46214 2206 46266
rect 2206 46214 2252 46266
rect 1956 46212 2012 46214
rect 2036 46212 2092 46214
rect 2116 46212 2172 46214
rect 2196 46212 2252 46214
rect 1956 45178 2012 45180
rect 2036 45178 2092 45180
rect 2116 45178 2172 45180
rect 2196 45178 2252 45180
rect 1956 45126 2002 45178
rect 2002 45126 2012 45178
rect 2036 45126 2066 45178
rect 2066 45126 2078 45178
rect 2078 45126 2092 45178
rect 2116 45126 2130 45178
rect 2130 45126 2142 45178
rect 2142 45126 2172 45178
rect 2196 45126 2206 45178
rect 2206 45126 2252 45178
rect 1956 45124 2012 45126
rect 2036 45124 2092 45126
rect 2116 45124 2172 45126
rect 2196 45124 2252 45126
rect 1956 44090 2012 44092
rect 2036 44090 2092 44092
rect 2116 44090 2172 44092
rect 2196 44090 2252 44092
rect 1956 44038 2002 44090
rect 2002 44038 2012 44090
rect 2036 44038 2066 44090
rect 2066 44038 2078 44090
rect 2078 44038 2092 44090
rect 2116 44038 2130 44090
rect 2130 44038 2142 44090
rect 2142 44038 2172 44090
rect 2196 44038 2206 44090
rect 2206 44038 2252 44090
rect 1956 44036 2012 44038
rect 2036 44036 2092 44038
rect 2116 44036 2172 44038
rect 2196 44036 2252 44038
rect 1956 43002 2012 43004
rect 2036 43002 2092 43004
rect 2116 43002 2172 43004
rect 2196 43002 2252 43004
rect 1956 42950 2002 43002
rect 2002 42950 2012 43002
rect 2036 42950 2066 43002
rect 2066 42950 2078 43002
rect 2078 42950 2092 43002
rect 2116 42950 2130 43002
rect 2130 42950 2142 43002
rect 2142 42950 2172 43002
rect 2196 42950 2206 43002
rect 2206 42950 2252 43002
rect 1956 42948 2012 42950
rect 2036 42948 2092 42950
rect 2116 42948 2172 42950
rect 2196 42948 2252 42950
rect 1956 41914 2012 41916
rect 2036 41914 2092 41916
rect 2116 41914 2172 41916
rect 2196 41914 2252 41916
rect 1956 41862 2002 41914
rect 2002 41862 2012 41914
rect 2036 41862 2066 41914
rect 2066 41862 2078 41914
rect 2078 41862 2092 41914
rect 2116 41862 2130 41914
rect 2130 41862 2142 41914
rect 2142 41862 2172 41914
rect 2196 41862 2206 41914
rect 2206 41862 2252 41914
rect 1956 41860 2012 41862
rect 2036 41860 2092 41862
rect 2116 41860 2172 41862
rect 2196 41860 2252 41862
rect 1956 40826 2012 40828
rect 2036 40826 2092 40828
rect 2116 40826 2172 40828
rect 2196 40826 2252 40828
rect 1956 40774 2002 40826
rect 2002 40774 2012 40826
rect 2036 40774 2066 40826
rect 2066 40774 2078 40826
rect 2078 40774 2092 40826
rect 2116 40774 2130 40826
rect 2130 40774 2142 40826
rect 2142 40774 2172 40826
rect 2196 40774 2206 40826
rect 2206 40774 2252 40826
rect 1956 40772 2012 40774
rect 2036 40772 2092 40774
rect 2116 40772 2172 40774
rect 2196 40772 2252 40774
rect 1956 39738 2012 39740
rect 2036 39738 2092 39740
rect 2116 39738 2172 39740
rect 2196 39738 2252 39740
rect 1956 39686 2002 39738
rect 2002 39686 2012 39738
rect 2036 39686 2066 39738
rect 2066 39686 2078 39738
rect 2078 39686 2092 39738
rect 2116 39686 2130 39738
rect 2130 39686 2142 39738
rect 2142 39686 2172 39738
rect 2196 39686 2206 39738
rect 2206 39686 2252 39738
rect 1956 39684 2012 39686
rect 2036 39684 2092 39686
rect 2116 39684 2172 39686
rect 2196 39684 2252 39686
rect 1956 38650 2012 38652
rect 2036 38650 2092 38652
rect 2116 38650 2172 38652
rect 2196 38650 2252 38652
rect 1956 38598 2002 38650
rect 2002 38598 2012 38650
rect 2036 38598 2066 38650
rect 2066 38598 2078 38650
rect 2078 38598 2092 38650
rect 2116 38598 2130 38650
rect 2130 38598 2142 38650
rect 2142 38598 2172 38650
rect 2196 38598 2206 38650
rect 2206 38598 2252 38650
rect 1956 38596 2012 38598
rect 2036 38596 2092 38598
rect 2116 38596 2172 38598
rect 2196 38596 2252 38598
rect 1956 37562 2012 37564
rect 2036 37562 2092 37564
rect 2116 37562 2172 37564
rect 2196 37562 2252 37564
rect 1956 37510 2002 37562
rect 2002 37510 2012 37562
rect 2036 37510 2066 37562
rect 2066 37510 2078 37562
rect 2078 37510 2092 37562
rect 2116 37510 2130 37562
rect 2130 37510 2142 37562
rect 2142 37510 2172 37562
rect 2196 37510 2206 37562
rect 2206 37510 2252 37562
rect 1956 37508 2012 37510
rect 2036 37508 2092 37510
rect 2116 37508 2172 37510
rect 2196 37508 2252 37510
rect 1956 36474 2012 36476
rect 2036 36474 2092 36476
rect 2116 36474 2172 36476
rect 2196 36474 2252 36476
rect 1956 36422 2002 36474
rect 2002 36422 2012 36474
rect 2036 36422 2066 36474
rect 2066 36422 2078 36474
rect 2078 36422 2092 36474
rect 2116 36422 2130 36474
rect 2130 36422 2142 36474
rect 2142 36422 2172 36474
rect 2196 36422 2206 36474
rect 2206 36422 2252 36474
rect 1956 36420 2012 36422
rect 2036 36420 2092 36422
rect 2116 36420 2172 36422
rect 2196 36420 2252 36422
rect 1956 35386 2012 35388
rect 2036 35386 2092 35388
rect 2116 35386 2172 35388
rect 2196 35386 2252 35388
rect 1956 35334 2002 35386
rect 2002 35334 2012 35386
rect 2036 35334 2066 35386
rect 2066 35334 2078 35386
rect 2078 35334 2092 35386
rect 2116 35334 2130 35386
rect 2130 35334 2142 35386
rect 2142 35334 2172 35386
rect 2196 35334 2206 35386
rect 2206 35334 2252 35386
rect 1956 35332 2012 35334
rect 2036 35332 2092 35334
rect 2116 35332 2172 35334
rect 2196 35332 2252 35334
rect 1956 34298 2012 34300
rect 2036 34298 2092 34300
rect 2116 34298 2172 34300
rect 2196 34298 2252 34300
rect 1956 34246 2002 34298
rect 2002 34246 2012 34298
rect 2036 34246 2066 34298
rect 2066 34246 2078 34298
rect 2078 34246 2092 34298
rect 2116 34246 2130 34298
rect 2130 34246 2142 34298
rect 2142 34246 2172 34298
rect 2196 34246 2206 34298
rect 2206 34246 2252 34298
rect 1956 34244 2012 34246
rect 2036 34244 2092 34246
rect 2116 34244 2172 34246
rect 2196 34244 2252 34246
rect 1956 33210 2012 33212
rect 2036 33210 2092 33212
rect 2116 33210 2172 33212
rect 2196 33210 2252 33212
rect 1956 33158 2002 33210
rect 2002 33158 2012 33210
rect 2036 33158 2066 33210
rect 2066 33158 2078 33210
rect 2078 33158 2092 33210
rect 2116 33158 2130 33210
rect 2130 33158 2142 33210
rect 2142 33158 2172 33210
rect 2196 33158 2206 33210
rect 2206 33158 2252 33210
rect 1956 33156 2012 33158
rect 2036 33156 2092 33158
rect 2116 33156 2172 33158
rect 2196 33156 2252 33158
rect 1956 32122 2012 32124
rect 2036 32122 2092 32124
rect 2116 32122 2172 32124
rect 2196 32122 2252 32124
rect 1956 32070 2002 32122
rect 2002 32070 2012 32122
rect 2036 32070 2066 32122
rect 2066 32070 2078 32122
rect 2078 32070 2092 32122
rect 2116 32070 2130 32122
rect 2130 32070 2142 32122
rect 2142 32070 2172 32122
rect 2196 32070 2206 32122
rect 2206 32070 2252 32122
rect 1956 32068 2012 32070
rect 2036 32068 2092 32070
rect 2116 32068 2172 32070
rect 2196 32068 2252 32070
rect 1956 31034 2012 31036
rect 2036 31034 2092 31036
rect 2116 31034 2172 31036
rect 2196 31034 2252 31036
rect 1956 30982 2002 31034
rect 2002 30982 2012 31034
rect 2036 30982 2066 31034
rect 2066 30982 2078 31034
rect 2078 30982 2092 31034
rect 2116 30982 2130 31034
rect 2130 30982 2142 31034
rect 2142 30982 2172 31034
rect 2196 30982 2206 31034
rect 2206 30982 2252 31034
rect 1956 30980 2012 30982
rect 2036 30980 2092 30982
rect 2116 30980 2172 30982
rect 2196 30980 2252 30982
rect 1956 29946 2012 29948
rect 2036 29946 2092 29948
rect 2116 29946 2172 29948
rect 2196 29946 2252 29948
rect 1956 29894 2002 29946
rect 2002 29894 2012 29946
rect 2036 29894 2066 29946
rect 2066 29894 2078 29946
rect 2078 29894 2092 29946
rect 2116 29894 2130 29946
rect 2130 29894 2142 29946
rect 2142 29894 2172 29946
rect 2196 29894 2206 29946
rect 2206 29894 2252 29946
rect 1956 29892 2012 29894
rect 2036 29892 2092 29894
rect 2116 29892 2172 29894
rect 2196 29892 2252 29894
rect 1956 28858 2012 28860
rect 2036 28858 2092 28860
rect 2116 28858 2172 28860
rect 2196 28858 2252 28860
rect 1956 28806 2002 28858
rect 2002 28806 2012 28858
rect 2036 28806 2066 28858
rect 2066 28806 2078 28858
rect 2078 28806 2092 28858
rect 2116 28806 2130 28858
rect 2130 28806 2142 28858
rect 2142 28806 2172 28858
rect 2196 28806 2206 28858
rect 2206 28806 2252 28858
rect 1956 28804 2012 28806
rect 2036 28804 2092 28806
rect 2116 28804 2172 28806
rect 2196 28804 2252 28806
rect 1956 27770 2012 27772
rect 2036 27770 2092 27772
rect 2116 27770 2172 27772
rect 2196 27770 2252 27772
rect 1956 27718 2002 27770
rect 2002 27718 2012 27770
rect 2036 27718 2066 27770
rect 2066 27718 2078 27770
rect 2078 27718 2092 27770
rect 2116 27718 2130 27770
rect 2130 27718 2142 27770
rect 2142 27718 2172 27770
rect 2196 27718 2206 27770
rect 2206 27718 2252 27770
rect 1956 27716 2012 27718
rect 2036 27716 2092 27718
rect 2116 27716 2172 27718
rect 2196 27716 2252 27718
rect 1956 26682 2012 26684
rect 2036 26682 2092 26684
rect 2116 26682 2172 26684
rect 2196 26682 2252 26684
rect 1956 26630 2002 26682
rect 2002 26630 2012 26682
rect 2036 26630 2066 26682
rect 2066 26630 2078 26682
rect 2078 26630 2092 26682
rect 2116 26630 2130 26682
rect 2130 26630 2142 26682
rect 2142 26630 2172 26682
rect 2196 26630 2206 26682
rect 2206 26630 2252 26682
rect 1956 26628 2012 26630
rect 2036 26628 2092 26630
rect 2116 26628 2172 26630
rect 2196 26628 2252 26630
rect 1956 25594 2012 25596
rect 2036 25594 2092 25596
rect 2116 25594 2172 25596
rect 2196 25594 2252 25596
rect 1956 25542 2002 25594
rect 2002 25542 2012 25594
rect 2036 25542 2066 25594
rect 2066 25542 2078 25594
rect 2078 25542 2092 25594
rect 2116 25542 2130 25594
rect 2130 25542 2142 25594
rect 2142 25542 2172 25594
rect 2196 25542 2206 25594
rect 2206 25542 2252 25594
rect 1956 25540 2012 25542
rect 2036 25540 2092 25542
rect 2116 25540 2172 25542
rect 2196 25540 2252 25542
rect 1956 24506 2012 24508
rect 2036 24506 2092 24508
rect 2116 24506 2172 24508
rect 2196 24506 2252 24508
rect 1956 24454 2002 24506
rect 2002 24454 2012 24506
rect 2036 24454 2066 24506
rect 2066 24454 2078 24506
rect 2078 24454 2092 24506
rect 2116 24454 2130 24506
rect 2130 24454 2142 24506
rect 2142 24454 2172 24506
rect 2196 24454 2206 24506
rect 2206 24454 2252 24506
rect 1956 24452 2012 24454
rect 2036 24452 2092 24454
rect 2116 24452 2172 24454
rect 2196 24452 2252 24454
rect 1956 23418 2012 23420
rect 2036 23418 2092 23420
rect 2116 23418 2172 23420
rect 2196 23418 2252 23420
rect 1956 23366 2002 23418
rect 2002 23366 2012 23418
rect 2036 23366 2066 23418
rect 2066 23366 2078 23418
rect 2078 23366 2092 23418
rect 2116 23366 2130 23418
rect 2130 23366 2142 23418
rect 2142 23366 2172 23418
rect 2196 23366 2206 23418
rect 2206 23366 2252 23418
rect 1956 23364 2012 23366
rect 2036 23364 2092 23366
rect 2116 23364 2172 23366
rect 2196 23364 2252 23366
rect 1956 22330 2012 22332
rect 2036 22330 2092 22332
rect 2116 22330 2172 22332
rect 2196 22330 2252 22332
rect 1956 22278 2002 22330
rect 2002 22278 2012 22330
rect 2036 22278 2066 22330
rect 2066 22278 2078 22330
rect 2078 22278 2092 22330
rect 2116 22278 2130 22330
rect 2130 22278 2142 22330
rect 2142 22278 2172 22330
rect 2196 22278 2206 22330
rect 2206 22278 2252 22330
rect 1956 22276 2012 22278
rect 2036 22276 2092 22278
rect 2116 22276 2172 22278
rect 2196 22276 2252 22278
rect 1956 21242 2012 21244
rect 2036 21242 2092 21244
rect 2116 21242 2172 21244
rect 2196 21242 2252 21244
rect 1956 21190 2002 21242
rect 2002 21190 2012 21242
rect 2036 21190 2066 21242
rect 2066 21190 2078 21242
rect 2078 21190 2092 21242
rect 2116 21190 2130 21242
rect 2130 21190 2142 21242
rect 2142 21190 2172 21242
rect 2196 21190 2206 21242
rect 2206 21190 2252 21242
rect 1956 21188 2012 21190
rect 2036 21188 2092 21190
rect 2116 21188 2172 21190
rect 2196 21188 2252 21190
rect 1956 20154 2012 20156
rect 2036 20154 2092 20156
rect 2116 20154 2172 20156
rect 2196 20154 2252 20156
rect 1956 20102 2002 20154
rect 2002 20102 2012 20154
rect 2036 20102 2066 20154
rect 2066 20102 2078 20154
rect 2078 20102 2092 20154
rect 2116 20102 2130 20154
rect 2130 20102 2142 20154
rect 2142 20102 2172 20154
rect 2196 20102 2206 20154
rect 2206 20102 2252 20154
rect 1956 20100 2012 20102
rect 2036 20100 2092 20102
rect 2116 20100 2172 20102
rect 2196 20100 2252 20102
rect 1956 19066 2012 19068
rect 2036 19066 2092 19068
rect 2116 19066 2172 19068
rect 2196 19066 2252 19068
rect 1956 19014 2002 19066
rect 2002 19014 2012 19066
rect 2036 19014 2066 19066
rect 2066 19014 2078 19066
rect 2078 19014 2092 19066
rect 2116 19014 2130 19066
rect 2130 19014 2142 19066
rect 2142 19014 2172 19066
rect 2196 19014 2206 19066
rect 2206 19014 2252 19066
rect 1956 19012 2012 19014
rect 2036 19012 2092 19014
rect 2116 19012 2172 19014
rect 2196 19012 2252 19014
rect 1956 17978 2012 17980
rect 2036 17978 2092 17980
rect 2116 17978 2172 17980
rect 2196 17978 2252 17980
rect 1956 17926 2002 17978
rect 2002 17926 2012 17978
rect 2036 17926 2066 17978
rect 2066 17926 2078 17978
rect 2078 17926 2092 17978
rect 2116 17926 2130 17978
rect 2130 17926 2142 17978
rect 2142 17926 2172 17978
rect 2196 17926 2206 17978
rect 2206 17926 2252 17978
rect 1956 17924 2012 17926
rect 2036 17924 2092 17926
rect 2116 17924 2172 17926
rect 2196 17924 2252 17926
rect 1956 16890 2012 16892
rect 2036 16890 2092 16892
rect 2116 16890 2172 16892
rect 2196 16890 2252 16892
rect 1956 16838 2002 16890
rect 2002 16838 2012 16890
rect 2036 16838 2066 16890
rect 2066 16838 2078 16890
rect 2078 16838 2092 16890
rect 2116 16838 2130 16890
rect 2130 16838 2142 16890
rect 2142 16838 2172 16890
rect 2196 16838 2206 16890
rect 2206 16838 2252 16890
rect 1956 16836 2012 16838
rect 2036 16836 2092 16838
rect 2116 16836 2172 16838
rect 2196 16836 2252 16838
rect 2616 46810 2672 46812
rect 2696 46810 2752 46812
rect 2776 46810 2832 46812
rect 2856 46810 2912 46812
rect 2616 46758 2662 46810
rect 2662 46758 2672 46810
rect 2696 46758 2726 46810
rect 2726 46758 2738 46810
rect 2738 46758 2752 46810
rect 2776 46758 2790 46810
rect 2790 46758 2802 46810
rect 2802 46758 2832 46810
rect 2856 46758 2866 46810
rect 2866 46758 2912 46810
rect 2616 46756 2672 46758
rect 2696 46756 2752 46758
rect 2776 46756 2832 46758
rect 2856 46756 2912 46758
rect 2616 45722 2672 45724
rect 2696 45722 2752 45724
rect 2776 45722 2832 45724
rect 2856 45722 2912 45724
rect 2616 45670 2662 45722
rect 2662 45670 2672 45722
rect 2696 45670 2726 45722
rect 2726 45670 2738 45722
rect 2738 45670 2752 45722
rect 2776 45670 2790 45722
rect 2790 45670 2802 45722
rect 2802 45670 2832 45722
rect 2856 45670 2866 45722
rect 2866 45670 2912 45722
rect 2616 45668 2672 45670
rect 2696 45668 2752 45670
rect 2776 45668 2832 45670
rect 2856 45668 2912 45670
rect 2616 44634 2672 44636
rect 2696 44634 2752 44636
rect 2776 44634 2832 44636
rect 2856 44634 2912 44636
rect 2616 44582 2662 44634
rect 2662 44582 2672 44634
rect 2696 44582 2726 44634
rect 2726 44582 2738 44634
rect 2738 44582 2752 44634
rect 2776 44582 2790 44634
rect 2790 44582 2802 44634
rect 2802 44582 2832 44634
rect 2856 44582 2866 44634
rect 2866 44582 2912 44634
rect 2616 44580 2672 44582
rect 2696 44580 2752 44582
rect 2776 44580 2832 44582
rect 2856 44580 2912 44582
rect 2616 43546 2672 43548
rect 2696 43546 2752 43548
rect 2776 43546 2832 43548
rect 2856 43546 2912 43548
rect 2616 43494 2662 43546
rect 2662 43494 2672 43546
rect 2696 43494 2726 43546
rect 2726 43494 2738 43546
rect 2738 43494 2752 43546
rect 2776 43494 2790 43546
rect 2790 43494 2802 43546
rect 2802 43494 2832 43546
rect 2856 43494 2866 43546
rect 2866 43494 2912 43546
rect 2616 43492 2672 43494
rect 2696 43492 2752 43494
rect 2776 43492 2832 43494
rect 2856 43492 2912 43494
rect 2616 42458 2672 42460
rect 2696 42458 2752 42460
rect 2776 42458 2832 42460
rect 2856 42458 2912 42460
rect 2616 42406 2662 42458
rect 2662 42406 2672 42458
rect 2696 42406 2726 42458
rect 2726 42406 2738 42458
rect 2738 42406 2752 42458
rect 2776 42406 2790 42458
rect 2790 42406 2802 42458
rect 2802 42406 2832 42458
rect 2856 42406 2866 42458
rect 2866 42406 2912 42458
rect 2616 42404 2672 42406
rect 2696 42404 2752 42406
rect 2776 42404 2832 42406
rect 2856 42404 2912 42406
rect 2616 41370 2672 41372
rect 2696 41370 2752 41372
rect 2776 41370 2832 41372
rect 2856 41370 2912 41372
rect 2616 41318 2662 41370
rect 2662 41318 2672 41370
rect 2696 41318 2726 41370
rect 2726 41318 2738 41370
rect 2738 41318 2752 41370
rect 2776 41318 2790 41370
rect 2790 41318 2802 41370
rect 2802 41318 2832 41370
rect 2856 41318 2866 41370
rect 2866 41318 2912 41370
rect 2616 41316 2672 41318
rect 2696 41316 2752 41318
rect 2776 41316 2832 41318
rect 2856 41316 2912 41318
rect 2616 40282 2672 40284
rect 2696 40282 2752 40284
rect 2776 40282 2832 40284
rect 2856 40282 2912 40284
rect 2616 40230 2662 40282
rect 2662 40230 2672 40282
rect 2696 40230 2726 40282
rect 2726 40230 2738 40282
rect 2738 40230 2752 40282
rect 2776 40230 2790 40282
rect 2790 40230 2802 40282
rect 2802 40230 2832 40282
rect 2856 40230 2866 40282
rect 2866 40230 2912 40282
rect 2616 40228 2672 40230
rect 2696 40228 2752 40230
rect 2776 40228 2832 40230
rect 2856 40228 2912 40230
rect 2616 39194 2672 39196
rect 2696 39194 2752 39196
rect 2776 39194 2832 39196
rect 2856 39194 2912 39196
rect 2616 39142 2662 39194
rect 2662 39142 2672 39194
rect 2696 39142 2726 39194
rect 2726 39142 2738 39194
rect 2738 39142 2752 39194
rect 2776 39142 2790 39194
rect 2790 39142 2802 39194
rect 2802 39142 2832 39194
rect 2856 39142 2866 39194
rect 2866 39142 2912 39194
rect 2616 39140 2672 39142
rect 2696 39140 2752 39142
rect 2776 39140 2832 39142
rect 2856 39140 2912 39142
rect 2616 38106 2672 38108
rect 2696 38106 2752 38108
rect 2776 38106 2832 38108
rect 2856 38106 2912 38108
rect 2616 38054 2662 38106
rect 2662 38054 2672 38106
rect 2696 38054 2726 38106
rect 2726 38054 2738 38106
rect 2738 38054 2752 38106
rect 2776 38054 2790 38106
rect 2790 38054 2802 38106
rect 2802 38054 2832 38106
rect 2856 38054 2866 38106
rect 2866 38054 2912 38106
rect 2616 38052 2672 38054
rect 2696 38052 2752 38054
rect 2776 38052 2832 38054
rect 2856 38052 2912 38054
rect 2616 37018 2672 37020
rect 2696 37018 2752 37020
rect 2776 37018 2832 37020
rect 2856 37018 2912 37020
rect 2616 36966 2662 37018
rect 2662 36966 2672 37018
rect 2696 36966 2726 37018
rect 2726 36966 2738 37018
rect 2738 36966 2752 37018
rect 2776 36966 2790 37018
rect 2790 36966 2802 37018
rect 2802 36966 2832 37018
rect 2856 36966 2866 37018
rect 2866 36966 2912 37018
rect 2616 36964 2672 36966
rect 2696 36964 2752 36966
rect 2776 36964 2832 36966
rect 2856 36964 2912 36966
rect 2616 35930 2672 35932
rect 2696 35930 2752 35932
rect 2776 35930 2832 35932
rect 2856 35930 2912 35932
rect 2616 35878 2662 35930
rect 2662 35878 2672 35930
rect 2696 35878 2726 35930
rect 2726 35878 2738 35930
rect 2738 35878 2752 35930
rect 2776 35878 2790 35930
rect 2790 35878 2802 35930
rect 2802 35878 2832 35930
rect 2856 35878 2866 35930
rect 2866 35878 2912 35930
rect 2616 35876 2672 35878
rect 2696 35876 2752 35878
rect 2776 35876 2832 35878
rect 2856 35876 2912 35878
rect 2616 34842 2672 34844
rect 2696 34842 2752 34844
rect 2776 34842 2832 34844
rect 2856 34842 2912 34844
rect 2616 34790 2662 34842
rect 2662 34790 2672 34842
rect 2696 34790 2726 34842
rect 2726 34790 2738 34842
rect 2738 34790 2752 34842
rect 2776 34790 2790 34842
rect 2790 34790 2802 34842
rect 2802 34790 2832 34842
rect 2856 34790 2866 34842
rect 2866 34790 2912 34842
rect 2616 34788 2672 34790
rect 2696 34788 2752 34790
rect 2776 34788 2832 34790
rect 2856 34788 2912 34790
rect 2616 33754 2672 33756
rect 2696 33754 2752 33756
rect 2776 33754 2832 33756
rect 2856 33754 2912 33756
rect 2616 33702 2662 33754
rect 2662 33702 2672 33754
rect 2696 33702 2726 33754
rect 2726 33702 2738 33754
rect 2738 33702 2752 33754
rect 2776 33702 2790 33754
rect 2790 33702 2802 33754
rect 2802 33702 2832 33754
rect 2856 33702 2866 33754
rect 2866 33702 2912 33754
rect 2616 33700 2672 33702
rect 2696 33700 2752 33702
rect 2776 33700 2832 33702
rect 2856 33700 2912 33702
rect 2616 32666 2672 32668
rect 2696 32666 2752 32668
rect 2776 32666 2832 32668
rect 2856 32666 2912 32668
rect 2616 32614 2662 32666
rect 2662 32614 2672 32666
rect 2696 32614 2726 32666
rect 2726 32614 2738 32666
rect 2738 32614 2752 32666
rect 2776 32614 2790 32666
rect 2790 32614 2802 32666
rect 2802 32614 2832 32666
rect 2856 32614 2866 32666
rect 2866 32614 2912 32666
rect 2616 32612 2672 32614
rect 2696 32612 2752 32614
rect 2776 32612 2832 32614
rect 2856 32612 2912 32614
rect 2616 31578 2672 31580
rect 2696 31578 2752 31580
rect 2776 31578 2832 31580
rect 2856 31578 2912 31580
rect 2616 31526 2662 31578
rect 2662 31526 2672 31578
rect 2696 31526 2726 31578
rect 2726 31526 2738 31578
rect 2738 31526 2752 31578
rect 2776 31526 2790 31578
rect 2790 31526 2802 31578
rect 2802 31526 2832 31578
rect 2856 31526 2866 31578
rect 2866 31526 2912 31578
rect 2616 31524 2672 31526
rect 2696 31524 2752 31526
rect 2776 31524 2832 31526
rect 2856 31524 2912 31526
rect 2616 30490 2672 30492
rect 2696 30490 2752 30492
rect 2776 30490 2832 30492
rect 2856 30490 2912 30492
rect 2616 30438 2662 30490
rect 2662 30438 2672 30490
rect 2696 30438 2726 30490
rect 2726 30438 2738 30490
rect 2738 30438 2752 30490
rect 2776 30438 2790 30490
rect 2790 30438 2802 30490
rect 2802 30438 2832 30490
rect 2856 30438 2866 30490
rect 2866 30438 2912 30490
rect 2616 30436 2672 30438
rect 2696 30436 2752 30438
rect 2776 30436 2832 30438
rect 2856 30436 2912 30438
rect 2616 29402 2672 29404
rect 2696 29402 2752 29404
rect 2776 29402 2832 29404
rect 2856 29402 2912 29404
rect 2616 29350 2662 29402
rect 2662 29350 2672 29402
rect 2696 29350 2726 29402
rect 2726 29350 2738 29402
rect 2738 29350 2752 29402
rect 2776 29350 2790 29402
rect 2790 29350 2802 29402
rect 2802 29350 2832 29402
rect 2856 29350 2866 29402
rect 2866 29350 2912 29402
rect 2616 29348 2672 29350
rect 2696 29348 2752 29350
rect 2776 29348 2832 29350
rect 2856 29348 2912 29350
rect 2616 28314 2672 28316
rect 2696 28314 2752 28316
rect 2776 28314 2832 28316
rect 2856 28314 2912 28316
rect 2616 28262 2662 28314
rect 2662 28262 2672 28314
rect 2696 28262 2726 28314
rect 2726 28262 2738 28314
rect 2738 28262 2752 28314
rect 2776 28262 2790 28314
rect 2790 28262 2802 28314
rect 2802 28262 2832 28314
rect 2856 28262 2866 28314
rect 2866 28262 2912 28314
rect 2616 28260 2672 28262
rect 2696 28260 2752 28262
rect 2776 28260 2832 28262
rect 2856 28260 2912 28262
rect 2616 27226 2672 27228
rect 2696 27226 2752 27228
rect 2776 27226 2832 27228
rect 2856 27226 2912 27228
rect 2616 27174 2662 27226
rect 2662 27174 2672 27226
rect 2696 27174 2726 27226
rect 2726 27174 2738 27226
rect 2738 27174 2752 27226
rect 2776 27174 2790 27226
rect 2790 27174 2802 27226
rect 2802 27174 2832 27226
rect 2856 27174 2866 27226
rect 2866 27174 2912 27226
rect 2616 27172 2672 27174
rect 2696 27172 2752 27174
rect 2776 27172 2832 27174
rect 2856 27172 2912 27174
rect 2616 26138 2672 26140
rect 2696 26138 2752 26140
rect 2776 26138 2832 26140
rect 2856 26138 2912 26140
rect 2616 26086 2662 26138
rect 2662 26086 2672 26138
rect 2696 26086 2726 26138
rect 2726 26086 2738 26138
rect 2738 26086 2752 26138
rect 2776 26086 2790 26138
rect 2790 26086 2802 26138
rect 2802 26086 2832 26138
rect 2856 26086 2866 26138
rect 2866 26086 2912 26138
rect 2616 26084 2672 26086
rect 2696 26084 2752 26086
rect 2776 26084 2832 26086
rect 2856 26084 2912 26086
rect 1956 15802 2012 15804
rect 2036 15802 2092 15804
rect 2116 15802 2172 15804
rect 2196 15802 2252 15804
rect 1956 15750 2002 15802
rect 2002 15750 2012 15802
rect 2036 15750 2066 15802
rect 2066 15750 2078 15802
rect 2078 15750 2092 15802
rect 2116 15750 2130 15802
rect 2130 15750 2142 15802
rect 2142 15750 2172 15802
rect 2196 15750 2206 15802
rect 2206 15750 2252 15802
rect 1956 15748 2012 15750
rect 2036 15748 2092 15750
rect 2116 15748 2172 15750
rect 2196 15748 2252 15750
rect 1956 14714 2012 14716
rect 2036 14714 2092 14716
rect 2116 14714 2172 14716
rect 2196 14714 2252 14716
rect 1956 14662 2002 14714
rect 2002 14662 2012 14714
rect 2036 14662 2066 14714
rect 2066 14662 2078 14714
rect 2078 14662 2092 14714
rect 2116 14662 2130 14714
rect 2130 14662 2142 14714
rect 2142 14662 2172 14714
rect 2196 14662 2206 14714
rect 2206 14662 2252 14714
rect 1956 14660 2012 14662
rect 2036 14660 2092 14662
rect 2116 14660 2172 14662
rect 2196 14660 2252 14662
rect 1956 13626 2012 13628
rect 2036 13626 2092 13628
rect 2116 13626 2172 13628
rect 2196 13626 2252 13628
rect 1956 13574 2002 13626
rect 2002 13574 2012 13626
rect 2036 13574 2066 13626
rect 2066 13574 2078 13626
rect 2078 13574 2092 13626
rect 2116 13574 2130 13626
rect 2130 13574 2142 13626
rect 2142 13574 2172 13626
rect 2196 13574 2206 13626
rect 2206 13574 2252 13626
rect 1956 13572 2012 13574
rect 2036 13572 2092 13574
rect 2116 13572 2172 13574
rect 2196 13572 2252 13574
rect 1956 12538 2012 12540
rect 2036 12538 2092 12540
rect 2116 12538 2172 12540
rect 2196 12538 2252 12540
rect 1956 12486 2002 12538
rect 2002 12486 2012 12538
rect 2036 12486 2066 12538
rect 2066 12486 2078 12538
rect 2078 12486 2092 12538
rect 2116 12486 2130 12538
rect 2130 12486 2142 12538
rect 2142 12486 2172 12538
rect 2196 12486 2206 12538
rect 2206 12486 2252 12538
rect 1956 12484 2012 12486
rect 2036 12484 2092 12486
rect 2116 12484 2172 12486
rect 2196 12484 2252 12486
rect 1956 11450 2012 11452
rect 2036 11450 2092 11452
rect 2116 11450 2172 11452
rect 2196 11450 2252 11452
rect 1956 11398 2002 11450
rect 2002 11398 2012 11450
rect 2036 11398 2066 11450
rect 2066 11398 2078 11450
rect 2078 11398 2092 11450
rect 2116 11398 2130 11450
rect 2130 11398 2142 11450
rect 2142 11398 2172 11450
rect 2196 11398 2206 11450
rect 2206 11398 2252 11450
rect 1956 11396 2012 11398
rect 2036 11396 2092 11398
rect 2116 11396 2172 11398
rect 2196 11396 2252 11398
rect 1858 11056 1914 11112
rect 1956 10362 2012 10364
rect 2036 10362 2092 10364
rect 2116 10362 2172 10364
rect 2196 10362 2252 10364
rect 1956 10310 2002 10362
rect 2002 10310 2012 10362
rect 2036 10310 2066 10362
rect 2066 10310 2078 10362
rect 2078 10310 2092 10362
rect 2116 10310 2130 10362
rect 2130 10310 2142 10362
rect 2142 10310 2172 10362
rect 2196 10310 2206 10362
rect 2206 10310 2252 10362
rect 1956 10308 2012 10310
rect 2036 10308 2092 10310
rect 2116 10308 2172 10310
rect 2196 10308 2252 10310
rect 1956 9274 2012 9276
rect 2036 9274 2092 9276
rect 2116 9274 2172 9276
rect 2196 9274 2252 9276
rect 1956 9222 2002 9274
rect 2002 9222 2012 9274
rect 2036 9222 2066 9274
rect 2066 9222 2078 9274
rect 2078 9222 2092 9274
rect 2116 9222 2130 9274
rect 2130 9222 2142 9274
rect 2142 9222 2172 9274
rect 2196 9222 2206 9274
rect 2206 9222 2252 9274
rect 1956 9220 2012 9222
rect 2036 9220 2092 9222
rect 2116 9220 2172 9222
rect 2196 9220 2252 9222
rect 1956 8186 2012 8188
rect 2036 8186 2092 8188
rect 2116 8186 2172 8188
rect 2196 8186 2252 8188
rect 1956 8134 2002 8186
rect 2002 8134 2012 8186
rect 2036 8134 2066 8186
rect 2066 8134 2078 8186
rect 2078 8134 2092 8186
rect 2116 8134 2130 8186
rect 2130 8134 2142 8186
rect 2142 8134 2172 8186
rect 2196 8134 2206 8186
rect 2206 8134 2252 8186
rect 1956 8132 2012 8134
rect 2036 8132 2092 8134
rect 2116 8132 2172 8134
rect 2196 8132 2252 8134
rect 1956 7098 2012 7100
rect 2036 7098 2092 7100
rect 2116 7098 2172 7100
rect 2196 7098 2252 7100
rect 1956 7046 2002 7098
rect 2002 7046 2012 7098
rect 2036 7046 2066 7098
rect 2066 7046 2078 7098
rect 2078 7046 2092 7098
rect 2116 7046 2130 7098
rect 2130 7046 2142 7098
rect 2142 7046 2172 7098
rect 2196 7046 2206 7098
rect 2206 7046 2252 7098
rect 1956 7044 2012 7046
rect 2036 7044 2092 7046
rect 2116 7044 2172 7046
rect 2196 7044 2252 7046
rect 1956 6010 2012 6012
rect 2036 6010 2092 6012
rect 2116 6010 2172 6012
rect 2196 6010 2252 6012
rect 1956 5958 2002 6010
rect 2002 5958 2012 6010
rect 2036 5958 2066 6010
rect 2066 5958 2078 6010
rect 2078 5958 2092 6010
rect 2116 5958 2130 6010
rect 2130 5958 2142 6010
rect 2142 5958 2172 6010
rect 2196 5958 2206 6010
rect 2206 5958 2252 6010
rect 1956 5956 2012 5958
rect 2036 5956 2092 5958
rect 2116 5956 2172 5958
rect 2196 5956 2252 5958
rect 1956 4922 2012 4924
rect 2036 4922 2092 4924
rect 2116 4922 2172 4924
rect 2196 4922 2252 4924
rect 1956 4870 2002 4922
rect 2002 4870 2012 4922
rect 2036 4870 2066 4922
rect 2066 4870 2078 4922
rect 2078 4870 2092 4922
rect 2116 4870 2130 4922
rect 2130 4870 2142 4922
rect 2142 4870 2172 4922
rect 2196 4870 2206 4922
rect 2206 4870 2252 4922
rect 1956 4868 2012 4870
rect 2036 4868 2092 4870
rect 2116 4868 2172 4870
rect 2196 4868 2252 4870
rect 846 4564 848 4584
rect 848 4564 900 4584
rect 900 4564 902 4584
rect 846 4528 902 4564
rect 1956 3834 2012 3836
rect 2036 3834 2092 3836
rect 2116 3834 2172 3836
rect 2196 3834 2252 3836
rect 1956 3782 2002 3834
rect 2002 3782 2012 3834
rect 2036 3782 2066 3834
rect 2066 3782 2078 3834
rect 2078 3782 2092 3834
rect 2116 3782 2130 3834
rect 2130 3782 2142 3834
rect 2142 3782 2172 3834
rect 2196 3782 2206 3834
rect 2206 3782 2252 3834
rect 1956 3780 2012 3782
rect 2036 3780 2092 3782
rect 2116 3780 2172 3782
rect 2196 3780 2252 3782
rect 1956 2746 2012 2748
rect 2036 2746 2092 2748
rect 2116 2746 2172 2748
rect 2196 2746 2252 2748
rect 1956 2694 2002 2746
rect 2002 2694 2012 2746
rect 2036 2694 2066 2746
rect 2066 2694 2078 2746
rect 2078 2694 2092 2746
rect 2116 2694 2130 2746
rect 2130 2694 2142 2746
rect 2142 2694 2172 2746
rect 2196 2694 2206 2746
rect 2206 2694 2252 2746
rect 1956 2692 2012 2694
rect 2036 2692 2092 2694
rect 2116 2692 2172 2694
rect 2196 2692 2252 2694
rect 2616 25050 2672 25052
rect 2696 25050 2752 25052
rect 2776 25050 2832 25052
rect 2856 25050 2912 25052
rect 2616 24998 2662 25050
rect 2662 24998 2672 25050
rect 2696 24998 2726 25050
rect 2726 24998 2738 25050
rect 2738 24998 2752 25050
rect 2776 24998 2790 25050
rect 2790 24998 2802 25050
rect 2802 24998 2832 25050
rect 2856 24998 2866 25050
rect 2866 24998 2912 25050
rect 2616 24996 2672 24998
rect 2696 24996 2752 24998
rect 2776 24996 2832 24998
rect 2856 24996 2912 24998
rect 2616 23962 2672 23964
rect 2696 23962 2752 23964
rect 2776 23962 2832 23964
rect 2856 23962 2912 23964
rect 2616 23910 2662 23962
rect 2662 23910 2672 23962
rect 2696 23910 2726 23962
rect 2726 23910 2738 23962
rect 2738 23910 2752 23962
rect 2776 23910 2790 23962
rect 2790 23910 2802 23962
rect 2802 23910 2832 23962
rect 2856 23910 2866 23962
rect 2866 23910 2912 23962
rect 2616 23908 2672 23910
rect 2696 23908 2752 23910
rect 2776 23908 2832 23910
rect 2856 23908 2912 23910
rect 2616 22874 2672 22876
rect 2696 22874 2752 22876
rect 2776 22874 2832 22876
rect 2856 22874 2912 22876
rect 2616 22822 2662 22874
rect 2662 22822 2672 22874
rect 2696 22822 2726 22874
rect 2726 22822 2738 22874
rect 2738 22822 2752 22874
rect 2776 22822 2790 22874
rect 2790 22822 2802 22874
rect 2802 22822 2832 22874
rect 2856 22822 2866 22874
rect 2866 22822 2912 22874
rect 2616 22820 2672 22822
rect 2696 22820 2752 22822
rect 2776 22820 2832 22822
rect 2856 22820 2912 22822
rect 2616 21786 2672 21788
rect 2696 21786 2752 21788
rect 2776 21786 2832 21788
rect 2856 21786 2912 21788
rect 2616 21734 2662 21786
rect 2662 21734 2672 21786
rect 2696 21734 2726 21786
rect 2726 21734 2738 21786
rect 2738 21734 2752 21786
rect 2776 21734 2790 21786
rect 2790 21734 2802 21786
rect 2802 21734 2832 21786
rect 2856 21734 2866 21786
rect 2866 21734 2912 21786
rect 2616 21732 2672 21734
rect 2696 21732 2752 21734
rect 2776 21732 2832 21734
rect 2856 21732 2912 21734
rect 2616 20698 2672 20700
rect 2696 20698 2752 20700
rect 2776 20698 2832 20700
rect 2856 20698 2912 20700
rect 2616 20646 2662 20698
rect 2662 20646 2672 20698
rect 2696 20646 2726 20698
rect 2726 20646 2738 20698
rect 2738 20646 2752 20698
rect 2776 20646 2790 20698
rect 2790 20646 2802 20698
rect 2802 20646 2832 20698
rect 2856 20646 2866 20698
rect 2866 20646 2912 20698
rect 2616 20644 2672 20646
rect 2696 20644 2752 20646
rect 2776 20644 2832 20646
rect 2856 20644 2912 20646
rect 2616 19610 2672 19612
rect 2696 19610 2752 19612
rect 2776 19610 2832 19612
rect 2856 19610 2912 19612
rect 2616 19558 2662 19610
rect 2662 19558 2672 19610
rect 2696 19558 2726 19610
rect 2726 19558 2738 19610
rect 2738 19558 2752 19610
rect 2776 19558 2790 19610
rect 2790 19558 2802 19610
rect 2802 19558 2832 19610
rect 2856 19558 2866 19610
rect 2866 19558 2912 19610
rect 2616 19556 2672 19558
rect 2696 19556 2752 19558
rect 2776 19556 2832 19558
rect 2856 19556 2912 19558
rect 2616 18522 2672 18524
rect 2696 18522 2752 18524
rect 2776 18522 2832 18524
rect 2856 18522 2912 18524
rect 2616 18470 2662 18522
rect 2662 18470 2672 18522
rect 2696 18470 2726 18522
rect 2726 18470 2738 18522
rect 2738 18470 2752 18522
rect 2776 18470 2790 18522
rect 2790 18470 2802 18522
rect 2802 18470 2832 18522
rect 2856 18470 2866 18522
rect 2866 18470 2912 18522
rect 2616 18468 2672 18470
rect 2696 18468 2752 18470
rect 2776 18468 2832 18470
rect 2856 18468 2912 18470
rect 2616 17434 2672 17436
rect 2696 17434 2752 17436
rect 2776 17434 2832 17436
rect 2856 17434 2912 17436
rect 2616 17382 2662 17434
rect 2662 17382 2672 17434
rect 2696 17382 2726 17434
rect 2726 17382 2738 17434
rect 2738 17382 2752 17434
rect 2776 17382 2790 17434
rect 2790 17382 2802 17434
rect 2802 17382 2832 17434
rect 2856 17382 2866 17434
rect 2866 17382 2912 17434
rect 2616 17380 2672 17382
rect 2696 17380 2752 17382
rect 2776 17380 2832 17382
rect 2856 17380 2912 17382
rect 2616 16346 2672 16348
rect 2696 16346 2752 16348
rect 2776 16346 2832 16348
rect 2856 16346 2912 16348
rect 2616 16294 2662 16346
rect 2662 16294 2672 16346
rect 2696 16294 2726 16346
rect 2726 16294 2738 16346
rect 2738 16294 2752 16346
rect 2776 16294 2790 16346
rect 2790 16294 2802 16346
rect 2802 16294 2832 16346
rect 2856 16294 2866 16346
rect 2866 16294 2912 16346
rect 2616 16292 2672 16294
rect 2696 16292 2752 16294
rect 2776 16292 2832 16294
rect 2856 16292 2912 16294
rect 2616 15258 2672 15260
rect 2696 15258 2752 15260
rect 2776 15258 2832 15260
rect 2856 15258 2912 15260
rect 2616 15206 2662 15258
rect 2662 15206 2672 15258
rect 2696 15206 2726 15258
rect 2726 15206 2738 15258
rect 2738 15206 2752 15258
rect 2776 15206 2790 15258
rect 2790 15206 2802 15258
rect 2802 15206 2832 15258
rect 2856 15206 2866 15258
rect 2866 15206 2912 15258
rect 2616 15204 2672 15206
rect 2696 15204 2752 15206
rect 2776 15204 2832 15206
rect 2856 15204 2912 15206
rect 2616 14170 2672 14172
rect 2696 14170 2752 14172
rect 2776 14170 2832 14172
rect 2856 14170 2912 14172
rect 2616 14118 2662 14170
rect 2662 14118 2672 14170
rect 2696 14118 2726 14170
rect 2726 14118 2738 14170
rect 2738 14118 2752 14170
rect 2776 14118 2790 14170
rect 2790 14118 2802 14170
rect 2802 14118 2832 14170
rect 2856 14118 2866 14170
rect 2866 14118 2912 14170
rect 2616 14116 2672 14118
rect 2696 14116 2752 14118
rect 2776 14116 2832 14118
rect 2856 14116 2912 14118
rect 2616 13082 2672 13084
rect 2696 13082 2752 13084
rect 2776 13082 2832 13084
rect 2856 13082 2912 13084
rect 2616 13030 2662 13082
rect 2662 13030 2672 13082
rect 2696 13030 2726 13082
rect 2726 13030 2738 13082
rect 2738 13030 2752 13082
rect 2776 13030 2790 13082
rect 2790 13030 2802 13082
rect 2802 13030 2832 13082
rect 2856 13030 2866 13082
rect 2866 13030 2912 13082
rect 2616 13028 2672 13030
rect 2696 13028 2752 13030
rect 2776 13028 2832 13030
rect 2856 13028 2912 13030
rect 2616 11994 2672 11996
rect 2696 11994 2752 11996
rect 2776 11994 2832 11996
rect 2856 11994 2912 11996
rect 2616 11942 2662 11994
rect 2662 11942 2672 11994
rect 2696 11942 2726 11994
rect 2726 11942 2738 11994
rect 2738 11942 2752 11994
rect 2776 11942 2790 11994
rect 2790 11942 2802 11994
rect 2802 11942 2832 11994
rect 2856 11942 2866 11994
rect 2866 11942 2912 11994
rect 2616 11940 2672 11942
rect 2696 11940 2752 11942
rect 2776 11940 2832 11942
rect 2856 11940 2912 11942
rect 2616 10906 2672 10908
rect 2696 10906 2752 10908
rect 2776 10906 2832 10908
rect 2856 10906 2912 10908
rect 2616 10854 2662 10906
rect 2662 10854 2672 10906
rect 2696 10854 2726 10906
rect 2726 10854 2738 10906
rect 2738 10854 2752 10906
rect 2776 10854 2790 10906
rect 2790 10854 2802 10906
rect 2802 10854 2832 10906
rect 2856 10854 2866 10906
rect 2866 10854 2912 10906
rect 2616 10852 2672 10854
rect 2696 10852 2752 10854
rect 2776 10852 2832 10854
rect 2856 10852 2912 10854
rect 2616 9818 2672 9820
rect 2696 9818 2752 9820
rect 2776 9818 2832 9820
rect 2856 9818 2912 9820
rect 2616 9766 2662 9818
rect 2662 9766 2672 9818
rect 2696 9766 2726 9818
rect 2726 9766 2738 9818
rect 2738 9766 2752 9818
rect 2776 9766 2790 9818
rect 2790 9766 2802 9818
rect 2802 9766 2832 9818
rect 2856 9766 2866 9818
rect 2866 9766 2912 9818
rect 2616 9764 2672 9766
rect 2696 9764 2752 9766
rect 2776 9764 2832 9766
rect 2856 9764 2912 9766
rect 2616 8730 2672 8732
rect 2696 8730 2752 8732
rect 2776 8730 2832 8732
rect 2856 8730 2912 8732
rect 2616 8678 2662 8730
rect 2662 8678 2672 8730
rect 2696 8678 2726 8730
rect 2726 8678 2738 8730
rect 2738 8678 2752 8730
rect 2776 8678 2790 8730
rect 2790 8678 2802 8730
rect 2802 8678 2832 8730
rect 2856 8678 2866 8730
rect 2866 8678 2912 8730
rect 2616 8676 2672 8678
rect 2696 8676 2752 8678
rect 2776 8676 2832 8678
rect 2856 8676 2912 8678
rect 2616 7642 2672 7644
rect 2696 7642 2752 7644
rect 2776 7642 2832 7644
rect 2856 7642 2912 7644
rect 2616 7590 2662 7642
rect 2662 7590 2672 7642
rect 2696 7590 2726 7642
rect 2726 7590 2738 7642
rect 2738 7590 2752 7642
rect 2776 7590 2790 7642
rect 2790 7590 2802 7642
rect 2802 7590 2832 7642
rect 2856 7590 2866 7642
rect 2866 7590 2912 7642
rect 2616 7588 2672 7590
rect 2696 7588 2752 7590
rect 2776 7588 2832 7590
rect 2856 7588 2912 7590
rect 2616 6554 2672 6556
rect 2696 6554 2752 6556
rect 2776 6554 2832 6556
rect 2856 6554 2912 6556
rect 2616 6502 2662 6554
rect 2662 6502 2672 6554
rect 2696 6502 2726 6554
rect 2726 6502 2738 6554
rect 2738 6502 2752 6554
rect 2776 6502 2790 6554
rect 2790 6502 2802 6554
rect 2802 6502 2832 6554
rect 2856 6502 2866 6554
rect 2866 6502 2912 6554
rect 2616 6500 2672 6502
rect 2696 6500 2752 6502
rect 2776 6500 2832 6502
rect 2856 6500 2912 6502
rect 2616 5466 2672 5468
rect 2696 5466 2752 5468
rect 2776 5466 2832 5468
rect 2856 5466 2912 5468
rect 2616 5414 2662 5466
rect 2662 5414 2672 5466
rect 2696 5414 2726 5466
rect 2726 5414 2738 5466
rect 2738 5414 2752 5466
rect 2776 5414 2790 5466
rect 2790 5414 2802 5466
rect 2802 5414 2832 5466
rect 2856 5414 2866 5466
rect 2866 5414 2912 5466
rect 2616 5412 2672 5414
rect 2696 5412 2752 5414
rect 2776 5412 2832 5414
rect 2856 5412 2912 5414
rect 4158 36624 4214 36680
rect 3790 11600 3846 11656
rect 2616 4378 2672 4380
rect 2696 4378 2752 4380
rect 2776 4378 2832 4380
rect 2856 4378 2912 4380
rect 2616 4326 2662 4378
rect 2662 4326 2672 4378
rect 2696 4326 2726 4378
rect 2726 4326 2738 4378
rect 2738 4326 2752 4378
rect 2776 4326 2790 4378
rect 2790 4326 2802 4378
rect 2802 4326 2832 4378
rect 2856 4326 2866 4378
rect 2866 4326 2912 4378
rect 2616 4324 2672 4326
rect 2696 4324 2752 4326
rect 2776 4324 2832 4326
rect 2856 4324 2912 4326
rect 7616 67482 7672 67484
rect 7696 67482 7752 67484
rect 7776 67482 7832 67484
rect 7856 67482 7912 67484
rect 7616 67430 7662 67482
rect 7662 67430 7672 67482
rect 7696 67430 7726 67482
rect 7726 67430 7738 67482
rect 7738 67430 7752 67482
rect 7776 67430 7790 67482
rect 7790 67430 7802 67482
rect 7802 67430 7832 67482
rect 7856 67430 7866 67482
rect 7866 67430 7912 67482
rect 7616 67428 7672 67430
rect 7696 67428 7752 67430
rect 7776 67428 7832 67430
rect 7856 67428 7912 67430
rect 6956 66938 7012 66940
rect 7036 66938 7092 66940
rect 7116 66938 7172 66940
rect 7196 66938 7252 66940
rect 6956 66886 7002 66938
rect 7002 66886 7012 66938
rect 7036 66886 7066 66938
rect 7066 66886 7078 66938
rect 7078 66886 7092 66938
rect 7116 66886 7130 66938
rect 7130 66886 7142 66938
rect 7142 66886 7172 66938
rect 7196 66886 7206 66938
rect 7206 66886 7252 66938
rect 6956 66884 7012 66886
rect 7036 66884 7092 66886
rect 7116 66884 7172 66886
rect 7196 66884 7252 66886
rect 6956 65850 7012 65852
rect 7036 65850 7092 65852
rect 7116 65850 7172 65852
rect 7196 65850 7252 65852
rect 6956 65798 7002 65850
rect 7002 65798 7012 65850
rect 7036 65798 7066 65850
rect 7066 65798 7078 65850
rect 7078 65798 7092 65850
rect 7116 65798 7130 65850
rect 7130 65798 7142 65850
rect 7142 65798 7172 65850
rect 7196 65798 7206 65850
rect 7206 65798 7252 65850
rect 6956 65796 7012 65798
rect 7036 65796 7092 65798
rect 7116 65796 7172 65798
rect 7196 65796 7252 65798
rect 6956 64762 7012 64764
rect 7036 64762 7092 64764
rect 7116 64762 7172 64764
rect 7196 64762 7252 64764
rect 6956 64710 7002 64762
rect 7002 64710 7012 64762
rect 7036 64710 7066 64762
rect 7066 64710 7078 64762
rect 7078 64710 7092 64762
rect 7116 64710 7130 64762
rect 7130 64710 7142 64762
rect 7142 64710 7172 64762
rect 7196 64710 7206 64762
rect 7206 64710 7252 64762
rect 6956 64708 7012 64710
rect 7036 64708 7092 64710
rect 7116 64708 7172 64710
rect 7196 64708 7252 64710
rect 6956 63674 7012 63676
rect 7036 63674 7092 63676
rect 7116 63674 7172 63676
rect 7196 63674 7252 63676
rect 6956 63622 7002 63674
rect 7002 63622 7012 63674
rect 7036 63622 7066 63674
rect 7066 63622 7078 63674
rect 7078 63622 7092 63674
rect 7116 63622 7130 63674
rect 7130 63622 7142 63674
rect 7142 63622 7172 63674
rect 7196 63622 7206 63674
rect 7206 63622 7252 63674
rect 6956 63620 7012 63622
rect 7036 63620 7092 63622
rect 7116 63620 7172 63622
rect 7196 63620 7252 63622
rect 6956 62586 7012 62588
rect 7036 62586 7092 62588
rect 7116 62586 7172 62588
rect 7196 62586 7252 62588
rect 6956 62534 7002 62586
rect 7002 62534 7012 62586
rect 7036 62534 7066 62586
rect 7066 62534 7078 62586
rect 7078 62534 7092 62586
rect 7116 62534 7130 62586
rect 7130 62534 7142 62586
rect 7142 62534 7172 62586
rect 7196 62534 7206 62586
rect 7206 62534 7252 62586
rect 6956 62532 7012 62534
rect 7036 62532 7092 62534
rect 7116 62532 7172 62534
rect 7196 62532 7252 62534
rect 6956 61498 7012 61500
rect 7036 61498 7092 61500
rect 7116 61498 7172 61500
rect 7196 61498 7252 61500
rect 6956 61446 7002 61498
rect 7002 61446 7012 61498
rect 7036 61446 7066 61498
rect 7066 61446 7078 61498
rect 7078 61446 7092 61498
rect 7116 61446 7130 61498
rect 7130 61446 7142 61498
rect 7142 61446 7172 61498
rect 7196 61446 7206 61498
rect 7206 61446 7252 61498
rect 6956 61444 7012 61446
rect 7036 61444 7092 61446
rect 7116 61444 7172 61446
rect 7196 61444 7252 61446
rect 6956 60410 7012 60412
rect 7036 60410 7092 60412
rect 7116 60410 7172 60412
rect 7196 60410 7252 60412
rect 6956 60358 7002 60410
rect 7002 60358 7012 60410
rect 7036 60358 7066 60410
rect 7066 60358 7078 60410
rect 7078 60358 7092 60410
rect 7116 60358 7130 60410
rect 7130 60358 7142 60410
rect 7142 60358 7172 60410
rect 7196 60358 7206 60410
rect 7206 60358 7252 60410
rect 6956 60356 7012 60358
rect 7036 60356 7092 60358
rect 7116 60356 7172 60358
rect 7196 60356 7252 60358
rect 6956 59322 7012 59324
rect 7036 59322 7092 59324
rect 7116 59322 7172 59324
rect 7196 59322 7252 59324
rect 6956 59270 7002 59322
rect 7002 59270 7012 59322
rect 7036 59270 7066 59322
rect 7066 59270 7078 59322
rect 7078 59270 7092 59322
rect 7116 59270 7130 59322
rect 7130 59270 7142 59322
rect 7142 59270 7172 59322
rect 7196 59270 7206 59322
rect 7206 59270 7252 59322
rect 6956 59268 7012 59270
rect 7036 59268 7092 59270
rect 7116 59268 7172 59270
rect 7196 59268 7252 59270
rect 6956 58234 7012 58236
rect 7036 58234 7092 58236
rect 7116 58234 7172 58236
rect 7196 58234 7252 58236
rect 6956 58182 7002 58234
rect 7002 58182 7012 58234
rect 7036 58182 7066 58234
rect 7066 58182 7078 58234
rect 7078 58182 7092 58234
rect 7116 58182 7130 58234
rect 7130 58182 7142 58234
rect 7142 58182 7172 58234
rect 7196 58182 7206 58234
rect 7206 58182 7252 58234
rect 6956 58180 7012 58182
rect 7036 58180 7092 58182
rect 7116 58180 7172 58182
rect 7196 58180 7252 58182
rect 6956 57146 7012 57148
rect 7036 57146 7092 57148
rect 7116 57146 7172 57148
rect 7196 57146 7252 57148
rect 6956 57094 7002 57146
rect 7002 57094 7012 57146
rect 7036 57094 7066 57146
rect 7066 57094 7078 57146
rect 7078 57094 7092 57146
rect 7116 57094 7130 57146
rect 7130 57094 7142 57146
rect 7142 57094 7172 57146
rect 7196 57094 7206 57146
rect 7206 57094 7252 57146
rect 6956 57092 7012 57094
rect 7036 57092 7092 57094
rect 7116 57092 7172 57094
rect 7196 57092 7252 57094
rect 6956 56058 7012 56060
rect 7036 56058 7092 56060
rect 7116 56058 7172 56060
rect 7196 56058 7252 56060
rect 6956 56006 7002 56058
rect 7002 56006 7012 56058
rect 7036 56006 7066 56058
rect 7066 56006 7078 56058
rect 7078 56006 7092 56058
rect 7116 56006 7130 56058
rect 7130 56006 7142 56058
rect 7142 56006 7172 56058
rect 7196 56006 7206 56058
rect 7206 56006 7252 56058
rect 6956 56004 7012 56006
rect 7036 56004 7092 56006
rect 7116 56004 7172 56006
rect 7196 56004 7252 56006
rect 6956 54970 7012 54972
rect 7036 54970 7092 54972
rect 7116 54970 7172 54972
rect 7196 54970 7252 54972
rect 6956 54918 7002 54970
rect 7002 54918 7012 54970
rect 7036 54918 7066 54970
rect 7066 54918 7078 54970
rect 7078 54918 7092 54970
rect 7116 54918 7130 54970
rect 7130 54918 7142 54970
rect 7142 54918 7172 54970
rect 7196 54918 7206 54970
rect 7206 54918 7252 54970
rect 6956 54916 7012 54918
rect 7036 54916 7092 54918
rect 7116 54916 7172 54918
rect 7196 54916 7252 54918
rect 6956 53882 7012 53884
rect 7036 53882 7092 53884
rect 7116 53882 7172 53884
rect 7196 53882 7252 53884
rect 6956 53830 7002 53882
rect 7002 53830 7012 53882
rect 7036 53830 7066 53882
rect 7066 53830 7078 53882
rect 7078 53830 7092 53882
rect 7116 53830 7130 53882
rect 7130 53830 7142 53882
rect 7142 53830 7172 53882
rect 7196 53830 7206 53882
rect 7206 53830 7252 53882
rect 6956 53828 7012 53830
rect 7036 53828 7092 53830
rect 7116 53828 7172 53830
rect 7196 53828 7252 53830
rect 6956 52794 7012 52796
rect 7036 52794 7092 52796
rect 7116 52794 7172 52796
rect 7196 52794 7252 52796
rect 6956 52742 7002 52794
rect 7002 52742 7012 52794
rect 7036 52742 7066 52794
rect 7066 52742 7078 52794
rect 7078 52742 7092 52794
rect 7116 52742 7130 52794
rect 7130 52742 7142 52794
rect 7142 52742 7172 52794
rect 7196 52742 7206 52794
rect 7206 52742 7252 52794
rect 6956 52740 7012 52742
rect 7036 52740 7092 52742
rect 7116 52740 7172 52742
rect 7196 52740 7252 52742
rect 6956 51706 7012 51708
rect 7036 51706 7092 51708
rect 7116 51706 7172 51708
rect 7196 51706 7252 51708
rect 6956 51654 7002 51706
rect 7002 51654 7012 51706
rect 7036 51654 7066 51706
rect 7066 51654 7078 51706
rect 7078 51654 7092 51706
rect 7116 51654 7130 51706
rect 7130 51654 7142 51706
rect 7142 51654 7172 51706
rect 7196 51654 7206 51706
rect 7206 51654 7252 51706
rect 6956 51652 7012 51654
rect 7036 51652 7092 51654
rect 7116 51652 7172 51654
rect 7196 51652 7252 51654
rect 6734 35128 6790 35184
rect 6956 50618 7012 50620
rect 7036 50618 7092 50620
rect 7116 50618 7172 50620
rect 7196 50618 7252 50620
rect 6956 50566 7002 50618
rect 7002 50566 7012 50618
rect 7036 50566 7066 50618
rect 7066 50566 7078 50618
rect 7078 50566 7092 50618
rect 7116 50566 7130 50618
rect 7130 50566 7142 50618
rect 7142 50566 7172 50618
rect 7196 50566 7206 50618
rect 7206 50566 7252 50618
rect 6956 50564 7012 50566
rect 7036 50564 7092 50566
rect 7116 50564 7172 50566
rect 7196 50564 7252 50566
rect 6956 49530 7012 49532
rect 7036 49530 7092 49532
rect 7116 49530 7172 49532
rect 7196 49530 7252 49532
rect 6956 49478 7002 49530
rect 7002 49478 7012 49530
rect 7036 49478 7066 49530
rect 7066 49478 7078 49530
rect 7078 49478 7092 49530
rect 7116 49478 7130 49530
rect 7130 49478 7142 49530
rect 7142 49478 7172 49530
rect 7196 49478 7206 49530
rect 7206 49478 7252 49530
rect 6956 49476 7012 49478
rect 7036 49476 7092 49478
rect 7116 49476 7172 49478
rect 7196 49476 7252 49478
rect 6956 48442 7012 48444
rect 7036 48442 7092 48444
rect 7116 48442 7172 48444
rect 7196 48442 7252 48444
rect 6956 48390 7002 48442
rect 7002 48390 7012 48442
rect 7036 48390 7066 48442
rect 7066 48390 7078 48442
rect 7078 48390 7092 48442
rect 7116 48390 7130 48442
rect 7130 48390 7142 48442
rect 7142 48390 7172 48442
rect 7196 48390 7206 48442
rect 7206 48390 7252 48442
rect 6956 48388 7012 48390
rect 7036 48388 7092 48390
rect 7116 48388 7172 48390
rect 7196 48388 7252 48390
rect 6956 47354 7012 47356
rect 7036 47354 7092 47356
rect 7116 47354 7172 47356
rect 7196 47354 7252 47356
rect 6956 47302 7002 47354
rect 7002 47302 7012 47354
rect 7036 47302 7066 47354
rect 7066 47302 7078 47354
rect 7078 47302 7092 47354
rect 7116 47302 7130 47354
rect 7130 47302 7142 47354
rect 7142 47302 7172 47354
rect 7196 47302 7206 47354
rect 7206 47302 7252 47354
rect 6956 47300 7012 47302
rect 7036 47300 7092 47302
rect 7116 47300 7172 47302
rect 7196 47300 7252 47302
rect 6956 46266 7012 46268
rect 7036 46266 7092 46268
rect 7116 46266 7172 46268
rect 7196 46266 7252 46268
rect 6956 46214 7002 46266
rect 7002 46214 7012 46266
rect 7036 46214 7066 46266
rect 7066 46214 7078 46266
rect 7078 46214 7092 46266
rect 7116 46214 7130 46266
rect 7130 46214 7142 46266
rect 7142 46214 7172 46266
rect 7196 46214 7206 46266
rect 7206 46214 7252 46266
rect 6956 46212 7012 46214
rect 7036 46212 7092 46214
rect 7116 46212 7172 46214
rect 7196 46212 7252 46214
rect 6956 45178 7012 45180
rect 7036 45178 7092 45180
rect 7116 45178 7172 45180
rect 7196 45178 7252 45180
rect 6956 45126 7002 45178
rect 7002 45126 7012 45178
rect 7036 45126 7066 45178
rect 7066 45126 7078 45178
rect 7078 45126 7092 45178
rect 7116 45126 7130 45178
rect 7130 45126 7142 45178
rect 7142 45126 7172 45178
rect 7196 45126 7206 45178
rect 7206 45126 7252 45178
rect 6956 45124 7012 45126
rect 7036 45124 7092 45126
rect 7116 45124 7172 45126
rect 7196 45124 7252 45126
rect 6956 44090 7012 44092
rect 7036 44090 7092 44092
rect 7116 44090 7172 44092
rect 7196 44090 7252 44092
rect 6956 44038 7002 44090
rect 7002 44038 7012 44090
rect 7036 44038 7066 44090
rect 7066 44038 7078 44090
rect 7078 44038 7092 44090
rect 7116 44038 7130 44090
rect 7130 44038 7142 44090
rect 7142 44038 7172 44090
rect 7196 44038 7206 44090
rect 7206 44038 7252 44090
rect 6956 44036 7012 44038
rect 7036 44036 7092 44038
rect 7116 44036 7172 44038
rect 7196 44036 7252 44038
rect 6956 43002 7012 43004
rect 7036 43002 7092 43004
rect 7116 43002 7172 43004
rect 7196 43002 7252 43004
rect 6956 42950 7002 43002
rect 7002 42950 7012 43002
rect 7036 42950 7066 43002
rect 7066 42950 7078 43002
rect 7078 42950 7092 43002
rect 7116 42950 7130 43002
rect 7130 42950 7142 43002
rect 7142 42950 7172 43002
rect 7196 42950 7206 43002
rect 7206 42950 7252 43002
rect 6956 42948 7012 42950
rect 7036 42948 7092 42950
rect 7116 42948 7172 42950
rect 7196 42948 7252 42950
rect 6956 41914 7012 41916
rect 7036 41914 7092 41916
rect 7116 41914 7172 41916
rect 7196 41914 7252 41916
rect 6956 41862 7002 41914
rect 7002 41862 7012 41914
rect 7036 41862 7066 41914
rect 7066 41862 7078 41914
rect 7078 41862 7092 41914
rect 7116 41862 7130 41914
rect 7130 41862 7142 41914
rect 7142 41862 7172 41914
rect 7196 41862 7206 41914
rect 7206 41862 7252 41914
rect 6956 41860 7012 41862
rect 7036 41860 7092 41862
rect 7116 41860 7172 41862
rect 7196 41860 7252 41862
rect 6956 40826 7012 40828
rect 7036 40826 7092 40828
rect 7116 40826 7172 40828
rect 7196 40826 7252 40828
rect 6956 40774 7002 40826
rect 7002 40774 7012 40826
rect 7036 40774 7066 40826
rect 7066 40774 7078 40826
rect 7078 40774 7092 40826
rect 7116 40774 7130 40826
rect 7130 40774 7142 40826
rect 7142 40774 7172 40826
rect 7196 40774 7206 40826
rect 7206 40774 7252 40826
rect 6956 40772 7012 40774
rect 7036 40772 7092 40774
rect 7116 40772 7172 40774
rect 7196 40772 7252 40774
rect 6956 39738 7012 39740
rect 7036 39738 7092 39740
rect 7116 39738 7172 39740
rect 7196 39738 7252 39740
rect 6956 39686 7002 39738
rect 7002 39686 7012 39738
rect 7036 39686 7066 39738
rect 7066 39686 7078 39738
rect 7078 39686 7092 39738
rect 7116 39686 7130 39738
rect 7130 39686 7142 39738
rect 7142 39686 7172 39738
rect 7196 39686 7206 39738
rect 7206 39686 7252 39738
rect 6956 39684 7012 39686
rect 7036 39684 7092 39686
rect 7116 39684 7172 39686
rect 7196 39684 7252 39686
rect 6956 38650 7012 38652
rect 7036 38650 7092 38652
rect 7116 38650 7172 38652
rect 7196 38650 7252 38652
rect 6956 38598 7002 38650
rect 7002 38598 7012 38650
rect 7036 38598 7066 38650
rect 7066 38598 7078 38650
rect 7078 38598 7092 38650
rect 7116 38598 7130 38650
rect 7130 38598 7142 38650
rect 7142 38598 7172 38650
rect 7196 38598 7206 38650
rect 7206 38598 7252 38650
rect 6956 38596 7012 38598
rect 7036 38596 7092 38598
rect 7116 38596 7172 38598
rect 7196 38596 7252 38598
rect 6956 37562 7012 37564
rect 7036 37562 7092 37564
rect 7116 37562 7172 37564
rect 7196 37562 7252 37564
rect 6956 37510 7002 37562
rect 7002 37510 7012 37562
rect 7036 37510 7066 37562
rect 7066 37510 7078 37562
rect 7078 37510 7092 37562
rect 7116 37510 7130 37562
rect 7130 37510 7142 37562
rect 7142 37510 7172 37562
rect 7196 37510 7206 37562
rect 7206 37510 7252 37562
rect 6956 37508 7012 37510
rect 7036 37508 7092 37510
rect 7116 37508 7172 37510
rect 7196 37508 7252 37510
rect 6956 36474 7012 36476
rect 7036 36474 7092 36476
rect 7116 36474 7172 36476
rect 7196 36474 7252 36476
rect 6956 36422 7002 36474
rect 7002 36422 7012 36474
rect 7036 36422 7066 36474
rect 7066 36422 7078 36474
rect 7078 36422 7092 36474
rect 7116 36422 7130 36474
rect 7130 36422 7142 36474
rect 7142 36422 7172 36474
rect 7196 36422 7206 36474
rect 7206 36422 7252 36474
rect 6956 36420 7012 36422
rect 7036 36420 7092 36422
rect 7116 36420 7172 36422
rect 7196 36420 7252 36422
rect 6956 35386 7012 35388
rect 7036 35386 7092 35388
rect 7116 35386 7172 35388
rect 7196 35386 7252 35388
rect 6956 35334 7002 35386
rect 7002 35334 7012 35386
rect 7036 35334 7066 35386
rect 7066 35334 7078 35386
rect 7078 35334 7092 35386
rect 7116 35334 7130 35386
rect 7130 35334 7142 35386
rect 7142 35334 7172 35386
rect 7196 35334 7206 35386
rect 7206 35334 7252 35386
rect 6956 35332 7012 35334
rect 7036 35332 7092 35334
rect 7116 35332 7172 35334
rect 7196 35332 7252 35334
rect 6956 34298 7012 34300
rect 7036 34298 7092 34300
rect 7116 34298 7172 34300
rect 7196 34298 7252 34300
rect 6956 34246 7002 34298
rect 7002 34246 7012 34298
rect 7036 34246 7066 34298
rect 7066 34246 7078 34298
rect 7078 34246 7092 34298
rect 7116 34246 7130 34298
rect 7130 34246 7142 34298
rect 7142 34246 7172 34298
rect 7196 34246 7206 34298
rect 7206 34246 7252 34298
rect 6956 34244 7012 34246
rect 7036 34244 7092 34246
rect 7116 34244 7172 34246
rect 7196 34244 7252 34246
rect 6956 33210 7012 33212
rect 7036 33210 7092 33212
rect 7116 33210 7172 33212
rect 7196 33210 7252 33212
rect 6956 33158 7002 33210
rect 7002 33158 7012 33210
rect 7036 33158 7066 33210
rect 7066 33158 7078 33210
rect 7078 33158 7092 33210
rect 7116 33158 7130 33210
rect 7130 33158 7142 33210
rect 7142 33158 7172 33210
rect 7196 33158 7206 33210
rect 7206 33158 7252 33210
rect 6956 33156 7012 33158
rect 7036 33156 7092 33158
rect 7116 33156 7172 33158
rect 7196 33156 7252 33158
rect 6956 32122 7012 32124
rect 7036 32122 7092 32124
rect 7116 32122 7172 32124
rect 7196 32122 7252 32124
rect 6956 32070 7002 32122
rect 7002 32070 7012 32122
rect 7036 32070 7066 32122
rect 7066 32070 7078 32122
rect 7078 32070 7092 32122
rect 7116 32070 7130 32122
rect 7130 32070 7142 32122
rect 7142 32070 7172 32122
rect 7196 32070 7206 32122
rect 7206 32070 7252 32122
rect 6956 32068 7012 32070
rect 7036 32068 7092 32070
rect 7116 32068 7172 32070
rect 7196 32068 7252 32070
rect 6956 31034 7012 31036
rect 7036 31034 7092 31036
rect 7116 31034 7172 31036
rect 7196 31034 7252 31036
rect 6956 30982 7002 31034
rect 7002 30982 7012 31034
rect 7036 30982 7066 31034
rect 7066 30982 7078 31034
rect 7078 30982 7092 31034
rect 7116 30982 7130 31034
rect 7130 30982 7142 31034
rect 7142 30982 7172 31034
rect 7196 30982 7206 31034
rect 7206 30982 7252 31034
rect 6956 30980 7012 30982
rect 7036 30980 7092 30982
rect 7116 30980 7172 30982
rect 7196 30980 7252 30982
rect 6956 29946 7012 29948
rect 7036 29946 7092 29948
rect 7116 29946 7172 29948
rect 7196 29946 7252 29948
rect 6956 29894 7002 29946
rect 7002 29894 7012 29946
rect 7036 29894 7066 29946
rect 7066 29894 7078 29946
rect 7078 29894 7092 29946
rect 7116 29894 7130 29946
rect 7130 29894 7142 29946
rect 7142 29894 7172 29946
rect 7196 29894 7206 29946
rect 7206 29894 7252 29946
rect 6956 29892 7012 29894
rect 7036 29892 7092 29894
rect 7116 29892 7172 29894
rect 7196 29892 7252 29894
rect 6956 28858 7012 28860
rect 7036 28858 7092 28860
rect 7116 28858 7172 28860
rect 7196 28858 7252 28860
rect 6956 28806 7002 28858
rect 7002 28806 7012 28858
rect 7036 28806 7066 28858
rect 7066 28806 7078 28858
rect 7078 28806 7092 28858
rect 7116 28806 7130 28858
rect 7130 28806 7142 28858
rect 7142 28806 7172 28858
rect 7196 28806 7206 28858
rect 7206 28806 7252 28858
rect 6956 28804 7012 28806
rect 7036 28804 7092 28806
rect 7116 28804 7172 28806
rect 7196 28804 7252 28806
rect 6956 27770 7012 27772
rect 7036 27770 7092 27772
rect 7116 27770 7172 27772
rect 7196 27770 7252 27772
rect 6956 27718 7002 27770
rect 7002 27718 7012 27770
rect 7036 27718 7066 27770
rect 7066 27718 7078 27770
rect 7078 27718 7092 27770
rect 7116 27718 7130 27770
rect 7130 27718 7142 27770
rect 7142 27718 7172 27770
rect 7196 27718 7206 27770
rect 7206 27718 7252 27770
rect 6956 27716 7012 27718
rect 7036 27716 7092 27718
rect 7116 27716 7172 27718
rect 7196 27716 7252 27718
rect 6956 26682 7012 26684
rect 7036 26682 7092 26684
rect 7116 26682 7172 26684
rect 7196 26682 7252 26684
rect 6956 26630 7002 26682
rect 7002 26630 7012 26682
rect 7036 26630 7066 26682
rect 7066 26630 7078 26682
rect 7078 26630 7092 26682
rect 7116 26630 7130 26682
rect 7130 26630 7142 26682
rect 7142 26630 7172 26682
rect 7196 26630 7206 26682
rect 7206 26630 7252 26682
rect 6956 26628 7012 26630
rect 7036 26628 7092 26630
rect 7116 26628 7172 26630
rect 7196 26628 7252 26630
rect 6956 25594 7012 25596
rect 7036 25594 7092 25596
rect 7116 25594 7172 25596
rect 7196 25594 7252 25596
rect 6956 25542 7002 25594
rect 7002 25542 7012 25594
rect 7036 25542 7066 25594
rect 7066 25542 7078 25594
rect 7078 25542 7092 25594
rect 7116 25542 7130 25594
rect 7130 25542 7142 25594
rect 7142 25542 7172 25594
rect 7196 25542 7206 25594
rect 7206 25542 7252 25594
rect 6956 25540 7012 25542
rect 7036 25540 7092 25542
rect 7116 25540 7172 25542
rect 7196 25540 7252 25542
rect 7616 66394 7672 66396
rect 7696 66394 7752 66396
rect 7776 66394 7832 66396
rect 7856 66394 7912 66396
rect 7616 66342 7662 66394
rect 7662 66342 7672 66394
rect 7696 66342 7726 66394
rect 7726 66342 7738 66394
rect 7738 66342 7752 66394
rect 7776 66342 7790 66394
rect 7790 66342 7802 66394
rect 7802 66342 7832 66394
rect 7856 66342 7866 66394
rect 7866 66342 7912 66394
rect 7616 66340 7672 66342
rect 7696 66340 7752 66342
rect 7776 66340 7832 66342
rect 7856 66340 7912 66342
rect 8114 65456 8170 65512
rect 7616 65306 7672 65308
rect 7696 65306 7752 65308
rect 7776 65306 7832 65308
rect 7856 65306 7912 65308
rect 7616 65254 7662 65306
rect 7662 65254 7672 65306
rect 7696 65254 7726 65306
rect 7726 65254 7738 65306
rect 7738 65254 7752 65306
rect 7776 65254 7790 65306
rect 7790 65254 7802 65306
rect 7802 65254 7832 65306
rect 7856 65254 7866 65306
rect 7866 65254 7912 65306
rect 7616 65252 7672 65254
rect 7696 65252 7752 65254
rect 7776 65252 7832 65254
rect 7856 65252 7912 65254
rect 7616 64218 7672 64220
rect 7696 64218 7752 64220
rect 7776 64218 7832 64220
rect 7856 64218 7912 64220
rect 7616 64166 7662 64218
rect 7662 64166 7672 64218
rect 7696 64166 7726 64218
rect 7726 64166 7738 64218
rect 7738 64166 7752 64218
rect 7776 64166 7790 64218
rect 7790 64166 7802 64218
rect 7802 64166 7832 64218
rect 7856 64166 7866 64218
rect 7866 64166 7912 64218
rect 7616 64164 7672 64166
rect 7696 64164 7752 64166
rect 7776 64164 7832 64166
rect 7856 64164 7912 64166
rect 7616 63130 7672 63132
rect 7696 63130 7752 63132
rect 7776 63130 7832 63132
rect 7856 63130 7912 63132
rect 7616 63078 7662 63130
rect 7662 63078 7672 63130
rect 7696 63078 7726 63130
rect 7726 63078 7738 63130
rect 7738 63078 7752 63130
rect 7776 63078 7790 63130
rect 7790 63078 7802 63130
rect 7802 63078 7832 63130
rect 7856 63078 7866 63130
rect 7866 63078 7912 63130
rect 7616 63076 7672 63078
rect 7696 63076 7752 63078
rect 7776 63076 7832 63078
rect 7856 63076 7912 63078
rect 7616 62042 7672 62044
rect 7696 62042 7752 62044
rect 7776 62042 7832 62044
rect 7856 62042 7912 62044
rect 7616 61990 7662 62042
rect 7662 61990 7672 62042
rect 7696 61990 7726 62042
rect 7726 61990 7738 62042
rect 7738 61990 7752 62042
rect 7776 61990 7790 62042
rect 7790 61990 7802 62042
rect 7802 61990 7832 62042
rect 7856 61990 7866 62042
rect 7866 61990 7912 62042
rect 7616 61988 7672 61990
rect 7696 61988 7752 61990
rect 7776 61988 7832 61990
rect 7856 61988 7912 61990
rect 7616 60954 7672 60956
rect 7696 60954 7752 60956
rect 7776 60954 7832 60956
rect 7856 60954 7912 60956
rect 7616 60902 7662 60954
rect 7662 60902 7672 60954
rect 7696 60902 7726 60954
rect 7726 60902 7738 60954
rect 7738 60902 7752 60954
rect 7776 60902 7790 60954
rect 7790 60902 7802 60954
rect 7802 60902 7832 60954
rect 7856 60902 7866 60954
rect 7866 60902 7912 60954
rect 7616 60900 7672 60902
rect 7696 60900 7752 60902
rect 7776 60900 7832 60902
rect 7856 60900 7912 60902
rect 7616 59866 7672 59868
rect 7696 59866 7752 59868
rect 7776 59866 7832 59868
rect 7856 59866 7912 59868
rect 7616 59814 7662 59866
rect 7662 59814 7672 59866
rect 7696 59814 7726 59866
rect 7726 59814 7738 59866
rect 7738 59814 7752 59866
rect 7776 59814 7790 59866
rect 7790 59814 7802 59866
rect 7802 59814 7832 59866
rect 7856 59814 7866 59866
rect 7866 59814 7912 59866
rect 7616 59812 7672 59814
rect 7696 59812 7752 59814
rect 7776 59812 7832 59814
rect 7856 59812 7912 59814
rect 7616 58778 7672 58780
rect 7696 58778 7752 58780
rect 7776 58778 7832 58780
rect 7856 58778 7912 58780
rect 7616 58726 7662 58778
rect 7662 58726 7672 58778
rect 7696 58726 7726 58778
rect 7726 58726 7738 58778
rect 7738 58726 7752 58778
rect 7776 58726 7790 58778
rect 7790 58726 7802 58778
rect 7802 58726 7832 58778
rect 7856 58726 7866 58778
rect 7866 58726 7912 58778
rect 7616 58724 7672 58726
rect 7696 58724 7752 58726
rect 7776 58724 7832 58726
rect 7856 58724 7912 58726
rect 7616 57690 7672 57692
rect 7696 57690 7752 57692
rect 7776 57690 7832 57692
rect 7856 57690 7912 57692
rect 7616 57638 7662 57690
rect 7662 57638 7672 57690
rect 7696 57638 7726 57690
rect 7726 57638 7738 57690
rect 7738 57638 7752 57690
rect 7776 57638 7790 57690
rect 7790 57638 7802 57690
rect 7802 57638 7832 57690
rect 7856 57638 7866 57690
rect 7866 57638 7912 57690
rect 7616 57636 7672 57638
rect 7696 57636 7752 57638
rect 7776 57636 7832 57638
rect 7856 57636 7912 57638
rect 7616 56602 7672 56604
rect 7696 56602 7752 56604
rect 7776 56602 7832 56604
rect 7856 56602 7912 56604
rect 7616 56550 7662 56602
rect 7662 56550 7672 56602
rect 7696 56550 7726 56602
rect 7726 56550 7738 56602
rect 7738 56550 7752 56602
rect 7776 56550 7790 56602
rect 7790 56550 7802 56602
rect 7802 56550 7832 56602
rect 7856 56550 7866 56602
rect 7866 56550 7912 56602
rect 7616 56548 7672 56550
rect 7696 56548 7752 56550
rect 7776 56548 7832 56550
rect 7856 56548 7912 56550
rect 7616 55514 7672 55516
rect 7696 55514 7752 55516
rect 7776 55514 7832 55516
rect 7856 55514 7912 55516
rect 7616 55462 7662 55514
rect 7662 55462 7672 55514
rect 7696 55462 7726 55514
rect 7726 55462 7738 55514
rect 7738 55462 7752 55514
rect 7776 55462 7790 55514
rect 7790 55462 7802 55514
rect 7802 55462 7832 55514
rect 7856 55462 7866 55514
rect 7866 55462 7912 55514
rect 7616 55460 7672 55462
rect 7696 55460 7752 55462
rect 7776 55460 7832 55462
rect 7856 55460 7912 55462
rect 7616 54426 7672 54428
rect 7696 54426 7752 54428
rect 7776 54426 7832 54428
rect 7856 54426 7912 54428
rect 7616 54374 7662 54426
rect 7662 54374 7672 54426
rect 7696 54374 7726 54426
rect 7726 54374 7738 54426
rect 7738 54374 7752 54426
rect 7776 54374 7790 54426
rect 7790 54374 7802 54426
rect 7802 54374 7832 54426
rect 7856 54374 7866 54426
rect 7866 54374 7912 54426
rect 7616 54372 7672 54374
rect 7696 54372 7752 54374
rect 7776 54372 7832 54374
rect 7856 54372 7912 54374
rect 7616 53338 7672 53340
rect 7696 53338 7752 53340
rect 7776 53338 7832 53340
rect 7856 53338 7912 53340
rect 7616 53286 7662 53338
rect 7662 53286 7672 53338
rect 7696 53286 7726 53338
rect 7726 53286 7738 53338
rect 7738 53286 7752 53338
rect 7776 53286 7790 53338
rect 7790 53286 7802 53338
rect 7802 53286 7832 53338
rect 7856 53286 7866 53338
rect 7866 53286 7912 53338
rect 7616 53284 7672 53286
rect 7696 53284 7752 53286
rect 7776 53284 7832 53286
rect 7856 53284 7912 53286
rect 7616 52250 7672 52252
rect 7696 52250 7752 52252
rect 7776 52250 7832 52252
rect 7856 52250 7912 52252
rect 7616 52198 7662 52250
rect 7662 52198 7672 52250
rect 7696 52198 7726 52250
rect 7726 52198 7738 52250
rect 7738 52198 7752 52250
rect 7776 52198 7790 52250
rect 7790 52198 7802 52250
rect 7802 52198 7832 52250
rect 7856 52198 7866 52250
rect 7866 52198 7912 52250
rect 7616 52196 7672 52198
rect 7696 52196 7752 52198
rect 7776 52196 7832 52198
rect 7856 52196 7912 52198
rect 7616 51162 7672 51164
rect 7696 51162 7752 51164
rect 7776 51162 7832 51164
rect 7856 51162 7912 51164
rect 7616 51110 7662 51162
rect 7662 51110 7672 51162
rect 7696 51110 7726 51162
rect 7726 51110 7738 51162
rect 7738 51110 7752 51162
rect 7776 51110 7790 51162
rect 7790 51110 7802 51162
rect 7802 51110 7832 51162
rect 7856 51110 7866 51162
rect 7866 51110 7912 51162
rect 7616 51108 7672 51110
rect 7696 51108 7752 51110
rect 7776 51108 7832 51110
rect 7856 51108 7912 51110
rect 11956 69114 12012 69116
rect 12036 69114 12092 69116
rect 12116 69114 12172 69116
rect 12196 69114 12252 69116
rect 11956 69062 12002 69114
rect 12002 69062 12012 69114
rect 12036 69062 12066 69114
rect 12066 69062 12078 69114
rect 12078 69062 12092 69114
rect 12116 69062 12130 69114
rect 12130 69062 12142 69114
rect 12142 69062 12172 69114
rect 12196 69062 12206 69114
rect 12206 69062 12252 69114
rect 11956 69060 12012 69062
rect 12036 69060 12092 69062
rect 12116 69060 12172 69062
rect 12196 69060 12252 69062
rect 16956 69114 17012 69116
rect 17036 69114 17092 69116
rect 17116 69114 17172 69116
rect 17196 69114 17252 69116
rect 16956 69062 17002 69114
rect 17002 69062 17012 69114
rect 17036 69062 17066 69114
rect 17066 69062 17078 69114
rect 17078 69062 17092 69114
rect 17116 69062 17130 69114
rect 17130 69062 17142 69114
rect 17142 69062 17172 69114
rect 17196 69062 17206 69114
rect 17206 69062 17252 69114
rect 16956 69060 17012 69062
rect 17036 69060 17092 69062
rect 17116 69060 17172 69062
rect 17196 69060 17252 69062
rect 21956 69114 22012 69116
rect 22036 69114 22092 69116
rect 22116 69114 22172 69116
rect 22196 69114 22252 69116
rect 21956 69062 22002 69114
rect 22002 69062 22012 69114
rect 22036 69062 22066 69114
rect 22066 69062 22078 69114
rect 22078 69062 22092 69114
rect 22116 69062 22130 69114
rect 22130 69062 22142 69114
rect 22142 69062 22172 69114
rect 22196 69062 22206 69114
rect 22206 69062 22252 69114
rect 21956 69060 22012 69062
rect 22036 69060 22092 69062
rect 22116 69060 22172 69062
rect 22196 69060 22252 69062
rect 7616 50074 7672 50076
rect 7696 50074 7752 50076
rect 7776 50074 7832 50076
rect 7856 50074 7912 50076
rect 7616 50022 7662 50074
rect 7662 50022 7672 50074
rect 7696 50022 7726 50074
rect 7726 50022 7738 50074
rect 7738 50022 7752 50074
rect 7776 50022 7790 50074
rect 7790 50022 7802 50074
rect 7802 50022 7832 50074
rect 7856 50022 7866 50074
rect 7866 50022 7912 50074
rect 7616 50020 7672 50022
rect 7696 50020 7752 50022
rect 7776 50020 7832 50022
rect 7856 50020 7912 50022
rect 7616 48986 7672 48988
rect 7696 48986 7752 48988
rect 7776 48986 7832 48988
rect 7856 48986 7912 48988
rect 7616 48934 7662 48986
rect 7662 48934 7672 48986
rect 7696 48934 7726 48986
rect 7726 48934 7738 48986
rect 7738 48934 7752 48986
rect 7776 48934 7790 48986
rect 7790 48934 7802 48986
rect 7802 48934 7832 48986
rect 7856 48934 7866 48986
rect 7866 48934 7912 48986
rect 7616 48932 7672 48934
rect 7696 48932 7752 48934
rect 7776 48932 7832 48934
rect 7856 48932 7912 48934
rect 7616 47898 7672 47900
rect 7696 47898 7752 47900
rect 7776 47898 7832 47900
rect 7856 47898 7912 47900
rect 7616 47846 7662 47898
rect 7662 47846 7672 47898
rect 7696 47846 7726 47898
rect 7726 47846 7738 47898
rect 7738 47846 7752 47898
rect 7776 47846 7790 47898
rect 7790 47846 7802 47898
rect 7802 47846 7832 47898
rect 7856 47846 7866 47898
rect 7866 47846 7912 47898
rect 7616 47844 7672 47846
rect 7696 47844 7752 47846
rect 7776 47844 7832 47846
rect 7856 47844 7912 47846
rect 7616 46810 7672 46812
rect 7696 46810 7752 46812
rect 7776 46810 7832 46812
rect 7856 46810 7912 46812
rect 7616 46758 7662 46810
rect 7662 46758 7672 46810
rect 7696 46758 7726 46810
rect 7726 46758 7738 46810
rect 7738 46758 7752 46810
rect 7776 46758 7790 46810
rect 7790 46758 7802 46810
rect 7802 46758 7832 46810
rect 7856 46758 7866 46810
rect 7866 46758 7912 46810
rect 7616 46756 7672 46758
rect 7696 46756 7752 46758
rect 7776 46756 7832 46758
rect 7856 46756 7912 46758
rect 7616 45722 7672 45724
rect 7696 45722 7752 45724
rect 7776 45722 7832 45724
rect 7856 45722 7912 45724
rect 7616 45670 7662 45722
rect 7662 45670 7672 45722
rect 7696 45670 7726 45722
rect 7726 45670 7738 45722
rect 7738 45670 7752 45722
rect 7776 45670 7790 45722
rect 7790 45670 7802 45722
rect 7802 45670 7832 45722
rect 7856 45670 7866 45722
rect 7866 45670 7912 45722
rect 7616 45668 7672 45670
rect 7696 45668 7752 45670
rect 7776 45668 7832 45670
rect 7856 45668 7912 45670
rect 7616 44634 7672 44636
rect 7696 44634 7752 44636
rect 7776 44634 7832 44636
rect 7856 44634 7912 44636
rect 7616 44582 7662 44634
rect 7662 44582 7672 44634
rect 7696 44582 7726 44634
rect 7726 44582 7738 44634
rect 7738 44582 7752 44634
rect 7776 44582 7790 44634
rect 7790 44582 7802 44634
rect 7802 44582 7832 44634
rect 7856 44582 7866 44634
rect 7866 44582 7912 44634
rect 7616 44580 7672 44582
rect 7696 44580 7752 44582
rect 7776 44580 7832 44582
rect 7856 44580 7912 44582
rect 7616 43546 7672 43548
rect 7696 43546 7752 43548
rect 7776 43546 7832 43548
rect 7856 43546 7912 43548
rect 7616 43494 7662 43546
rect 7662 43494 7672 43546
rect 7696 43494 7726 43546
rect 7726 43494 7738 43546
rect 7738 43494 7752 43546
rect 7776 43494 7790 43546
rect 7790 43494 7802 43546
rect 7802 43494 7832 43546
rect 7856 43494 7866 43546
rect 7866 43494 7912 43546
rect 7616 43492 7672 43494
rect 7696 43492 7752 43494
rect 7776 43492 7832 43494
rect 7856 43492 7912 43494
rect 7616 42458 7672 42460
rect 7696 42458 7752 42460
rect 7776 42458 7832 42460
rect 7856 42458 7912 42460
rect 7616 42406 7662 42458
rect 7662 42406 7672 42458
rect 7696 42406 7726 42458
rect 7726 42406 7738 42458
rect 7738 42406 7752 42458
rect 7776 42406 7790 42458
rect 7790 42406 7802 42458
rect 7802 42406 7832 42458
rect 7856 42406 7866 42458
rect 7866 42406 7912 42458
rect 7616 42404 7672 42406
rect 7696 42404 7752 42406
rect 7776 42404 7832 42406
rect 7856 42404 7912 42406
rect 7616 41370 7672 41372
rect 7696 41370 7752 41372
rect 7776 41370 7832 41372
rect 7856 41370 7912 41372
rect 7616 41318 7662 41370
rect 7662 41318 7672 41370
rect 7696 41318 7726 41370
rect 7726 41318 7738 41370
rect 7738 41318 7752 41370
rect 7776 41318 7790 41370
rect 7790 41318 7802 41370
rect 7802 41318 7832 41370
rect 7856 41318 7866 41370
rect 7866 41318 7912 41370
rect 7616 41316 7672 41318
rect 7696 41316 7752 41318
rect 7776 41316 7832 41318
rect 7856 41316 7912 41318
rect 7616 40282 7672 40284
rect 7696 40282 7752 40284
rect 7776 40282 7832 40284
rect 7856 40282 7912 40284
rect 7616 40230 7662 40282
rect 7662 40230 7672 40282
rect 7696 40230 7726 40282
rect 7726 40230 7738 40282
rect 7738 40230 7752 40282
rect 7776 40230 7790 40282
rect 7790 40230 7802 40282
rect 7802 40230 7832 40282
rect 7856 40230 7866 40282
rect 7866 40230 7912 40282
rect 7616 40228 7672 40230
rect 7696 40228 7752 40230
rect 7776 40228 7832 40230
rect 7856 40228 7912 40230
rect 7616 39194 7672 39196
rect 7696 39194 7752 39196
rect 7776 39194 7832 39196
rect 7856 39194 7912 39196
rect 7616 39142 7662 39194
rect 7662 39142 7672 39194
rect 7696 39142 7726 39194
rect 7726 39142 7738 39194
rect 7738 39142 7752 39194
rect 7776 39142 7790 39194
rect 7790 39142 7802 39194
rect 7802 39142 7832 39194
rect 7856 39142 7866 39194
rect 7866 39142 7912 39194
rect 7616 39140 7672 39142
rect 7696 39140 7752 39142
rect 7776 39140 7832 39142
rect 7856 39140 7912 39142
rect 7616 38106 7672 38108
rect 7696 38106 7752 38108
rect 7776 38106 7832 38108
rect 7856 38106 7912 38108
rect 7616 38054 7662 38106
rect 7662 38054 7672 38106
rect 7696 38054 7726 38106
rect 7726 38054 7738 38106
rect 7738 38054 7752 38106
rect 7776 38054 7790 38106
rect 7790 38054 7802 38106
rect 7802 38054 7832 38106
rect 7856 38054 7866 38106
rect 7866 38054 7912 38106
rect 7616 38052 7672 38054
rect 7696 38052 7752 38054
rect 7776 38052 7832 38054
rect 7856 38052 7912 38054
rect 7616 37018 7672 37020
rect 7696 37018 7752 37020
rect 7776 37018 7832 37020
rect 7856 37018 7912 37020
rect 7616 36966 7662 37018
rect 7662 36966 7672 37018
rect 7696 36966 7726 37018
rect 7726 36966 7738 37018
rect 7738 36966 7752 37018
rect 7776 36966 7790 37018
rect 7790 36966 7802 37018
rect 7802 36966 7832 37018
rect 7856 36966 7866 37018
rect 7866 36966 7912 37018
rect 7616 36964 7672 36966
rect 7696 36964 7752 36966
rect 7776 36964 7832 36966
rect 7856 36964 7912 36966
rect 7616 35930 7672 35932
rect 7696 35930 7752 35932
rect 7776 35930 7832 35932
rect 7856 35930 7912 35932
rect 7616 35878 7662 35930
rect 7662 35878 7672 35930
rect 7696 35878 7726 35930
rect 7726 35878 7738 35930
rect 7738 35878 7752 35930
rect 7776 35878 7790 35930
rect 7790 35878 7802 35930
rect 7802 35878 7832 35930
rect 7856 35878 7866 35930
rect 7866 35878 7912 35930
rect 7616 35876 7672 35878
rect 7696 35876 7752 35878
rect 7776 35876 7832 35878
rect 7856 35876 7912 35878
rect 7378 34720 7434 34776
rect 7616 34842 7672 34844
rect 7696 34842 7752 34844
rect 7776 34842 7832 34844
rect 7856 34842 7912 34844
rect 7616 34790 7662 34842
rect 7662 34790 7672 34842
rect 7696 34790 7726 34842
rect 7726 34790 7738 34842
rect 7738 34790 7752 34842
rect 7776 34790 7790 34842
rect 7790 34790 7802 34842
rect 7802 34790 7832 34842
rect 7856 34790 7866 34842
rect 7866 34790 7912 34842
rect 7616 34788 7672 34790
rect 7696 34788 7752 34790
rect 7776 34788 7832 34790
rect 7856 34788 7912 34790
rect 7470 34448 7526 34504
rect 7616 33754 7672 33756
rect 7696 33754 7752 33756
rect 7776 33754 7832 33756
rect 7856 33754 7912 33756
rect 7616 33702 7662 33754
rect 7662 33702 7672 33754
rect 7696 33702 7726 33754
rect 7726 33702 7738 33754
rect 7738 33702 7752 33754
rect 7776 33702 7790 33754
rect 7790 33702 7802 33754
rect 7802 33702 7832 33754
rect 7856 33702 7866 33754
rect 7866 33702 7912 33754
rect 7616 33700 7672 33702
rect 7696 33700 7752 33702
rect 7776 33700 7832 33702
rect 7856 33700 7912 33702
rect 7616 32666 7672 32668
rect 7696 32666 7752 32668
rect 7776 32666 7832 32668
rect 7856 32666 7912 32668
rect 7616 32614 7662 32666
rect 7662 32614 7672 32666
rect 7696 32614 7726 32666
rect 7726 32614 7738 32666
rect 7738 32614 7752 32666
rect 7776 32614 7790 32666
rect 7790 32614 7802 32666
rect 7802 32614 7832 32666
rect 7856 32614 7866 32666
rect 7866 32614 7912 32666
rect 7616 32612 7672 32614
rect 7696 32612 7752 32614
rect 7776 32612 7832 32614
rect 7856 32612 7912 32614
rect 6956 24506 7012 24508
rect 7036 24506 7092 24508
rect 7116 24506 7172 24508
rect 7196 24506 7252 24508
rect 6956 24454 7002 24506
rect 7002 24454 7012 24506
rect 7036 24454 7066 24506
rect 7066 24454 7078 24506
rect 7078 24454 7092 24506
rect 7116 24454 7130 24506
rect 7130 24454 7142 24506
rect 7142 24454 7172 24506
rect 7196 24454 7206 24506
rect 7206 24454 7252 24506
rect 6956 24452 7012 24454
rect 7036 24452 7092 24454
rect 7116 24452 7172 24454
rect 7196 24452 7252 24454
rect 6956 23418 7012 23420
rect 7036 23418 7092 23420
rect 7116 23418 7172 23420
rect 7196 23418 7252 23420
rect 6956 23366 7002 23418
rect 7002 23366 7012 23418
rect 7036 23366 7066 23418
rect 7066 23366 7078 23418
rect 7078 23366 7092 23418
rect 7116 23366 7130 23418
rect 7130 23366 7142 23418
rect 7142 23366 7172 23418
rect 7196 23366 7206 23418
rect 7206 23366 7252 23418
rect 6956 23364 7012 23366
rect 7036 23364 7092 23366
rect 7116 23364 7172 23366
rect 7196 23364 7252 23366
rect 6956 22330 7012 22332
rect 7036 22330 7092 22332
rect 7116 22330 7172 22332
rect 7196 22330 7252 22332
rect 6956 22278 7002 22330
rect 7002 22278 7012 22330
rect 7036 22278 7066 22330
rect 7066 22278 7078 22330
rect 7078 22278 7092 22330
rect 7116 22278 7130 22330
rect 7130 22278 7142 22330
rect 7142 22278 7172 22330
rect 7196 22278 7206 22330
rect 7206 22278 7252 22330
rect 6956 22276 7012 22278
rect 7036 22276 7092 22278
rect 7116 22276 7172 22278
rect 7196 22276 7252 22278
rect 6956 21242 7012 21244
rect 7036 21242 7092 21244
rect 7116 21242 7172 21244
rect 7196 21242 7252 21244
rect 6956 21190 7002 21242
rect 7002 21190 7012 21242
rect 7036 21190 7066 21242
rect 7066 21190 7078 21242
rect 7078 21190 7092 21242
rect 7116 21190 7130 21242
rect 7130 21190 7142 21242
rect 7142 21190 7172 21242
rect 7196 21190 7206 21242
rect 7206 21190 7252 21242
rect 6956 21188 7012 21190
rect 7036 21188 7092 21190
rect 7116 21188 7172 21190
rect 7196 21188 7252 21190
rect 6956 20154 7012 20156
rect 7036 20154 7092 20156
rect 7116 20154 7172 20156
rect 7196 20154 7252 20156
rect 6956 20102 7002 20154
rect 7002 20102 7012 20154
rect 7036 20102 7066 20154
rect 7066 20102 7078 20154
rect 7078 20102 7092 20154
rect 7116 20102 7130 20154
rect 7130 20102 7142 20154
rect 7142 20102 7172 20154
rect 7196 20102 7206 20154
rect 7206 20102 7252 20154
rect 6956 20100 7012 20102
rect 7036 20100 7092 20102
rect 7116 20100 7172 20102
rect 7196 20100 7252 20102
rect 6956 19066 7012 19068
rect 7036 19066 7092 19068
rect 7116 19066 7172 19068
rect 7196 19066 7252 19068
rect 6956 19014 7002 19066
rect 7002 19014 7012 19066
rect 7036 19014 7066 19066
rect 7066 19014 7078 19066
rect 7078 19014 7092 19066
rect 7116 19014 7130 19066
rect 7130 19014 7142 19066
rect 7142 19014 7172 19066
rect 7196 19014 7206 19066
rect 7206 19014 7252 19066
rect 6956 19012 7012 19014
rect 7036 19012 7092 19014
rect 7116 19012 7172 19014
rect 7196 19012 7252 19014
rect 6956 17978 7012 17980
rect 7036 17978 7092 17980
rect 7116 17978 7172 17980
rect 7196 17978 7252 17980
rect 6956 17926 7002 17978
rect 7002 17926 7012 17978
rect 7036 17926 7066 17978
rect 7066 17926 7078 17978
rect 7078 17926 7092 17978
rect 7116 17926 7130 17978
rect 7130 17926 7142 17978
rect 7142 17926 7172 17978
rect 7196 17926 7206 17978
rect 7206 17926 7252 17978
rect 6956 17924 7012 17926
rect 7036 17924 7092 17926
rect 7116 17924 7172 17926
rect 7196 17924 7252 17926
rect 6956 16890 7012 16892
rect 7036 16890 7092 16892
rect 7116 16890 7172 16892
rect 7196 16890 7252 16892
rect 6956 16838 7002 16890
rect 7002 16838 7012 16890
rect 7036 16838 7066 16890
rect 7066 16838 7078 16890
rect 7078 16838 7092 16890
rect 7116 16838 7130 16890
rect 7130 16838 7142 16890
rect 7142 16838 7172 16890
rect 7196 16838 7206 16890
rect 7206 16838 7252 16890
rect 6956 16836 7012 16838
rect 7036 16836 7092 16838
rect 7116 16836 7172 16838
rect 7196 16836 7252 16838
rect 6956 15802 7012 15804
rect 7036 15802 7092 15804
rect 7116 15802 7172 15804
rect 7196 15802 7252 15804
rect 6956 15750 7002 15802
rect 7002 15750 7012 15802
rect 7036 15750 7066 15802
rect 7066 15750 7078 15802
rect 7078 15750 7092 15802
rect 7116 15750 7130 15802
rect 7130 15750 7142 15802
rect 7142 15750 7172 15802
rect 7196 15750 7206 15802
rect 7206 15750 7252 15802
rect 6956 15748 7012 15750
rect 7036 15748 7092 15750
rect 7116 15748 7172 15750
rect 7196 15748 7252 15750
rect 6956 14714 7012 14716
rect 7036 14714 7092 14716
rect 7116 14714 7172 14716
rect 7196 14714 7252 14716
rect 6956 14662 7002 14714
rect 7002 14662 7012 14714
rect 7036 14662 7066 14714
rect 7066 14662 7078 14714
rect 7078 14662 7092 14714
rect 7116 14662 7130 14714
rect 7130 14662 7142 14714
rect 7142 14662 7172 14714
rect 7196 14662 7206 14714
rect 7206 14662 7252 14714
rect 6956 14660 7012 14662
rect 7036 14660 7092 14662
rect 7116 14660 7172 14662
rect 7196 14660 7252 14662
rect 6956 13626 7012 13628
rect 7036 13626 7092 13628
rect 7116 13626 7172 13628
rect 7196 13626 7252 13628
rect 6956 13574 7002 13626
rect 7002 13574 7012 13626
rect 7036 13574 7066 13626
rect 7066 13574 7078 13626
rect 7078 13574 7092 13626
rect 7116 13574 7130 13626
rect 7130 13574 7142 13626
rect 7142 13574 7172 13626
rect 7196 13574 7206 13626
rect 7206 13574 7252 13626
rect 6956 13572 7012 13574
rect 7036 13572 7092 13574
rect 7116 13572 7172 13574
rect 7196 13572 7252 13574
rect 6956 12538 7012 12540
rect 7036 12538 7092 12540
rect 7116 12538 7172 12540
rect 7196 12538 7252 12540
rect 6956 12486 7002 12538
rect 7002 12486 7012 12538
rect 7036 12486 7066 12538
rect 7066 12486 7078 12538
rect 7078 12486 7092 12538
rect 7116 12486 7130 12538
rect 7130 12486 7142 12538
rect 7142 12486 7172 12538
rect 7196 12486 7206 12538
rect 7206 12486 7252 12538
rect 6956 12484 7012 12486
rect 7036 12484 7092 12486
rect 7116 12484 7172 12486
rect 7196 12484 7252 12486
rect 6956 11450 7012 11452
rect 7036 11450 7092 11452
rect 7116 11450 7172 11452
rect 7196 11450 7252 11452
rect 6956 11398 7002 11450
rect 7002 11398 7012 11450
rect 7036 11398 7066 11450
rect 7066 11398 7078 11450
rect 7078 11398 7092 11450
rect 7116 11398 7130 11450
rect 7130 11398 7142 11450
rect 7142 11398 7172 11450
rect 7196 11398 7206 11450
rect 7206 11398 7252 11450
rect 6956 11396 7012 11398
rect 7036 11396 7092 11398
rect 7116 11396 7172 11398
rect 7196 11396 7252 11398
rect 6956 10362 7012 10364
rect 7036 10362 7092 10364
rect 7116 10362 7172 10364
rect 7196 10362 7252 10364
rect 6956 10310 7002 10362
rect 7002 10310 7012 10362
rect 7036 10310 7066 10362
rect 7066 10310 7078 10362
rect 7078 10310 7092 10362
rect 7116 10310 7130 10362
rect 7130 10310 7142 10362
rect 7142 10310 7172 10362
rect 7196 10310 7206 10362
rect 7206 10310 7252 10362
rect 6956 10308 7012 10310
rect 7036 10308 7092 10310
rect 7116 10308 7172 10310
rect 7196 10308 7252 10310
rect 6956 9274 7012 9276
rect 7036 9274 7092 9276
rect 7116 9274 7172 9276
rect 7196 9274 7252 9276
rect 6956 9222 7002 9274
rect 7002 9222 7012 9274
rect 7036 9222 7066 9274
rect 7066 9222 7078 9274
rect 7078 9222 7092 9274
rect 7116 9222 7130 9274
rect 7130 9222 7142 9274
rect 7142 9222 7172 9274
rect 7196 9222 7206 9274
rect 7206 9222 7252 9274
rect 6956 9220 7012 9222
rect 7036 9220 7092 9222
rect 7116 9220 7172 9222
rect 7196 9220 7252 9222
rect 6956 8186 7012 8188
rect 7036 8186 7092 8188
rect 7116 8186 7172 8188
rect 7196 8186 7252 8188
rect 6956 8134 7002 8186
rect 7002 8134 7012 8186
rect 7036 8134 7066 8186
rect 7066 8134 7078 8186
rect 7078 8134 7092 8186
rect 7116 8134 7130 8186
rect 7130 8134 7142 8186
rect 7142 8134 7172 8186
rect 7196 8134 7206 8186
rect 7206 8134 7252 8186
rect 6956 8132 7012 8134
rect 7036 8132 7092 8134
rect 7116 8132 7172 8134
rect 7196 8132 7252 8134
rect 6956 7098 7012 7100
rect 7036 7098 7092 7100
rect 7116 7098 7172 7100
rect 7196 7098 7252 7100
rect 6956 7046 7002 7098
rect 7002 7046 7012 7098
rect 7036 7046 7066 7098
rect 7066 7046 7078 7098
rect 7078 7046 7092 7098
rect 7116 7046 7130 7098
rect 7130 7046 7142 7098
rect 7142 7046 7172 7098
rect 7196 7046 7206 7098
rect 7206 7046 7252 7098
rect 6956 7044 7012 7046
rect 7036 7044 7092 7046
rect 7116 7044 7172 7046
rect 7196 7044 7252 7046
rect 6956 6010 7012 6012
rect 7036 6010 7092 6012
rect 7116 6010 7172 6012
rect 7196 6010 7252 6012
rect 6956 5958 7002 6010
rect 7002 5958 7012 6010
rect 7036 5958 7066 6010
rect 7066 5958 7078 6010
rect 7078 5958 7092 6010
rect 7116 5958 7130 6010
rect 7130 5958 7142 6010
rect 7142 5958 7172 6010
rect 7196 5958 7206 6010
rect 7206 5958 7252 6010
rect 6956 5956 7012 5958
rect 7036 5956 7092 5958
rect 7116 5956 7172 5958
rect 7196 5956 7252 5958
rect 7616 31578 7672 31580
rect 7696 31578 7752 31580
rect 7776 31578 7832 31580
rect 7856 31578 7912 31580
rect 7616 31526 7662 31578
rect 7662 31526 7672 31578
rect 7696 31526 7726 31578
rect 7726 31526 7738 31578
rect 7738 31526 7752 31578
rect 7776 31526 7790 31578
rect 7790 31526 7802 31578
rect 7802 31526 7832 31578
rect 7856 31526 7866 31578
rect 7866 31526 7912 31578
rect 7616 31524 7672 31526
rect 7696 31524 7752 31526
rect 7776 31524 7832 31526
rect 7856 31524 7912 31526
rect 7616 30490 7672 30492
rect 7696 30490 7752 30492
rect 7776 30490 7832 30492
rect 7856 30490 7912 30492
rect 7616 30438 7662 30490
rect 7662 30438 7672 30490
rect 7696 30438 7726 30490
rect 7726 30438 7738 30490
rect 7738 30438 7752 30490
rect 7776 30438 7790 30490
rect 7790 30438 7802 30490
rect 7802 30438 7832 30490
rect 7856 30438 7866 30490
rect 7866 30438 7912 30490
rect 7616 30436 7672 30438
rect 7696 30436 7752 30438
rect 7776 30436 7832 30438
rect 7856 30436 7912 30438
rect 7616 29402 7672 29404
rect 7696 29402 7752 29404
rect 7776 29402 7832 29404
rect 7856 29402 7912 29404
rect 7616 29350 7662 29402
rect 7662 29350 7672 29402
rect 7696 29350 7726 29402
rect 7726 29350 7738 29402
rect 7738 29350 7752 29402
rect 7776 29350 7790 29402
rect 7790 29350 7802 29402
rect 7802 29350 7832 29402
rect 7856 29350 7866 29402
rect 7866 29350 7912 29402
rect 7616 29348 7672 29350
rect 7696 29348 7752 29350
rect 7776 29348 7832 29350
rect 7856 29348 7912 29350
rect 7616 28314 7672 28316
rect 7696 28314 7752 28316
rect 7776 28314 7832 28316
rect 7856 28314 7912 28316
rect 7616 28262 7662 28314
rect 7662 28262 7672 28314
rect 7696 28262 7726 28314
rect 7726 28262 7738 28314
rect 7738 28262 7752 28314
rect 7776 28262 7790 28314
rect 7790 28262 7802 28314
rect 7802 28262 7832 28314
rect 7856 28262 7866 28314
rect 7866 28262 7912 28314
rect 7616 28260 7672 28262
rect 7696 28260 7752 28262
rect 7776 28260 7832 28262
rect 7856 28260 7912 28262
rect 7616 27226 7672 27228
rect 7696 27226 7752 27228
rect 7776 27226 7832 27228
rect 7856 27226 7912 27228
rect 7616 27174 7662 27226
rect 7662 27174 7672 27226
rect 7696 27174 7726 27226
rect 7726 27174 7738 27226
rect 7738 27174 7752 27226
rect 7776 27174 7790 27226
rect 7790 27174 7802 27226
rect 7802 27174 7832 27226
rect 7856 27174 7866 27226
rect 7866 27174 7912 27226
rect 7616 27172 7672 27174
rect 7696 27172 7752 27174
rect 7776 27172 7832 27174
rect 7856 27172 7912 27174
rect 7616 26138 7672 26140
rect 7696 26138 7752 26140
rect 7776 26138 7832 26140
rect 7856 26138 7912 26140
rect 7616 26086 7662 26138
rect 7662 26086 7672 26138
rect 7696 26086 7726 26138
rect 7726 26086 7738 26138
rect 7738 26086 7752 26138
rect 7776 26086 7790 26138
rect 7790 26086 7802 26138
rect 7802 26086 7832 26138
rect 7856 26086 7866 26138
rect 7866 26086 7912 26138
rect 7616 26084 7672 26086
rect 7696 26084 7752 26086
rect 7776 26084 7832 26086
rect 7856 26084 7912 26086
rect 7616 25050 7672 25052
rect 7696 25050 7752 25052
rect 7776 25050 7832 25052
rect 7856 25050 7912 25052
rect 7616 24998 7662 25050
rect 7662 24998 7672 25050
rect 7696 24998 7726 25050
rect 7726 24998 7738 25050
rect 7738 24998 7752 25050
rect 7776 24998 7790 25050
rect 7790 24998 7802 25050
rect 7802 24998 7832 25050
rect 7856 24998 7866 25050
rect 7866 24998 7912 25050
rect 7616 24996 7672 24998
rect 7696 24996 7752 24998
rect 7776 24996 7832 24998
rect 7856 24996 7912 24998
rect 8206 34992 8262 35048
rect 8206 34720 8262 34776
rect 7616 23962 7672 23964
rect 7696 23962 7752 23964
rect 7776 23962 7832 23964
rect 7856 23962 7912 23964
rect 7616 23910 7662 23962
rect 7662 23910 7672 23962
rect 7696 23910 7726 23962
rect 7726 23910 7738 23962
rect 7738 23910 7752 23962
rect 7776 23910 7790 23962
rect 7790 23910 7802 23962
rect 7802 23910 7832 23962
rect 7856 23910 7866 23962
rect 7866 23910 7912 23962
rect 7616 23908 7672 23910
rect 7696 23908 7752 23910
rect 7776 23908 7832 23910
rect 7856 23908 7912 23910
rect 7616 22874 7672 22876
rect 7696 22874 7752 22876
rect 7776 22874 7832 22876
rect 7856 22874 7912 22876
rect 7616 22822 7662 22874
rect 7662 22822 7672 22874
rect 7696 22822 7726 22874
rect 7726 22822 7738 22874
rect 7738 22822 7752 22874
rect 7776 22822 7790 22874
rect 7790 22822 7802 22874
rect 7802 22822 7832 22874
rect 7856 22822 7866 22874
rect 7866 22822 7912 22874
rect 7616 22820 7672 22822
rect 7696 22820 7752 22822
rect 7776 22820 7832 22822
rect 7856 22820 7912 22822
rect 7616 21786 7672 21788
rect 7696 21786 7752 21788
rect 7776 21786 7832 21788
rect 7856 21786 7912 21788
rect 7616 21734 7662 21786
rect 7662 21734 7672 21786
rect 7696 21734 7726 21786
rect 7726 21734 7738 21786
rect 7738 21734 7752 21786
rect 7776 21734 7790 21786
rect 7790 21734 7802 21786
rect 7802 21734 7832 21786
rect 7856 21734 7866 21786
rect 7866 21734 7912 21786
rect 7616 21732 7672 21734
rect 7696 21732 7752 21734
rect 7776 21732 7832 21734
rect 7856 21732 7912 21734
rect 7616 20698 7672 20700
rect 7696 20698 7752 20700
rect 7776 20698 7832 20700
rect 7856 20698 7912 20700
rect 7616 20646 7662 20698
rect 7662 20646 7672 20698
rect 7696 20646 7726 20698
rect 7726 20646 7738 20698
rect 7738 20646 7752 20698
rect 7776 20646 7790 20698
rect 7790 20646 7802 20698
rect 7802 20646 7832 20698
rect 7856 20646 7866 20698
rect 7866 20646 7912 20698
rect 7616 20644 7672 20646
rect 7696 20644 7752 20646
rect 7776 20644 7832 20646
rect 7856 20644 7912 20646
rect 7616 19610 7672 19612
rect 7696 19610 7752 19612
rect 7776 19610 7832 19612
rect 7856 19610 7912 19612
rect 7616 19558 7662 19610
rect 7662 19558 7672 19610
rect 7696 19558 7726 19610
rect 7726 19558 7738 19610
rect 7738 19558 7752 19610
rect 7776 19558 7790 19610
rect 7790 19558 7802 19610
rect 7802 19558 7832 19610
rect 7856 19558 7866 19610
rect 7866 19558 7912 19610
rect 7616 19556 7672 19558
rect 7696 19556 7752 19558
rect 7776 19556 7832 19558
rect 7856 19556 7912 19558
rect 7616 18522 7672 18524
rect 7696 18522 7752 18524
rect 7776 18522 7832 18524
rect 7856 18522 7912 18524
rect 7616 18470 7662 18522
rect 7662 18470 7672 18522
rect 7696 18470 7726 18522
rect 7726 18470 7738 18522
rect 7738 18470 7752 18522
rect 7776 18470 7790 18522
rect 7790 18470 7802 18522
rect 7802 18470 7832 18522
rect 7856 18470 7866 18522
rect 7866 18470 7912 18522
rect 7616 18468 7672 18470
rect 7696 18468 7752 18470
rect 7776 18468 7832 18470
rect 7856 18468 7912 18470
rect 7616 17434 7672 17436
rect 7696 17434 7752 17436
rect 7776 17434 7832 17436
rect 7856 17434 7912 17436
rect 7616 17382 7662 17434
rect 7662 17382 7672 17434
rect 7696 17382 7726 17434
rect 7726 17382 7738 17434
rect 7738 17382 7752 17434
rect 7776 17382 7790 17434
rect 7790 17382 7802 17434
rect 7802 17382 7832 17434
rect 7856 17382 7866 17434
rect 7866 17382 7912 17434
rect 7616 17380 7672 17382
rect 7696 17380 7752 17382
rect 7776 17380 7832 17382
rect 7856 17380 7912 17382
rect 6956 4922 7012 4924
rect 7036 4922 7092 4924
rect 7116 4922 7172 4924
rect 7196 4922 7252 4924
rect 6956 4870 7002 4922
rect 7002 4870 7012 4922
rect 7036 4870 7066 4922
rect 7066 4870 7078 4922
rect 7078 4870 7092 4922
rect 7116 4870 7130 4922
rect 7130 4870 7142 4922
rect 7142 4870 7172 4922
rect 7196 4870 7206 4922
rect 7206 4870 7252 4922
rect 6956 4868 7012 4870
rect 7036 4868 7092 4870
rect 7116 4868 7172 4870
rect 7196 4868 7252 4870
rect 7616 16346 7672 16348
rect 7696 16346 7752 16348
rect 7776 16346 7832 16348
rect 7856 16346 7912 16348
rect 7616 16294 7662 16346
rect 7662 16294 7672 16346
rect 7696 16294 7726 16346
rect 7726 16294 7738 16346
rect 7738 16294 7752 16346
rect 7776 16294 7790 16346
rect 7790 16294 7802 16346
rect 7802 16294 7832 16346
rect 7856 16294 7866 16346
rect 7866 16294 7912 16346
rect 7616 16292 7672 16294
rect 7696 16292 7752 16294
rect 7776 16292 7832 16294
rect 7856 16292 7912 16294
rect 7616 15258 7672 15260
rect 7696 15258 7752 15260
rect 7776 15258 7832 15260
rect 7856 15258 7912 15260
rect 7616 15206 7662 15258
rect 7662 15206 7672 15258
rect 7696 15206 7726 15258
rect 7726 15206 7738 15258
rect 7738 15206 7752 15258
rect 7776 15206 7790 15258
rect 7790 15206 7802 15258
rect 7802 15206 7832 15258
rect 7856 15206 7866 15258
rect 7866 15206 7912 15258
rect 7616 15204 7672 15206
rect 7696 15204 7752 15206
rect 7776 15204 7832 15206
rect 7856 15204 7912 15206
rect 7616 14170 7672 14172
rect 7696 14170 7752 14172
rect 7776 14170 7832 14172
rect 7856 14170 7912 14172
rect 7616 14118 7662 14170
rect 7662 14118 7672 14170
rect 7696 14118 7726 14170
rect 7726 14118 7738 14170
rect 7738 14118 7752 14170
rect 7776 14118 7790 14170
rect 7790 14118 7802 14170
rect 7802 14118 7832 14170
rect 7856 14118 7866 14170
rect 7866 14118 7912 14170
rect 7616 14116 7672 14118
rect 7696 14116 7752 14118
rect 7776 14116 7832 14118
rect 7856 14116 7912 14118
rect 7616 13082 7672 13084
rect 7696 13082 7752 13084
rect 7776 13082 7832 13084
rect 7856 13082 7912 13084
rect 7616 13030 7662 13082
rect 7662 13030 7672 13082
rect 7696 13030 7726 13082
rect 7726 13030 7738 13082
rect 7738 13030 7752 13082
rect 7776 13030 7790 13082
rect 7790 13030 7802 13082
rect 7802 13030 7832 13082
rect 7856 13030 7866 13082
rect 7866 13030 7912 13082
rect 7616 13028 7672 13030
rect 7696 13028 7752 13030
rect 7776 13028 7832 13030
rect 7856 13028 7912 13030
rect 7616 11994 7672 11996
rect 7696 11994 7752 11996
rect 7776 11994 7832 11996
rect 7856 11994 7912 11996
rect 7616 11942 7662 11994
rect 7662 11942 7672 11994
rect 7696 11942 7726 11994
rect 7726 11942 7738 11994
rect 7738 11942 7752 11994
rect 7776 11942 7790 11994
rect 7790 11942 7802 11994
rect 7802 11942 7832 11994
rect 7856 11942 7866 11994
rect 7866 11942 7912 11994
rect 7616 11940 7672 11942
rect 7696 11940 7752 11942
rect 7776 11940 7832 11942
rect 7856 11940 7912 11942
rect 7616 10906 7672 10908
rect 7696 10906 7752 10908
rect 7776 10906 7832 10908
rect 7856 10906 7912 10908
rect 7616 10854 7662 10906
rect 7662 10854 7672 10906
rect 7696 10854 7726 10906
rect 7726 10854 7738 10906
rect 7738 10854 7752 10906
rect 7776 10854 7790 10906
rect 7790 10854 7802 10906
rect 7802 10854 7832 10906
rect 7856 10854 7866 10906
rect 7866 10854 7912 10906
rect 7616 10852 7672 10854
rect 7696 10852 7752 10854
rect 7776 10852 7832 10854
rect 7856 10852 7912 10854
rect 7616 9818 7672 9820
rect 7696 9818 7752 9820
rect 7776 9818 7832 9820
rect 7856 9818 7912 9820
rect 7616 9766 7662 9818
rect 7662 9766 7672 9818
rect 7696 9766 7726 9818
rect 7726 9766 7738 9818
rect 7738 9766 7752 9818
rect 7776 9766 7790 9818
rect 7790 9766 7802 9818
rect 7802 9766 7832 9818
rect 7856 9766 7866 9818
rect 7866 9766 7912 9818
rect 7616 9764 7672 9766
rect 7696 9764 7752 9766
rect 7776 9764 7832 9766
rect 7856 9764 7912 9766
rect 7616 8730 7672 8732
rect 7696 8730 7752 8732
rect 7776 8730 7832 8732
rect 7856 8730 7912 8732
rect 7616 8678 7662 8730
rect 7662 8678 7672 8730
rect 7696 8678 7726 8730
rect 7726 8678 7738 8730
rect 7738 8678 7752 8730
rect 7776 8678 7790 8730
rect 7790 8678 7802 8730
rect 7802 8678 7832 8730
rect 7856 8678 7866 8730
rect 7866 8678 7912 8730
rect 7616 8676 7672 8678
rect 7696 8676 7752 8678
rect 7776 8676 7832 8678
rect 7856 8676 7912 8678
rect 7616 7642 7672 7644
rect 7696 7642 7752 7644
rect 7776 7642 7832 7644
rect 7856 7642 7912 7644
rect 7616 7590 7662 7642
rect 7662 7590 7672 7642
rect 7696 7590 7726 7642
rect 7726 7590 7738 7642
rect 7738 7590 7752 7642
rect 7776 7590 7790 7642
rect 7790 7590 7802 7642
rect 7802 7590 7832 7642
rect 7856 7590 7866 7642
rect 7866 7590 7912 7642
rect 7616 7588 7672 7590
rect 7696 7588 7752 7590
rect 7776 7588 7832 7590
rect 7856 7588 7912 7590
rect 7616 6554 7672 6556
rect 7696 6554 7752 6556
rect 7776 6554 7832 6556
rect 7856 6554 7912 6556
rect 7616 6502 7662 6554
rect 7662 6502 7672 6554
rect 7696 6502 7726 6554
rect 7726 6502 7738 6554
rect 7738 6502 7752 6554
rect 7776 6502 7790 6554
rect 7790 6502 7802 6554
rect 7802 6502 7832 6554
rect 7856 6502 7866 6554
rect 7866 6502 7912 6554
rect 7616 6500 7672 6502
rect 7696 6500 7752 6502
rect 7776 6500 7832 6502
rect 7856 6500 7912 6502
rect 7616 5466 7672 5468
rect 7696 5466 7752 5468
rect 7776 5466 7832 5468
rect 7856 5466 7912 5468
rect 7616 5414 7662 5466
rect 7662 5414 7672 5466
rect 7696 5414 7726 5466
rect 7726 5414 7738 5466
rect 7738 5414 7752 5466
rect 7776 5414 7790 5466
rect 7790 5414 7802 5466
rect 7802 5414 7832 5466
rect 7856 5414 7866 5466
rect 7866 5414 7912 5466
rect 7616 5412 7672 5414
rect 7696 5412 7752 5414
rect 7776 5412 7832 5414
rect 7856 5412 7912 5414
rect 7616 4378 7672 4380
rect 7696 4378 7752 4380
rect 7776 4378 7832 4380
rect 7856 4378 7912 4380
rect 7616 4326 7662 4378
rect 7662 4326 7672 4378
rect 7696 4326 7726 4378
rect 7726 4326 7738 4378
rect 7738 4326 7752 4378
rect 7776 4326 7790 4378
rect 7790 4326 7802 4378
rect 7802 4326 7832 4378
rect 7856 4326 7866 4378
rect 7866 4326 7912 4378
rect 7616 4324 7672 4326
rect 7696 4324 7752 4326
rect 7776 4324 7832 4326
rect 7856 4324 7912 4326
rect 6956 3834 7012 3836
rect 7036 3834 7092 3836
rect 7116 3834 7172 3836
rect 7196 3834 7252 3836
rect 6956 3782 7002 3834
rect 7002 3782 7012 3834
rect 7036 3782 7066 3834
rect 7066 3782 7078 3834
rect 7078 3782 7092 3834
rect 7116 3782 7130 3834
rect 7130 3782 7142 3834
rect 7142 3782 7172 3834
rect 7196 3782 7206 3834
rect 7206 3782 7252 3834
rect 6956 3780 7012 3782
rect 7036 3780 7092 3782
rect 7116 3780 7172 3782
rect 7196 3780 7252 3782
rect 2616 3290 2672 3292
rect 2696 3290 2752 3292
rect 2776 3290 2832 3292
rect 2856 3290 2912 3292
rect 2616 3238 2662 3290
rect 2662 3238 2672 3290
rect 2696 3238 2726 3290
rect 2726 3238 2738 3290
rect 2738 3238 2752 3290
rect 2776 3238 2790 3290
rect 2790 3238 2802 3290
rect 2802 3238 2832 3290
rect 2856 3238 2866 3290
rect 2866 3238 2912 3290
rect 2616 3236 2672 3238
rect 2696 3236 2752 3238
rect 2776 3236 2832 3238
rect 2856 3236 2912 3238
rect 7616 3290 7672 3292
rect 7696 3290 7752 3292
rect 7776 3290 7832 3292
rect 7856 3290 7912 3292
rect 7616 3238 7662 3290
rect 7662 3238 7672 3290
rect 7696 3238 7726 3290
rect 7726 3238 7738 3290
rect 7738 3238 7752 3290
rect 7776 3238 7790 3290
rect 7790 3238 7802 3290
rect 7802 3238 7832 3290
rect 7856 3238 7866 3290
rect 7866 3238 7912 3290
rect 7616 3236 7672 3238
rect 7696 3236 7752 3238
rect 7776 3236 7832 3238
rect 7856 3236 7912 3238
rect 9494 31184 9550 31240
rect 6956 2746 7012 2748
rect 7036 2746 7092 2748
rect 7116 2746 7172 2748
rect 7196 2746 7252 2748
rect 6956 2694 7002 2746
rect 7002 2694 7012 2746
rect 7036 2694 7066 2746
rect 7066 2694 7078 2746
rect 7078 2694 7092 2746
rect 7116 2694 7130 2746
rect 7130 2694 7142 2746
rect 7142 2694 7172 2746
rect 7196 2694 7206 2746
rect 7206 2694 7252 2746
rect 6956 2692 7012 2694
rect 7036 2692 7092 2694
rect 7116 2692 7172 2694
rect 7196 2692 7252 2694
rect 10782 56788 10784 56808
rect 10784 56788 10836 56808
rect 10836 56788 10838 56808
rect 10782 56752 10838 56788
rect 12616 68570 12672 68572
rect 12696 68570 12752 68572
rect 12776 68570 12832 68572
rect 12856 68570 12912 68572
rect 12616 68518 12662 68570
rect 12662 68518 12672 68570
rect 12696 68518 12726 68570
rect 12726 68518 12738 68570
rect 12738 68518 12752 68570
rect 12776 68518 12790 68570
rect 12790 68518 12802 68570
rect 12802 68518 12832 68570
rect 12856 68518 12866 68570
rect 12866 68518 12912 68570
rect 12616 68516 12672 68518
rect 12696 68516 12752 68518
rect 12776 68516 12832 68518
rect 12856 68516 12912 68518
rect 11956 68026 12012 68028
rect 12036 68026 12092 68028
rect 12116 68026 12172 68028
rect 12196 68026 12252 68028
rect 11956 67974 12002 68026
rect 12002 67974 12012 68026
rect 12036 67974 12066 68026
rect 12066 67974 12078 68026
rect 12078 67974 12092 68026
rect 12116 67974 12130 68026
rect 12130 67974 12142 68026
rect 12142 67974 12172 68026
rect 12196 67974 12206 68026
rect 12206 67974 12252 68026
rect 11956 67972 12012 67974
rect 12036 67972 12092 67974
rect 12116 67972 12172 67974
rect 12196 67972 12252 67974
rect 12616 67482 12672 67484
rect 12696 67482 12752 67484
rect 12776 67482 12832 67484
rect 12856 67482 12912 67484
rect 12616 67430 12662 67482
rect 12662 67430 12672 67482
rect 12696 67430 12726 67482
rect 12726 67430 12738 67482
rect 12738 67430 12752 67482
rect 12776 67430 12790 67482
rect 12790 67430 12802 67482
rect 12802 67430 12832 67482
rect 12856 67430 12866 67482
rect 12866 67430 12912 67482
rect 12616 67428 12672 67430
rect 12696 67428 12752 67430
rect 12776 67428 12832 67430
rect 12856 67428 12912 67430
rect 11956 66938 12012 66940
rect 12036 66938 12092 66940
rect 12116 66938 12172 66940
rect 12196 66938 12252 66940
rect 11956 66886 12002 66938
rect 12002 66886 12012 66938
rect 12036 66886 12066 66938
rect 12066 66886 12078 66938
rect 12078 66886 12092 66938
rect 12116 66886 12130 66938
rect 12130 66886 12142 66938
rect 12142 66886 12172 66938
rect 12196 66886 12206 66938
rect 12206 66886 12252 66938
rect 11956 66884 12012 66886
rect 12036 66884 12092 66886
rect 12116 66884 12172 66886
rect 12196 66884 12252 66886
rect 12616 66394 12672 66396
rect 12696 66394 12752 66396
rect 12776 66394 12832 66396
rect 12856 66394 12912 66396
rect 12616 66342 12662 66394
rect 12662 66342 12672 66394
rect 12696 66342 12726 66394
rect 12726 66342 12738 66394
rect 12738 66342 12752 66394
rect 12776 66342 12790 66394
rect 12790 66342 12802 66394
rect 12802 66342 12832 66394
rect 12856 66342 12866 66394
rect 12866 66342 12912 66394
rect 12616 66340 12672 66342
rect 12696 66340 12752 66342
rect 12776 66340 12832 66342
rect 12856 66340 12912 66342
rect 11956 65850 12012 65852
rect 12036 65850 12092 65852
rect 12116 65850 12172 65852
rect 12196 65850 12252 65852
rect 11956 65798 12002 65850
rect 12002 65798 12012 65850
rect 12036 65798 12066 65850
rect 12066 65798 12078 65850
rect 12078 65798 12092 65850
rect 12116 65798 12130 65850
rect 12130 65798 12142 65850
rect 12142 65798 12172 65850
rect 12196 65798 12206 65850
rect 12206 65798 12252 65850
rect 11956 65796 12012 65798
rect 12036 65796 12092 65798
rect 12116 65796 12172 65798
rect 12196 65796 12252 65798
rect 11956 64762 12012 64764
rect 12036 64762 12092 64764
rect 12116 64762 12172 64764
rect 12196 64762 12252 64764
rect 11956 64710 12002 64762
rect 12002 64710 12012 64762
rect 12036 64710 12066 64762
rect 12066 64710 12078 64762
rect 12078 64710 12092 64762
rect 12116 64710 12130 64762
rect 12130 64710 12142 64762
rect 12142 64710 12172 64762
rect 12196 64710 12206 64762
rect 12206 64710 12252 64762
rect 11956 64708 12012 64710
rect 12036 64708 12092 64710
rect 12116 64708 12172 64710
rect 12196 64708 12252 64710
rect 11956 63674 12012 63676
rect 12036 63674 12092 63676
rect 12116 63674 12172 63676
rect 12196 63674 12252 63676
rect 11956 63622 12002 63674
rect 12002 63622 12012 63674
rect 12036 63622 12066 63674
rect 12066 63622 12078 63674
rect 12078 63622 12092 63674
rect 12116 63622 12130 63674
rect 12130 63622 12142 63674
rect 12142 63622 12172 63674
rect 12196 63622 12206 63674
rect 12206 63622 12252 63674
rect 11956 63620 12012 63622
rect 12036 63620 12092 63622
rect 12116 63620 12172 63622
rect 12196 63620 12252 63622
rect 11956 62586 12012 62588
rect 12036 62586 12092 62588
rect 12116 62586 12172 62588
rect 12196 62586 12252 62588
rect 11956 62534 12002 62586
rect 12002 62534 12012 62586
rect 12036 62534 12066 62586
rect 12066 62534 12078 62586
rect 12078 62534 12092 62586
rect 12116 62534 12130 62586
rect 12130 62534 12142 62586
rect 12142 62534 12172 62586
rect 12196 62534 12206 62586
rect 12206 62534 12252 62586
rect 11956 62532 12012 62534
rect 12036 62532 12092 62534
rect 12116 62532 12172 62534
rect 12196 62532 12252 62534
rect 11956 61498 12012 61500
rect 12036 61498 12092 61500
rect 12116 61498 12172 61500
rect 12196 61498 12252 61500
rect 11956 61446 12002 61498
rect 12002 61446 12012 61498
rect 12036 61446 12066 61498
rect 12066 61446 12078 61498
rect 12078 61446 12092 61498
rect 12116 61446 12130 61498
rect 12130 61446 12142 61498
rect 12142 61446 12172 61498
rect 12196 61446 12206 61498
rect 12206 61446 12252 61498
rect 11956 61444 12012 61446
rect 12036 61444 12092 61446
rect 12116 61444 12172 61446
rect 12196 61444 12252 61446
rect 11956 60410 12012 60412
rect 12036 60410 12092 60412
rect 12116 60410 12172 60412
rect 12196 60410 12252 60412
rect 11956 60358 12002 60410
rect 12002 60358 12012 60410
rect 12036 60358 12066 60410
rect 12066 60358 12078 60410
rect 12078 60358 12092 60410
rect 12116 60358 12130 60410
rect 12130 60358 12142 60410
rect 12142 60358 12172 60410
rect 12196 60358 12206 60410
rect 12206 60358 12252 60410
rect 11956 60356 12012 60358
rect 12036 60356 12092 60358
rect 12116 60356 12172 60358
rect 12196 60356 12252 60358
rect 11956 59322 12012 59324
rect 12036 59322 12092 59324
rect 12116 59322 12172 59324
rect 12196 59322 12252 59324
rect 11956 59270 12002 59322
rect 12002 59270 12012 59322
rect 12036 59270 12066 59322
rect 12066 59270 12078 59322
rect 12078 59270 12092 59322
rect 12116 59270 12130 59322
rect 12130 59270 12142 59322
rect 12142 59270 12172 59322
rect 12196 59270 12206 59322
rect 12206 59270 12252 59322
rect 11956 59268 12012 59270
rect 12036 59268 12092 59270
rect 12116 59268 12172 59270
rect 12196 59268 12252 59270
rect 11956 58234 12012 58236
rect 12036 58234 12092 58236
rect 12116 58234 12172 58236
rect 12196 58234 12252 58236
rect 11956 58182 12002 58234
rect 12002 58182 12012 58234
rect 12036 58182 12066 58234
rect 12066 58182 12078 58234
rect 12078 58182 12092 58234
rect 12116 58182 12130 58234
rect 12130 58182 12142 58234
rect 12142 58182 12172 58234
rect 12196 58182 12206 58234
rect 12206 58182 12252 58234
rect 11956 58180 12012 58182
rect 12036 58180 12092 58182
rect 12116 58180 12172 58182
rect 12196 58180 12252 58182
rect 11956 57146 12012 57148
rect 12036 57146 12092 57148
rect 12116 57146 12172 57148
rect 12196 57146 12252 57148
rect 11956 57094 12002 57146
rect 12002 57094 12012 57146
rect 12036 57094 12066 57146
rect 12066 57094 12078 57146
rect 12078 57094 12092 57146
rect 12116 57094 12130 57146
rect 12130 57094 12142 57146
rect 12142 57094 12172 57146
rect 12196 57094 12206 57146
rect 12206 57094 12252 57146
rect 11956 57092 12012 57094
rect 12036 57092 12092 57094
rect 12116 57092 12172 57094
rect 12196 57092 12252 57094
rect 11956 56058 12012 56060
rect 12036 56058 12092 56060
rect 12116 56058 12172 56060
rect 12196 56058 12252 56060
rect 11956 56006 12002 56058
rect 12002 56006 12012 56058
rect 12036 56006 12066 56058
rect 12066 56006 12078 56058
rect 12078 56006 12092 56058
rect 12116 56006 12130 56058
rect 12130 56006 12142 56058
rect 12142 56006 12172 56058
rect 12196 56006 12206 56058
rect 12206 56006 12252 56058
rect 11956 56004 12012 56006
rect 12036 56004 12092 56006
rect 12116 56004 12172 56006
rect 12196 56004 12252 56006
rect 11956 54970 12012 54972
rect 12036 54970 12092 54972
rect 12116 54970 12172 54972
rect 12196 54970 12252 54972
rect 11956 54918 12002 54970
rect 12002 54918 12012 54970
rect 12036 54918 12066 54970
rect 12066 54918 12078 54970
rect 12078 54918 12092 54970
rect 12116 54918 12130 54970
rect 12130 54918 12142 54970
rect 12142 54918 12172 54970
rect 12196 54918 12206 54970
rect 12206 54918 12252 54970
rect 11956 54916 12012 54918
rect 12036 54916 12092 54918
rect 12116 54916 12172 54918
rect 12196 54916 12252 54918
rect 11956 53882 12012 53884
rect 12036 53882 12092 53884
rect 12116 53882 12172 53884
rect 12196 53882 12252 53884
rect 11956 53830 12002 53882
rect 12002 53830 12012 53882
rect 12036 53830 12066 53882
rect 12066 53830 12078 53882
rect 12078 53830 12092 53882
rect 12116 53830 12130 53882
rect 12130 53830 12142 53882
rect 12142 53830 12172 53882
rect 12196 53830 12206 53882
rect 12206 53830 12252 53882
rect 11956 53828 12012 53830
rect 12036 53828 12092 53830
rect 12116 53828 12172 53830
rect 12196 53828 12252 53830
rect 11956 52794 12012 52796
rect 12036 52794 12092 52796
rect 12116 52794 12172 52796
rect 12196 52794 12252 52796
rect 11956 52742 12002 52794
rect 12002 52742 12012 52794
rect 12036 52742 12066 52794
rect 12066 52742 12078 52794
rect 12078 52742 12092 52794
rect 12116 52742 12130 52794
rect 12130 52742 12142 52794
rect 12142 52742 12172 52794
rect 12196 52742 12206 52794
rect 12206 52742 12252 52794
rect 11956 52740 12012 52742
rect 12036 52740 12092 52742
rect 12116 52740 12172 52742
rect 12196 52740 12252 52742
rect 11956 51706 12012 51708
rect 12036 51706 12092 51708
rect 12116 51706 12172 51708
rect 12196 51706 12252 51708
rect 11956 51654 12002 51706
rect 12002 51654 12012 51706
rect 12036 51654 12066 51706
rect 12066 51654 12078 51706
rect 12078 51654 12092 51706
rect 12116 51654 12130 51706
rect 12130 51654 12142 51706
rect 12142 51654 12172 51706
rect 12196 51654 12206 51706
rect 12206 51654 12252 51706
rect 11956 51652 12012 51654
rect 12036 51652 12092 51654
rect 12116 51652 12172 51654
rect 12196 51652 12252 51654
rect 11956 50618 12012 50620
rect 12036 50618 12092 50620
rect 12116 50618 12172 50620
rect 12196 50618 12252 50620
rect 11956 50566 12002 50618
rect 12002 50566 12012 50618
rect 12036 50566 12066 50618
rect 12066 50566 12078 50618
rect 12078 50566 12092 50618
rect 12116 50566 12130 50618
rect 12130 50566 12142 50618
rect 12142 50566 12172 50618
rect 12196 50566 12206 50618
rect 12206 50566 12252 50618
rect 11956 50564 12012 50566
rect 12036 50564 12092 50566
rect 12116 50564 12172 50566
rect 12196 50564 12252 50566
rect 11956 49530 12012 49532
rect 12036 49530 12092 49532
rect 12116 49530 12172 49532
rect 12196 49530 12252 49532
rect 11956 49478 12002 49530
rect 12002 49478 12012 49530
rect 12036 49478 12066 49530
rect 12066 49478 12078 49530
rect 12078 49478 12092 49530
rect 12116 49478 12130 49530
rect 12130 49478 12142 49530
rect 12142 49478 12172 49530
rect 12196 49478 12206 49530
rect 12206 49478 12252 49530
rect 11956 49476 12012 49478
rect 12036 49476 12092 49478
rect 12116 49476 12172 49478
rect 12196 49476 12252 49478
rect 11956 48442 12012 48444
rect 12036 48442 12092 48444
rect 12116 48442 12172 48444
rect 12196 48442 12252 48444
rect 11956 48390 12002 48442
rect 12002 48390 12012 48442
rect 12036 48390 12066 48442
rect 12066 48390 12078 48442
rect 12078 48390 12092 48442
rect 12116 48390 12130 48442
rect 12130 48390 12142 48442
rect 12142 48390 12172 48442
rect 12196 48390 12206 48442
rect 12206 48390 12252 48442
rect 11956 48388 12012 48390
rect 12036 48388 12092 48390
rect 12116 48388 12172 48390
rect 12196 48388 12252 48390
rect 11956 47354 12012 47356
rect 12036 47354 12092 47356
rect 12116 47354 12172 47356
rect 12196 47354 12252 47356
rect 11956 47302 12002 47354
rect 12002 47302 12012 47354
rect 12036 47302 12066 47354
rect 12066 47302 12078 47354
rect 12078 47302 12092 47354
rect 12116 47302 12130 47354
rect 12130 47302 12142 47354
rect 12142 47302 12172 47354
rect 12196 47302 12206 47354
rect 12206 47302 12252 47354
rect 11956 47300 12012 47302
rect 12036 47300 12092 47302
rect 12116 47300 12172 47302
rect 12196 47300 12252 47302
rect 11956 46266 12012 46268
rect 12036 46266 12092 46268
rect 12116 46266 12172 46268
rect 12196 46266 12252 46268
rect 11956 46214 12002 46266
rect 12002 46214 12012 46266
rect 12036 46214 12066 46266
rect 12066 46214 12078 46266
rect 12078 46214 12092 46266
rect 12116 46214 12130 46266
rect 12130 46214 12142 46266
rect 12142 46214 12172 46266
rect 12196 46214 12206 46266
rect 12206 46214 12252 46266
rect 11956 46212 12012 46214
rect 12036 46212 12092 46214
rect 12116 46212 12172 46214
rect 12196 46212 12252 46214
rect 11956 45178 12012 45180
rect 12036 45178 12092 45180
rect 12116 45178 12172 45180
rect 12196 45178 12252 45180
rect 11956 45126 12002 45178
rect 12002 45126 12012 45178
rect 12036 45126 12066 45178
rect 12066 45126 12078 45178
rect 12078 45126 12092 45178
rect 12116 45126 12130 45178
rect 12130 45126 12142 45178
rect 12142 45126 12172 45178
rect 12196 45126 12206 45178
rect 12206 45126 12252 45178
rect 11956 45124 12012 45126
rect 12036 45124 12092 45126
rect 12116 45124 12172 45126
rect 12196 45124 12252 45126
rect 12616 65306 12672 65308
rect 12696 65306 12752 65308
rect 12776 65306 12832 65308
rect 12856 65306 12912 65308
rect 12616 65254 12662 65306
rect 12662 65254 12672 65306
rect 12696 65254 12726 65306
rect 12726 65254 12738 65306
rect 12738 65254 12752 65306
rect 12776 65254 12790 65306
rect 12790 65254 12802 65306
rect 12802 65254 12832 65306
rect 12856 65254 12866 65306
rect 12866 65254 12912 65306
rect 12616 65252 12672 65254
rect 12696 65252 12752 65254
rect 12776 65252 12832 65254
rect 12856 65252 12912 65254
rect 12616 64218 12672 64220
rect 12696 64218 12752 64220
rect 12776 64218 12832 64220
rect 12856 64218 12912 64220
rect 12616 64166 12662 64218
rect 12662 64166 12672 64218
rect 12696 64166 12726 64218
rect 12726 64166 12738 64218
rect 12738 64166 12752 64218
rect 12776 64166 12790 64218
rect 12790 64166 12802 64218
rect 12802 64166 12832 64218
rect 12856 64166 12866 64218
rect 12866 64166 12912 64218
rect 12616 64164 12672 64166
rect 12696 64164 12752 64166
rect 12776 64164 12832 64166
rect 12856 64164 12912 64166
rect 12616 63130 12672 63132
rect 12696 63130 12752 63132
rect 12776 63130 12832 63132
rect 12856 63130 12912 63132
rect 12616 63078 12662 63130
rect 12662 63078 12672 63130
rect 12696 63078 12726 63130
rect 12726 63078 12738 63130
rect 12738 63078 12752 63130
rect 12776 63078 12790 63130
rect 12790 63078 12802 63130
rect 12802 63078 12832 63130
rect 12856 63078 12866 63130
rect 12866 63078 12912 63130
rect 12616 63076 12672 63078
rect 12696 63076 12752 63078
rect 12776 63076 12832 63078
rect 12856 63076 12912 63078
rect 12616 62042 12672 62044
rect 12696 62042 12752 62044
rect 12776 62042 12832 62044
rect 12856 62042 12912 62044
rect 12616 61990 12662 62042
rect 12662 61990 12672 62042
rect 12696 61990 12726 62042
rect 12726 61990 12738 62042
rect 12738 61990 12752 62042
rect 12776 61990 12790 62042
rect 12790 61990 12802 62042
rect 12802 61990 12832 62042
rect 12856 61990 12866 62042
rect 12866 61990 12912 62042
rect 12616 61988 12672 61990
rect 12696 61988 12752 61990
rect 12776 61988 12832 61990
rect 12856 61988 12912 61990
rect 12616 60954 12672 60956
rect 12696 60954 12752 60956
rect 12776 60954 12832 60956
rect 12856 60954 12912 60956
rect 12616 60902 12662 60954
rect 12662 60902 12672 60954
rect 12696 60902 12726 60954
rect 12726 60902 12738 60954
rect 12738 60902 12752 60954
rect 12776 60902 12790 60954
rect 12790 60902 12802 60954
rect 12802 60902 12832 60954
rect 12856 60902 12866 60954
rect 12866 60902 12912 60954
rect 12616 60900 12672 60902
rect 12696 60900 12752 60902
rect 12776 60900 12832 60902
rect 12856 60900 12912 60902
rect 12616 59866 12672 59868
rect 12696 59866 12752 59868
rect 12776 59866 12832 59868
rect 12856 59866 12912 59868
rect 12616 59814 12662 59866
rect 12662 59814 12672 59866
rect 12696 59814 12726 59866
rect 12726 59814 12738 59866
rect 12738 59814 12752 59866
rect 12776 59814 12790 59866
rect 12790 59814 12802 59866
rect 12802 59814 12832 59866
rect 12856 59814 12866 59866
rect 12866 59814 12912 59866
rect 12616 59812 12672 59814
rect 12696 59812 12752 59814
rect 12776 59812 12832 59814
rect 12856 59812 12912 59814
rect 12616 58778 12672 58780
rect 12696 58778 12752 58780
rect 12776 58778 12832 58780
rect 12856 58778 12912 58780
rect 12616 58726 12662 58778
rect 12662 58726 12672 58778
rect 12696 58726 12726 58778
rect 12726 58726 12738 58778
rect 12738 58726 12752 58778
rect 12776 58726 12790 58778
rect 12790 58726 12802 58778
rect 12802 58726 12832 58778
rect 12856 58726 12866 58778
rect 12866 58726 12912 58778
rect 12616 58724 12672 58726
rect 12696 58724 12752 58726
rect 12776 58724 12832 58726
rect 12856 58724 12912 58726
rect 12616 57690 12672 57692
rect 12696 57690 12752 57692
rect 12776 57690 12832 57692
rect 12856 57690 12912 57692
rect 12616 57638 12662 57690
rect 12662 57638 12672 57690
rect 12696 57638 12726 57690
rect 12726 57638 12738 57690
rect 12738 57638 12752 57690
rect 12776 57638 12790 57690
rect 12790 57638 12802 57690
rect 12802 57638 12832 57690
rect 12856 57638 12866 57690
rect 12866 57638 12912 57690
rect 12616 57636 12672 57638
rect 12696 57636 12752 57638
rect 12776 57636 12832 57638
rect 12856 57636 12912 57638
rect 12616 56602 12672 56604
rect 12696 56602 12752 56604
rect 12776 56602 12832 56604
rect 12856 56602 12912 56604
rect 12616 56550 12662 56602
rect 12662 56550 12672 56602
rect 12696 56550 12726 56602
rect 12726 56550 12738 56602
rect 12738 56550 12752 56602
rect 12776 56550 12790 56602
rect 12790 56550 12802 56602
rect 12802 56550 12832 56602
rect 12856 56550 12866 56602
rect 12866 56550 12912 56602
rect 12616 56548 12672 56550
rect 12696 56548 12752 56550
rect 12776 56548 12832 56550
rect 12856 56548 12912 56550
rect 12616 55514 12672 55516
rect 12696 55514 12752 55516
rect 12776 55514 12832 55516
rect 12856 55514 12912 55516
rect 12616 55462 12662 55514
rect 12662 55462 12672 55514
rect 12696 55462 12726 55514
rect 12726 55462 12738 55514
rect 12738 55462 12752 55514
rect 12776 55462 12790 55514
rect 12790 55462 12802 55514
rect 12802 55462 12832 55514
rect 12856 55462 12866 55514
rect 12866 55462 12912 55514
rect 12616 55460 12672 55462
rect 12696 55460 12752 55462
rect 12776 55460 12832 55462
rect 12856 55460 12912 55462
rect 12616 54426 12672 54428
rect 12696 54426 12752 54428
rect 12776 54426 12832 54428
rect 12856 54426 12912 54428
rect 12616 54374 12662 54426
rect 12662 54374 12672 54426
rect 12696 54374 12726 54426
rect 12726 54374 12738 54426
rect 12738 54374 12752 54426
rect 12776 54374 12790 54426
rect 12790 54374 12802 54426
rect 12802 54374 12832 54426
rect 12856 54374 12866 54426
rect 12866 54374 12912 54426
rect 12616 54372 12672 54374
rect 12696 54372 12752 54374
rect 12776 54372 12832 54374
rect 12856 54372 12912 54374
rect 12616 53338 12672 53340
rect 12696 53338 12752 53340
rect 12776 53338 12832 53340
rect 12856 53338 12912 53340
rect 12616 53286 12662 53338
rect 12662 53286 12672 53338
rect 12696 53286 12726 53338
rect 12726 53286 12738 53338
rect 12738 53286 12752 53338
rect 12776 53286 12790 53338
rect 12790 53286 12802 53338
rect 12802 53286 12832 53338
rect 12856 53286 12866 53338
rect 12866 53286 12912 53338
rect 12616 53284 12672 53286
rect 12696 53284 12752 53286
rect 12776 53284 12832 53286
rect 12856 53284 12912 53286
rect 12616 52250 12672 52252
rect 12696 52250 12752 52252
rect 12776 52250 12832 52252
rect 12856 52250 12912 52252
rect 12616 52198 12662 52250
rect 12662 52198 12672 52250
rect 12696 52198 12726 52250
rect 12726 52198 12738 52250
rect 12738 52198 12752 52250
rect 12776 52198 12790 52250
rect 12790 52198 12802 52250
rect 12802 52198 12832 52250
rect 12856 52198 12866 52250
rect 12866 52198 12912 52250
rect 12616 52196 12672 52198
rect 12696 52196 12752 52198
rect 12776 52196 12832 52198
rect 12856 52196 12912 52198
rect 12616 51162 12672 51164
rect 12696 51162 12752 51164
rect 12776 51162 12832 51164
rect 12856 51162 12912 51164
rect 12616 51110 12662 51162
rect 12662 51110 12672 51162
rect 12696 51110 12726 51162
rect 12726 51110 12738 51162
rect 12738 51110 12752 51162
rect 12776 51110 12790 51162
rect 12790 51110 12802 51162
rect 12802 51110 12832 51162
rect 12856 51110 12866 51162
rect 12866 51110 12912 51162
rect 12616 51108 12672 51110
rect 12696 51108 12752 51110
rect 12776 51108 12832 51110
rect 12856 51108 12912 51110
rect 12616 50074 12672 50076
rect 12696 50074 12752 50076
rect 12776 50074 12832 50076
rect 12856 50074 12912 50076
rect 12616 50022 12662 50074
rect 12662 50022 12672 50074
rect 12696 50022 12726 50074
rect 12726 50022 12738 50074
rect 12738 50022 12752 50074
rect 12776 50022 12790 50074
rect 12790 50022 12802 50074
rect 12802 50022 12832 50074
rect 12856 50022 12866 50074
rect 12866 50022 12912 50074
rect 12616 50020 12672 50022
rect 12696 50020 12752 50022
rect 12776 50020 12832 50022
rect 12856 50020 12912 50022
rect 12616 48986 12672 48988
rect 12696 48986 12752 48988
rect 12776 48986 12832 48988
rect 12856 48986 12912 48988
rect 12616 48934 12662 48986
rect 12662 48934 12672 48986
rect 12696 48934 12726 48986
rect 12726 48934 12738 48986
rect 12738 48934 12752 48986
rect 12776 48934 12790 48986
rect 12790 48934 12802 48986
rect 12802 48934 12832 48986
rect 12856 48934 12866 48986
rect 12866 48934 12912 48986
rect 12616 48932 12672 48934
rect 12696 48932 12752 48934
rect 12776 48932 12832 48934
rect 12856 48932 12912 48934
rect 12616 47898 12672 47900
rect 12696 47898 12752 47900
rect 12776 47898 12832 47900
rect 12856 47898 12912 47900
rect 12616 47846 12662 47898
rect 12662 47846 12672 47898
rect 12696 47846 12726 47898
rect 12726 47846 12738 47898
rect 12738 47846 12752 47898
rect 12776 47846 12790 47898
rect 12790 47846 12802 47898
rect 12802 47846 12832 47898
rect 12856 47846 12866 47898
rect 12866 47846 12912 47898
rect 12616 47844 12672 47846
rect 12696 47844 12752 47846
rect 12776 47844 12832 47846
rect 12856 47844 12912 47846
rect 12616 46810 12672 46812
rect 12696 46810 12752 46812
rect 12776 46810 12832 46812
rect 12856 46810 12912 46812
rect 12616 46758 12662 46810
rect 12662 46758 12672 46810
rect 12696 46758 12726 46810
rect 12726 46758 12738 46810
rect 12738 46758 12752 46810
rect 12776 46758 12790 46810
rect 12790 46758 12802 46810
rect 12802 46758 12832 46810
rect 12856 46758 12866 46810
rect 12866 46758 12912 46810
rect 12616 46756 12672 46758
rect 12696 46756 12752 46758
rect 12776 46756 12832 46758
rect 12856 46756 12912 46758
rect 12616 45722 12672 45724
rect 12696 45722 12752 45724
rect 12776 45722 12832 45724
rect 12856 45722 12912 45724
rect 12616 45670 12662 45722
rect 12662 45670 12672 45722
rect 12696 45670 12726 45722
rect 12726 45670 12738 45722
rect 12738 45670 12752 45722
rect 12776 45670 12790 45722
rect 12790 45670 12802 45722
rect 12802 45670 12832 45722
rect 12856 45670 12866 45722
rect 12866 45670 12912 45722
rect 12616 45668 12672 45670
rect 12696 45668 12752 45670
rect 12776 45668 12832 45670
rect 12856 45668 12912 45670
rect 12616 44634 12672 44636
rect 12696 44634 12752 44636
rect 12776 44634 12832 44636
rect 12856 44634 12912 44636
rect 12616 44582 12662 44634
rect 12662 44582 12672 44634
rect 12696 44582 12726 44634
rect 12726 44582 12738 44634
rect 12738 44582 12752 44634
rect 12776 44582 12790 44634
rect 12790 44582 12802 44634
rect 12802 44582 12832 44634
rect 12856 44582 12866 44634
rect 12866 44582 12912 44634
rect 12616 44580 12672 44582
rect 12696 44580 12752 44582
rect 12776 44580 12832 44582
rect 12856 44580 12912 44582
rect 11956 44090 12012 44092
rect 12036 44090 12092 44092
rect 12116 44090 12172 44092
rect 12196 44090 12252 44092
rect 11956 44038 12002 44090
rect 12002 44038 12012 44090
rect 12036 44038 12066 44090
rect 12066 44038 12078 44090
rect 12078 44038 12092 44090
rect 12116 44038 12130 44090
rect 12130 44038 12142 44090
rect 12142 44038 12172 44090
rect 12196 44038 12206 44090
rect 12206 44038 12252 44090
rect 11956 44036 12012 44038
rect 12036 44036 12092 44038
rect 12116 44036 12172 44038
rect 12196 44036 12252 44038
rect 12616 43546 12672 43548
rect 12696 43546 12752 43548
rect 12776 43546 12832 43548
rect 12856 43546 12912 43548
rect 12616 43494 12662 43546
rect 12662 43494 12672 43546
rect 12696 43494 12726 43546
rect 12726 43494 12738 43546
rect 12738 43494 12752 43546
rect 12776 43494 12790 43546
rect 12790 43494 12802 43546
rect 12802 43494 12832 43546
rect 12856 43494 12866 43546
rect 12866 43494 12912 43546
rect 12616 43492 12672 43494
rect 12696 43492 12752 43494
rect 12776 43492 12832 43494
rect 12856 43492 12912 43494
rect 11956 43002 12012 43004
rect 12036 43002 12092 43004
rect 12116 43002 12172 43004
rect 12196 43002 12252 43004
rect 11956 42950 12002 43002
rect 12002 42950 12012 43002
rect 12036 42950 12066 43002
rect 12066 42950 12078 43002
rect 12078 42950 12092 43002
rect 12116 42950 12130 43002
rect 12130 42950 12142 43002
rect 12142 42950 12172 43002
rect 12196 42950 12206 43002
rect 12206 42950 12252 43002
rect 11956 42948 12012 42950
rect 12036 42948 12092 42950
rect 12116 42948 12172 42950
rect 12196 42948 12252 42950
rect 11956 41914 12012 41916
rect 12036 41914 12092 41916
rect 12116 41914 12172 41916
rect 12196 41914 12252 41916
rect 11956 41862 12002 41914
rect 12002 41862 12012 41914
rect 12036 41862 12066 41914
rect 12066 41862 12078 41914
rect 12078 41862 12092 41914
rect 12116 41862 12130 41914
rect 12130 41862 12142 41914
rect 12142 41862 12172 41914
rect 12196 41862 12206 41914
rect 12206 41862 12252 41914
rect 11956 41860 12012 41862
rect 12036 41860 12092 41862
rect 12116 41860 12172 41862
rect 12196 41860 12252 41862
rect 11956 40826 12012 40828
rect 12036 40826 12092 40828
rect 12116 40826 12172 40828
rect 12196 40826 12252 40828
rect 11956 40774 12002 40826
rect 12002 40774 12012 40826
rect 12036 40774 12066 40826
rect 12066 40774 12078 40826
rect 12078 40774 12092 40826
rect 12116 40774 12130 40826
rect 12130 40774 12142 40826
rect 12142 40774 12172 40826
rect 12196 40774 12206 40826
rect 12206 40774 12252 40826
rect 11956 40772 12012 40774
rect 12036 40772 12092 40774
rect 12116 40772 12172 40774
rect 12196 40772 12252 40774
rect 11956 39738 12012 39740
rect 12036 39738 12092 39740
rect 12116 39738 12172 39740
rect 12196 39738 12252 39740
rect 11956 39686 12002 39738
rect 12002 39686 12012 39738
rect 12036 39686 12066 39738
rect 12066 39686 12078 39738
rect 12078 39686 12092 39738
rect 12116 39686 12130 39738
rect 12130 39686 12142 39738
rect 12142 39686 12172 39738
rect 12196 39686 12206 39738
rect 12206 39686 12252 39738
rect 11956 39684 12012 39686
rect 12036 39684 12092 39686
rect 12116 39684 12172 39686
rect 12196 39684 12252 39686
rect 11956 38650 12012 38652
rect 12036 38650 12092 38652
rect 12116 38650 12172 38652
rect 12196 38650 12252 38652
rect 11956 38598 12002 38650
rect 12002 38598 12012 38650
rect 12036 38598 12066 38650
rect 12066 38598 12078 38650
rect 12078 38598 12092 38650
rect 12116 38598 12130 38650
rect 12130 38598 12142 38650
rect 12142 38598 12172 38650
rect 12196 38598 12206 38650
rect 12206 38598 12252 38650
rect 11956 38596 12012 38598
rect 12036 38596 12092 38598
rect 12116 38596 12172 38598
rect 12196 38596 12252 38598
rect 11956 37562 12012 37564
rect 12036 37562 12092 37564
rect 12116 37562 12172 37564
rect 12196 37562 12252 37564
rect 11956 37510 12002 37562
rect 12002 37510 12012 37562
rect 12036 37510 12066 37562
rect 12066 37510 12078 37562
rect 12078 37510 12092 37562
rect 12116 37510 12130 37562
rect 12130 37510 12142 37562
rect 12142 37510 12172 37562
rect 12196 37510 12206 37562
rect 12206 37510 12252 37562
rect 11956 37508 12012 37510
rect 12036 37508 12092 37510
rect 12116 37508 12172 37510
rect 12196 37508 12252 37510
rect 11956 36474 12012 36476
rect 12036 36474 12092 36476
rect 12116 36474 12172 36476
rect 12196 36474 12252 36476
rect 11956 36422 12002 36474
rect 12002 36422 12012 36474
rect 12036 36422 12066 36474
rect 12066 36422 12078 36474
rect 12078 36422 12092 36474
rect 12116 36422 12130 36474
rect 12130 36422 12142 36474
rect 12142 36422 12172 36474
rect 12196 36422 12206 36474
rect 12206 36422 12252 36474
rect 11956 36420 12012 36422
rect 12036 36420 12092 36422
rect 12116 36420 12172 36422
rect 12196 36420 12252 36422
rect 11956 35386 12012 35388
rect 12036 35386 12092 35388
rect 12116 35386 12172 35388
rect 12196 35386 12252 35388
rect 11956 35334 12002 35386
rect 12002 35334 12012 35386
rect 12036 35334 12066 35386
rect 12066 35334 12078 35386
rect 12078 35334 12092 35386
rect 12116 35334 12130 35386
rect 12130 35334 12142 35386
rect 12142 35334 12172 35386
rect 12196 35334 12206 35386
rect 12206 35334 12252 35386
rect 11956 35332 12012 35334
rect 12036 35332 12092 35334
rect 12116 35332 12172 35334
rect 12196 35332 12252 35334
rect 11956 34298 12012 34300
rect 12036 34298 12092 34300
rect 12116 34298 12172 34300
rect 12196 34298 12252 34300
rect 11956 34246 12002 34298
rect 12002 34246 12012 34298
rect 12036 34246 12066 34298
rect 12066 34246 12078 34298
rect 12078 34246 12092 34298
rect 12116 34246 12130 34298
rect 12130 34246 12142 34298
rect 12142 34246 12172 34298
rect 12196 34246 12206 34298
rect 12206 34246 12252 34298
rect 11956 34244 12012 34246
rect 12036 34244 12092 34246
rect 12116 34244 12172 34246
rect 12196 34244 12252 34246
rect 11956 33210 12012 33212
rect 12036 33210 12092 33212
rect 12116 33210 12172 33212
rect 12196 33210 12252 33212
rect 11956 33158 12002 33210
rect 12002 33158 12012 33210
rect 12036 33158 12066 33210
rect 12066 33158 12078 33210
rect 12078 33158 12092 33210
rect 12116 33158 12130 33210
rect 12130 33158 12142 33210
rect 12142 33158 12172 33210
rect 12196 33158 12206 33210
rect 12206 33158 12252 33210
rect 11956 33156 12012 33158
rect 12036 33156 12092 33158
rect 12116 33156 12172 33158
rect 12196 33156 12252 33158
rect 11956 32122 12012 32124
rect 12036 32122 12092 32124
rect 12116 32122 12172 32124
rect 12196 32122 12252 32124
rect 11956 32070 12002 32122
rect 12002 32070 12012 32122
rect 12036 32070 12066 32122
rect 12066 32070 12078 32122
rect 12078 32070 12092 32122
rect 12116 32070 12130 32122
rect 12130 32070 12142 32122
rect 12142 32070 12172 32122
rect 12196 32070 12206 32122
rect 12206 32070 12252 32122
rect 11956 32068 12012 32070
rect 12036 32068 12092 32070
rect 12116 32068 12172 32070
rect 12196 32068 12252 32070
rect 11956 31034 12012 31036
rect 12036 31034 12092 31036
rect 12116 31034 12172 31036
rect 12196 31034 12252 31036
rect 11956 30982 12002 31034
rect 12002 30982 12012 31034
rect 12036 30982 12066 31034
rect 12066 30982 12078 31034
rect 12078 30982 12092 31034
rect 12116 30982 12130 31034
rect 12130 30982 12142 31034
rect 12142 30982 12172 31034
rect 12196 30982 12206 31034
rect 12206 30982 12252 31034
rect 11956 30980 12012 30982
rect 12036 30980 12092 30982
rect 12116 30980 12172 30982
rect 12196 30980 12252 30982
rect 11956 29946 12012 29948
rect 12036 29946 12092 29948
rect 12116 29946 12172 29948
rect 12196 29946 12252 29948
rect 11956 29894 12002 29946
rect 12002 29894 12012 29946
rect 12036 29894 12066 29946
rect 12066 29894 12078 29946
rect 12078 29894 12092 29946
rect 12116 29894 12130 29946
rect 12130 29894 12142 29946
rect 12142 29894 12172 29946
rect 12196 29894 12206 29946
rect 12206 29894 12252 29946
rect 11956 29892 12012 29894
rect 12036 29892 12092 29894
rect 12116 29892 12172 29894
rect 12196 29892 12252 29894
rect 11956 28858 12012 28860
rect 12036 28858 12092 28860
rect 12116 28858 12172 28860
rect 12196 28858 12252 28860
rect 11956 28806 12002 28858
rect 12002 28806 12012 28858
rect 12036 28806 12066 28858
rect 12066 28806 12078 28858
rect 12078 28806 12092 28858
rect 12116 28806 12130 28858
rect 12130 28806 12142 28858
rect 12142 28806 12172 28858
rect 12196 28806 12206 28858
rect 12206 28806 12252 28858
rect 11956 28804 12012 28806
rect 12036 28804 12092 28806
rect 12116 28804 12172 28806
rect 12196 28804 12252 28806
rect 11956 27770 12012 27772
rect 12036 27770 12092 27772
rect 12116 27770 12172 27772
rect 12196 27770 12252 27772
rect 11956 27718 12002 27770
rect 12002 27718 12012 27770
rect 12036 27718 12066 27770
rect 12066 27718 12078 27770
rect 12078 27718 12092 27770
rect 12116 27718 12130 27770
rect 12130 27718 12142 27770
rect 12142 27718 12172 27770
rect 12196 27718 12206 27770
rect 12206 27718 12252 27770
rect 11956 27716 12012 27718
rect 12036 27716 12092 27718
rect 12116 27716 12172 27718
rect 12196 27716 12252 27718
rect 11956 26682 12012 26684
rect 12036 26682 12092 26684
rect 12116 26682 12172 26684
rect 12196 26682 12252 26684
rect 11956 26630 12002 26682
rect 12002 26630 12012 26682
rect 12036 26630 12066 26682
rect 12066 26630 12078 26682
rect 12078 26630 12092 26682
rect 12116 26630 12130 26682
rect 12130 26630 12142 26682
rect 12142 26630 12172 26682
rect 12196 26630 12206 26682
rect 12206 26630 12252 26682
rect 11956 26628 12012 26630
rect 12036 26628 12092 26630
rect 12116 26628 12172 26630
rect 12196 26628 12252 26630
rect 11956 25594 12012 25596
rect 12036 25594 12092 25596
rect 12116 25594 12172 25596
rect 12196 25594 12252 25596
rect 11956 25542 12002 25594
rect 12002 25542 12012 25594
rect 12036 25542 12066 25594
rect 12066 25542 12078 25594
rect 12078 25542 12092 25594
rect 12116 25542 12130 25594
rect 12130 25542 12142 25594
rect 12142 25542 12172 25594
rect 12196 25542 12206 25594
rect 12206 25542 12252 25594
rect 11956 25540 12012 25542
rect 12036 25540 12092 25542
rect 12116 25540 12172 25542
rect 12196 25540 12252 25542
rect 11956 24506 12012 24508
rect 12036 24506 12092 24508
rect 12116 24506 12172 24508
rect 12196 24506 12252 24508
rect 11956 24454 12002 24506
rect 12002 24454 12012 24506
rect 12036 24454 12066 24506
rect 12066 24454 12078 24506
rect 12078 24454 12092 24506
rect 12116 24454 12130 24506
rect 12130 24454 12142 24506
rect 12142 24454 12172 24506
rect 12196 24454 12206 24506
rect 12206 24454 12252 24506
rect 11956 24452 12012 24454
rect 12036 24452 12092 24454
rect 12116 24452 12172 24454
rect 12196 24452 12252 24454
rect 12616 42458 12672 42460
rect 12696 42458 12752 42460
rect 12776 42458 12832 42460
rect 12856 42458 12912 42460
rect 12616 42406 12662 42458
rect 12662 42406 12672 42458
rect 12696 42406 12726 42458
rect 12726 42406 12738 42458
rect 12738 42406 12752 42458
rect 12776 42406 12790 42458
rect 12790 42406 12802 42458
rect 12802 42406 12832 42458
rect 12856 42406 12866 42458
rect 12866 42406 12912 42458
rect 12616 42404 12672 42406
rect 12696 42404 12752 42406
rect 12776 42404 12832 42406
rect 12856 42404 12912 42406
rect 12616 41370 12672 41372
rect 12696 41370 12752 41372
rect 12776 41370 12832 41372
rect 12856 41370 12912 41372
rect 12616 41318 12662 41370
rect 12662 41318 12672 41370
rect 12696 41318 12726 41370
rect 12726 41318 12738 41370
rect 12738 41318 12752 41370
rect 12776 41318 12790 41370
rect 12790 41318 12802 41370
rect 12802 41318 12832 41370
rect 12856 41318 12866 41370
rect 12866 41318 12912 41370
rect 12616 41316 12672 41318
rect 12696 41316 12752 41318
rect 12776 41316 12832 41318
rect 12856 41316 12912 41318
rect 12616 40282 12672 40284
rect 12696 40282 12752 40284
rect 12776 40282 12832 40284
rect 12856 40282 12912 40284
rect 12616 40230 12662 40282
rect 12662 40230 12672 40282
rect 12696 40230 12726 40282
rect 12726 40230 12738 40282
rect 12738 40230 12752 40282
rect 12776 40230 12790 40282
rect 12790 40230 12802 40282
rect 12802 40230 12832 40282
rect 12856 40230 12866 40282
rect 12866 40230 12912 40282
rect 12616 40228 12672 40230
rect 12696 40228 12752 40230
rect 12776 40228 12832 40230
rect 12856 40228 12912 40230
rect 12616 39194 12672 39196
rect 12696 39194 12752 39196
rect 12776 39194 12832 39196
rect 12856 39194 12912 39196
rect 12616 39142 12662 39194
rect 12662 39142 12672 39194
rect 12696 39142 12726 39194
rect 12726 39142 12738 39194
rect 12738 39142 12752 39194
rect 12776 39142 12790 39194
rect 12790 39142 12802 39194
rect 12802 39142 12832 39194
rect 12856 39142 12866 39194
rect 12866 39142 12912 39194
rect 12616 39140 12672 39142
rect 12696 39140 12752 39142
rect 12776 39140 12832 39142
rect 12856 39140 12912 39142
rect 12616 38106 12672 38108
rect 12696 38106 12752 38108
rect 12776 38106 12832 38108
rect 12856 38106 12912 38108
rect 12616 38054 12662 38106
rect 12662 38054 12672 38106
rect 12696 38054 12726 38106
rect 12726 38054 12738 38106
rect 12738 38054 12752 38106
rect 12776 38054 12790 38106
rect 12790 38054 12802 38106
rect 12802 38054 12832 38106
rect 12856 38054 12866 38106
rect 12866 38054 12912 38106
rect 12616 38052 12672 38054
rect 12696 38052 12752 38054
rect 12776 38052 12832 38054
rect 12856 38052 12912 38054
rect 12616 37018 12672 37020
rect 12696 37018 12752 37020
rect 12776 37018 12832 37020
rect 12856 37018 12912 37020
rect 12616 36966 12662 37018
rect 12662 36966 12672 37018
rect 12696 36966 12726 37018
rect 12726 36966 12738 37018
rect 12738 36966 12752 37018
rect 12776 36966 12790 37018
rect 12790 36966 12802 37018
rect 12802 36966 12832 37018
rect 12856 36966 12866 37018
rect 12866 36966 12912 37018
rect 12616 36964 12672 36966
rect 12696 36964 12752 36966
rect 12776 36964 12832 36966
rect 12856 36964 12912 36966
rect 12616 35930 12672 35932
rect 12696 35930 12752 35932
rect 12776 35930 12832 35932
rect 12856 35930 12912 35932
rect 12616 35878 12662 35930
rect 12662 35878 12672 35930
rect 12696 35878 12726 35930
rect 12726 35878 12738 35930
rect 12738 35878 12752 35930
rect 12776 35878 12790 35930
rect 12790 35878 12802 35930
rect 12802 35878 12832 35930
rect 12856 35878 12866 35930
rect 12866 35878 12912 35930
rect 12616 35876 12672 35878
rect 12696 35876 12752 35878
rect 12776 35876 12832 35878
rect 12856 35876 12912 35878
rect 11956 23418 12012 23420
rect 12036 23418 12092 23420
rect 12116 23418 12172 23420
rect 12196 23418 12252 23420
rect 11956 23366 12002 23418
rect 12002 23366 12012 23418
rect 12036 23366 12066 23418
rect 12066 23366 12078 23418
rect 12078 23366 12092 23418
rect 12116 23366 12130 23418
rect 12130 23366 12142 23418
rect 12142 23366 12172 23418
rect 12196 23366 12206 23418
rect 12206 23366 12252 23418
rect 11956 23364 12012 23366
rect 12036 23364 12092 23366
rect 12116 23364 12172 23366
rect 12196 23364 12252 23366
rect 11956 22330 12012 22332
rect 12036 22330 12092 22332
rect 12116 22330 12172 22332
rect 12196 22330 12252 22332
rect 11956 22278 12002 22330
rect 12002 22278 12012 22330
rect 12036 22278 12066 22330
rect 12066 22278 12078 22330
rect 12078 22278 12092 22330
rect 12116 22278 12130 22330
rect 12130 22278 12142 22330
rect 12142 22278 12172 22330
rect 12196 22278 12206 22330
rect 12206 22278 12252 22330
rect 11956 22276 12012 22278
rect 12036 22276 12092 22278
rect 12116 22276 12172 22278
rect 12196 22276 12252 22278
rect 11956 21242 12012 21244
rect 12036 21242 12092 21244
rect 12116 21242 12172 21244
rect 12196 21242 12252 21244
rect 11956 21190 12002 21242
rect 12002 21190 12012 21242
rect 12036 21190 12066 21242
rect 12066 21190 12078 21242
rect 12078 21190 12092 21242
rect 12116 21190 12130 21242
rect 12130 21190 12142 21242
rect 12142 21190 12172 21242
rect 12196 21190 12206 21242
rect 12206 21190 12252 21242
rect 11956 21188 12012 21190
rect 12036 21188 12092 21190
rect 12116 21188 12172 21190
rect 12196 21188 12252 21190
rect 11956 20154 12012 20156
rect 12036 20154 12092 20156
rect 12116 20154 12172 20156
rect 12196 20154 12252 20156
rect 11956 20102 12002 20154
rect 12002 20102 12012 20154
rect 12036 20102 12066 20154
rect 12066 20102 12078 20154
rect 12078 20102 12092 20154
rect 12116 20102 12130 20154
rect 12130 20102 12142 20154
rect 12142 20102 12172 20154
rect 12196 20102 12206 20154
rect 12206 20102 12252 20154
rect 11956 20100 12012 20102
rect 12036 20100 12092 20102
rect 12116 20100 12172 20102
rect 12196 20100 12252 20102
rect 11956 19066 12012 19068
rect 12036 19066 12092 19068
rect 12116 19066 12172 19068
rect 12196 19066 12252 19068
rect 11956 19014 12002 19066
rect 12002 19014 12012 19066
rect 12036 19014 12066 19066
rect 12066 19014 12078 19066
rect 12078 19014 12092 19066
rect 12116 19014 12130 19066
rect 12130 19014 12142 19066
rect 12142 19014 12172 19066
rect 12196 19014 12206 19066
rect 12206 19014 12252 19066
rect 11956 19012 12012 19014
rect 12036 19012 12092 19014
rect 12116 19012 12172 19014
rect 12196 19012 12252 19014
rect 11956 17978 12012 17980
rect 12036 17978 12092 17980
rect 12116 17978 12172 17980
rect 12196 17978 12252 17980
rect 11956 17926 12002 17978
rect 12002 17926 12012 17978
rect 12036 17926 12066 17978
rect 12066 17926 12078 17978
rect 12078 17926 12092 17978
rect 12116 17926 12130 17978
rect 12130 17926 12142 17978
rect 12142 17926 12172 17978
rect 12196 17926 12206 17978
rect 12206 17926 12252 17978
rect 11956 17924 12012 17926
rect 12036 17924 12092 17926
rect 12116 17924 12172 17926
rect 12196 17924 12252 17926
rect 11956 16890 12012 16892
rect 12036 16890 12092 16892
rect 12116 16890 12172 16892
rect 12196 16890 12252 16892
rect 11956 16838 12002 16890
rect 12002 16838 12012 16890
rect 12036 16838 12066 16890
rect 12066 16838 12078 16890
rect 12078 16838 12092 16890
rect 12116 16838 12130 16890
rect 12130 16838 12142 16890
rect 12142 16838 12172 16890
rect 12196 16838 12206 16890
rect 12206 16838 12252 16890
rect 11956 16836 12012 16838
rect 12036 16836 12092 16838
rect 12116 16836 12172 16838
rect 12196 16836 12252 16838
rect 11956 15802 12012 15804
rect 12036 15802 12092 15804
rect 12116 15802 12172 15804
rect 12196 15802 12252 15804
rect 11956 15750 12002 15802
rect 12002 15750 12012 15802
rect 12036 15750 12066 15802
rect 12066 15750 12078 15802
rect 12078 15750 12092 15802
rect 12116 15750 12130 15802
rect 12130 15750 12142 15802
rect 12142 15750 12172 15802
rect 12196 15750 12206 15802
rect 12206 15750 12252 15802
rect 11956 15748 12012 15750
rect 12036 15748 12092 15750
rect 12116 15748 12172 15750
rect 12196 15748 12252 15750
rect 11956 14714 12012 14716
rect 12036 14714 12092 14716
rect 12116 14714 12172 14716
rect 12196 14714 12252 14716
rect 11956 14662 12002 14714
rect 12002 14662 12012 14714
rect 12036 14662 12066 14714
rect 12066 14662 12078 14714
rect 12078 14662 12092 14714
rect 12116 14662 12130 14714
rect 12130 14662 12142 14714
rect 12142 14662 12172 14714
rect 12196 14662 12206 14714
rect 12206 14662 12252 14714
rect 11956 14660 12012 14662
rect 12036 14660 12092 14662
rect 12116 14660 12172 14662
rect 12196 14660 12252 14662
rect 11956 13626 12012 13628
rect 12036 13626 12092 13628
rect 12116 13626 12172 13628
rect 12196 13626 12252 13628
rect 11956 13574 12002 13626
rect 12002 13574 12012 13626
rect 12036 13574 12066 13626
rect 12066 13574 12078 13626
rect 12078 13574 12092 13626
rect 12116 13574 12130 13626
rect 12130 13574 12142 13626
rect 12142 13574 12172 13626
rect 12196 13574 12206 13626
rect 12206 13574 12252 13626
rect 11956 13572 12012 13574
rect 12036 13572 12092 13574
rect 12116 13572 12172 13574
rect 12196 13572 12252 13574
rect 11956 12538 12012 12540
rect 12036 12538 12092 12540
rect 12116 12538 12172 12540
rect 12196 12538 12252 12540
rect 11956 12486 12002 12538
rect 12002 12486 12012 12538
rect 12036 12486 12066 12538
rect 12066 12486 12078 12538
rect 12078 12486 12092 12538
rect 12116 12486 12130 12538
rect 12130 12486 12142 12538
rect 12142 12486 12172 12538
rect 12196 12486 12206 12538
rect 12206 12486 12252 12538
rect 11956 12484 12012 12486
rect 12036 12484 12092 12486
rect 12116 12484 12172 12486
rect 12196 12484 12252 12486
rect 11956 11450 12012 11452
rect 12036 11450 12092 11452
rect 12116 11450 12172 11452
rect 12196 11450 12252 11452
rect 11956 11398 12002 11450
rect 12002 11398 12012 11450
rect 12036 11398 12066 11450
rect 12066 11398 12078 11450
rect 12078 11398 12092 11450
rect 12116 11398 12130 11450
rect 12130 11398 12142 11450
rect 12142 11398 12172 11450
rect 12196 11398 12206 11450
rect 12206 11398 12252 11450
rect 11956 11396 12012 11398
rect 12036 11396 12092 11398
rect 12116 11396 12172 11398
rect 12196 11396 12252 11398
rect 12616 34842 12672 34844
rect 12696 34842 12752 34844
rect 12776 34842 12832 34844
rect 12856 34842 12912 34844
rect 12616 34790 12662 34842
rect 12662 34790 12672 34842
rect 12696 34790 12726 34842
rect 12726 34790 12738 34842
rect 12738 34790 12752 34842
rect 12776 34790 12790 34842
rect 12790 34790 12802 34842
rect 12802 34790 12832 34842
rect 12856 34790 12866 34842
rect 12866 34790 12912 34842
rect 12616 34788 12672 34790
rect 12696 34788 12752 34790
rect 12776 34788 12832 34790
rect 12856 34788 12912 34790
rect 12616 33754 12672 33756
rect 12696 33754 12752 33756
rect 12776 33754 12832 33756
rect 12856 33754 12912 33756
rect 12616 33702 12662 33754
rect 12662 33702 12672 33754
rect 12696 33702 12726 33754
rect 12726 33702 12738 33754
rect 12738 33702 12752 33754
rect 12776 33702 12790 33754
rect 12790 33702 12802 33754
rect 12802 33702 12832 33754
rect 12856 33702 12866 33754
rect 12866 33702 12912 33754
rect 12616 33700 12672 33702
rect 12696 33700 12752 33702
rect 12776 33700 12832 33702
rect 12856 33700 12912 33702
rect 12616 32666 12672 32668
rect 12696 32666 12752 32668
rect 12776 32666 12832 32668
rect 12856 32666 12912 32668
rect 12616 32614 12662 32666
rect 12662 32614 12672 32666
rect 12696 32614 12726 32666
rect 12726 32614 12738 32666
rect 12738 32614 12752 32666
rect 12776 32614 12790 32666
rect 12790 32614 12802 32666
rect 12802 32614 12832 32666
rect 12856 32614 12866 32666
rect 12866 32614 12912 32666
rect 12616 32612 12672 32614
rect 12696 32612 12752 32614
rect 12776 32612 12832 32614
rect 12856 32612 12912 32614
rect 12616 31578 12672 31580
rect 12696 31578 12752 31580
rect 12776 31578 12832 31580
rect 12856 31578 12912 31580
rect 12616 31526 12662 31578
rect 12662 31526 12672 31578
rect 12696 31526 12726 31578
rect 12726 31526 12738 31578
rect 12738 31526 12752 31578
rect 12776 31526 12790 31578
rect 12790 31526 12802 31578
rect 12802 31526 12832 31578
rect 12856 31526 12866 31578
rect 12866 31526 12912 31578
rect 12616 31524 12672 31526
rect 12696 31524 12752 31526
rect 12776 31524 12832 31526
rect 12856 31524 12912 31526
rect 12616 30490 12672 30492
rect 12696 30490 12752 30492
rect 12776 30490 12832 30492
rect 12856 30490 12912 30492
rect 12616 30438 12662 30490
rect 12662 30438 12672 30490
rect 12696 30438 12726 30490
rect 12726 30438 12738 30490
rect 12738 30438 12752 30490
rect 12776 30438 12790 30490
rect 12790 30438 12802 30490
rect 12802 30438 12832 30490
rect 12856 30438 12866 30490
rect 12866 30438 12912 30490
rect 12616 30436 12672 30438
rect 12696 30436 12752 30438
rect 12776 30436 12832 30438
rect 12856 30436 12912 30438
rect 12616 29402 12672 29404
rect 12696 29402 12752 29404
rect 12776 29402 12832 29404
rect 12856 29402 12912 29404
rect 12616 29350 12662 29402
rect 12662 29350 12672 29402
rect 12696 29350 12726 29402
rect 12726 29350 12738 29402
rect 12738 29350 12752 29402
rect 12776 29350 12790 29402
rect 12790 29350 12802 29402
rect 12802 29350 12832 29402
rect 12856 29350 12866 29402
rect 12866 29350 12912 29402
rect 12616 29348 12672 29350
rect 12696 29348 12752 29350
rect 12776 29348 12832 29350
rect 12856 29348 12912 29350
rect 12616 28314 12672 28316
rect 12696 28314 12752 28316
rect 12776 28314 12832 28316
rect 12856 28314 12912 28316
rect 12616 28262 12662 28314
rect 12662 28262 12672 28314
rect 12696 28262 12726 28314
rect 12726 28262 12738 28314
rect 12738 28262 12752 28314
rect 12776 28262 12790 28314
rect 12790 28262 12802 28314
rect 12802 28262 12832 28314
rect 12856 28262 12866 28314
rect 12866 28262 12912 28314
rect 12616 28260 12672 28262
rect 12696 28260 12752 28262
rect 12776 28260 12832 28262
rect 12856 28260 12912 28262
rect 12616 27226 12672 27228
rect 12696 27226 12752 27228
rect 12776 27226 12832 27228
rect 12856 27226 12912 27228
rect 12616 27174 12662 27226
rect 12662 27174 12672 27226
rect 12696 27174 12726 27226
rect 12726 27174 12738 27226
rect 12738 27174 12752 27226
rect 12776 27174 12790 27226
rect 12790 27174 12802 27226
rect 12802 27174 12832 27226
rect 12856 27174 12866 27226
rect 12866 27174 12912 27226
rect 12616 27172 12672 27174
rect 12696 27172 12752 27174
rect 12776 27172 12832 27174
rect 12856 27172 12912 27174
rect 12616 26138 12672 26140
rect 12696 26138 12752 26140
rect 12776 26138 12832 26140
rect 12856 26138 12912 26140
rect 12616 26086 12662 26138
rect 12662 26086 12672 26138
rect 12696 26086 12726 26138
rect 12726 26086 12738 26138
rect 12738 26086 12752 26138
rect 12776 26086 12790 26138
rect 12790 26086 12802 26138
rect 12802 26086 12832 26138
rect 12856 26086 12866 26138
rect 12866 26086 12912 26138
rect 12616 26084 12672 26086
rect 12696 26084 12752 26086
rect 12776 26084 12832 26086
rect 12856 26084 12912 26086
rect 12616 25050 12672 25052
rect 12696 25050 12752 25052
rect 12776 25050 12832 25052
rect 12856 25050 12912 25052
rect 12616 24998 12662 25050
rect 12662 24998 12672 25050
rect 12696 24998 12726 25050
rect 12726 24998 12738 25050
rect 12738 24998 12752 25050
rect 12776 24998 12790 25050
rect 12790 24998 12802 25050
rect 12802 24998 12832 25050
rect 12856 24998 12866 25050
rect 12866 24998 12912 25050
rect 12616 24996 12672 24998
rect 12696 24996 12752 24998
rect 12776 24996 12832 24998
rect 12856 24996 12912 24998
rect 12616 23962 12672 23964
rect 12696 23962 12752 23964
rect 12776 23962 12832 23964
rect 12856 23962 12912 23964
rect 12616 23910 12662 23962
rect 12662 23910 12672 23962
rect 12696 23910 12726 23962
rect 12726 23910 12738 23962
rect 12738 23910 12752 23962
rect 12776 23910 12790 23962
rect 12790 23910 12802 23962
rect 12802 23910 12832 23962
rect 12856 23910 12866 23962
rect 12866 23910 12912 23962
rect 12616 23908 12672 23910
rect 12696 23908 12752 23910
rect 12776 23908 12832 23910
rect 12856 23908 12912 23910
rect 12616 22874 12672 22876
rect 12696 22874 12752 22876
rect 12776 22874 12832 22876
rect 12856 22874 12912 22876
rect 12616 22822 12662 22874
rect 12662 22822 12672 22874
rect 12696 22822 12726 22874
rect 12726 22822 12738 22874
rect 12738 22822 12752 22874
rect 12776 22822 12790 22874
rect 12790 22822 12802 22874
rect 12802 22822 12832 22874
rect 12856 22822 12866 22874
rect 12866 22822 12912 22874
rect 12616 22820 12672 22822
rect 12696 22820 12752 22822
rect 12776 22820 12832 22822
rect 12856 22820 12912 22822
rect 12616 21786 12672 21788
rect 12696 21786 12752 21788
rect 12776 21786 12832 21788
rect 12856 21786 12912 21788
rect 12616 21734 12662 21786
rect 12662 21734 12672 21786
rect 12696 21734 12726 21786
rect 12726 21734 12738 21786
rect 12738 21734 12752 21786
rect 12776 21734 12790 21786
rect 12790 21734 12802 21786
rect 12802 21734 12832 21786
rect 12856 21734 12866 21786
rect 12866 21734 12912 21786
rect 12616 21732 12672 21734
rect 12696 21732 12752 21734
rect 12776 21732 12832 21734
rect 12856 21732 12912 21734
rect 12616 20698 12672 20700
rect 12696 20698 12752 20700
rect 12776 20698 12832 20700
rect 12856 20698 12912 20700
rect 12616 20646 12662 20698
rect 12662 20646 12672 20698
rect 12696 20646 12726 20698
rect 12726 20646 12738 20698
rect 12738 20646 12752 20698
rect 12776 20646 12790 20698
rect 12790 20646 12802 20698
rect 12802 20646 12832 20698
rect 12856 20646 12866 20698
rect 12866 20646 12912 20698
rect 12616 20644 12672 20646
rect 12696 20644 12752 20646
rect 12776 20644 12832 20646
rect 12856 20644 12912 20646
rect 12616 19610 12672 19612
rect 12696 19610 12752 19612
rect 12776 19610 12832 19612
rect 12856 19610 12912 19612
rect 12616 19558 12662 19610
rect 12662 19558 12672 19610
rect 12696 19558 12726 19610
rect 12726 19558 12738 19610
rect 12738 19558 12752 19610
rect 12776 19558 12790 19610
rect 12790 19558 12802 19610
rect 12802 19558 12832 19610
rect 12856 19558 12866 19610
rect 12866 19558 12912 19610
rect 12616 19556 12672 19558
rect 12696 19556 12752 19558
rect 12776 19556 12832 19558
rect 12856 19556 12912 19558
rect 12616 18522 12672 18524
rect 12696 18522 12752 18524
rect 12776 18522 12832 18524
rect 12856 18522 12912 18524
rect 12616 18470 12662 18522
rect 12662 18470 12672 18522
rect 12696 18470 12726 18522
rect 12726 18470 12738 18522
rect 12738 18470 12752 18522
rect 12776 18470 12790 18522
rect 12790 18470 12802 18522
rect 12802 18470 12832 18522
rect 12856 18470 12866 18522
rect 12866 18470 12912 18522
rect 12616 18468 12672 18470
rect 12696 18468 12752 18470
rect 12776 18468 12832 18470
rect 12856 18468 12912 18470
rect 12616 17434 12672 17436
rect 12696 17434 12752 17436
rect 12776 17434 12832 17436
rect 12856 17434 12912 17436
rect 12616 17382 12662 17434
rect 12662 17382 12672 17434
rect 12696 17382 12726 17434
rect 12726 17382 12738 17434
rect 12738 17382 12752 17434
rect 12776 17382 12790 17434
rect 12790 17382 12802 17434
rect 12802 17382 12832 17434
rect 12856 17382 12866 17434
rect 12866 17382 12912 17434
rect 12616 17380 12672 17382
rect 12696 17380 12752 17382
rect 12776 17380 12832 17382
rect 12856 17380 12912 17382
rect 12616 16346 12672 16348
rect 12696 16346 12752 16348
rect 12776 16346 12832 16348
rect 12856 16346 12912 16348
rect 12616 16294 12662 16346
rect 12662 16294 12672 16346
rect 12696 16294 12726 16346
rect 12726 16294 12738 16346
rect 12738 16294 12752 16346
rect 12776 16294 12790 16346
rect 12790 16294 12802 16346
rect 12802 16294 12832 16346
rect 12856 16294 12866 16346
rect 12866 16294 12912 16346
rect 12616 16292 12672 16294
rect 12696 16292 12752 16294
rect 12776 16292 12832 16294
rect 12856 16292 12912 16294
rect 12616 15258 12672 15260
rect 12696 15258 12752 15260
rect 12776 15258 12832 15260
rect 12856 15258 12912 15260
rect 12616 15206 12662 15258
rect 12662 15206 12672 15258
rect 12696 15206 12726 15258
rect 12726 15206 12738 15258
rect 12738 15206 12752 15258
rect 12776 15206 12790 15258
rect 12790 15206 12802 15258
rect 12802 15206 12832 15258
rect 12856 15206 12866 15258
rect 12866 15206 12912 15258
rect 12616 15204 12672 15206
rect 12696 15204 12752 15206
rect 12776 15204 12832 15206
rect 12856 15204 12912 15206
rect 12616 14170 12672 14172
rect 12696 14170 12752 14172
rect 12776 14170 12832 14172
rect 12856 14170 12912 14172
rect 12616 14118 12662 14170
rect 12662 14118 12672 14170
rect 12696 14118 12726 14170
rect 12726 14118 12738 14170
rect 12738 14118 12752 14170
rect 12776 14118 12790 14170
rect 12790 14118 12802 14170
rect 12802 14118 12832 14170
rect 12856 14118 12866 14170
rect 12866 14118 12912 14170
rect 12616 14116 12672 14118
rect 12696 14116 12752 14118
rect 12776 14116 12832 14118
rect 12856 14116 12912 14118
rect 12616 13082 12672 13084
rect 12696 13082 12752 13084
rect 12776 13082 12832 13084
rect 12856 13082 12912 13084
rect 12616 13030 12662 13082
rect 12662 13030 12672 13082
rect 12696 13030 12726 13082
rect 12726 13030 12738 13082
rect 12738 13030 12752 13082
rect 12776 13030 12790 13082
rect 12790 13030 12802 13082
rect 12802 13030 12832 13082
rect 12856 13030 12866 13082
rect 12866 13030 12912 13082
rect 12616 13028 12672 13030
rect 12696 13028 12752 13030
rect 12776 13028 12832 13030
rect 12856 13028 12912 13030
rect 12616 11994 12672 11996
rect 12696 11994 12752 11996
rect 12776 11994 12832 11996
rect 12856 11994 12912 11996
rect 12616 11942 12662 11994
rect 12662 11942 12672 11994
rect 12696 11942 12726 11994
rect 12726 11942 12738 11994
rect 12738 11942 12752 11994
rect 12776 11942 12790 11994
rect 12790 11942 12802 11994
rect 12802 11942 12832 11994
rect 12856 11942 12866 11994
rect 12866 11942 12912 11994
rect 12616 11940 12672 11942
rect 12696 11940 12752 11942
rect 12776 11940 12832 11942
rect 12856 11940 12912 11942
rect 12616 10906 12672 10908
rect 12696 10906 12752 10908
rect 12776 10906 12832 10908
rect 12856 10906 12912 10908
rect 12616 10854 12662 10906
rect 12662 10854 12672 10906
rect 12696 10854 12726 10906
rect 12726 10854 12738 10906
rect 12738 10854 12752 10906
rect 12776 10854 12790 10906
rect 12790 10854 12802 10906
rect 12802 10854 12832 10906
rect 12856 10854 12866 10906
rect 12866 10854 12912 10906
rect 12616 10852 12672 10854
rect 12696 10852 12752 10854
rect 12776 10852 12832 10854
rect 12856 10852 12912 10854
rect 11956 10362 12012 10364
rect 12036 10362 12092 10364
rect 12116 10362 12172 10364
rect 12196 10362 12252 10364
rect 11956 10310 12002 10362
rect 12002 10310 12012 10362
rect 12036 10310 12066 10362
rect 12066 10310 12078 10362
rect 12078 10310 12092 10362
rect 12116 10310 12130 10362
rect 12130 10310 12142 10362
rect 12142 10310 12172 10362
rect 12196 10310 12206 10362
rect 12206 10310 12252 10362
rect 11956 10308 12012 10310
rect 12036 10308 12092 10310
rect 12116 10308 12172 10310
rect 12196 10308 12252 10310
rect 12616 9818 12672 9820
rect 12696 9818 12752 9820
rect 12776 9818 12832 9820
rect 12856 9818 12912 9820
rect 12616 9766 12662 9818
rect 12662 9766 12672 9818
rect 12696 9766 12726 9818
rect 12726 9766 12738 9818
rect 12738 9766 12752 9818
rect 12776 9766 12790 9818
rect 12790 9766 12802 9818
rect 12802 9766 12832 9818
rect 12856 9766 12866 9818
rect 12866 9766 12912 9818
rect 12616 9764 12672 9766
rect 12696 9764 12752 9766
rect 12776 9764 12832 9766
rect 12856 9764 12912 9766
rect 11956 9274 12012 9276
rect 12036 9274 12092 9276
rect 12116 9274 12172 9276
rect 12196 9274 12252 9276
rect 11956 9222 12002 9274
rect 12002 9222 12012 9274
rect 12036 9222 12066 9274
rect 12066 9222 12078 9274
rect 12078 9222 12092 9274
rect 12116 9222 12130 9274
rect 12130 9222 12142 9274
rect 12142 9222 12172 9274
rect 12196 9222 12206 9274
rect 12206 9222 12252 9274
rect 11956 9220 12012 9222
rect 12036 9220 12092 9222
rect 12116 9220 12172 9222
rect 12196 9220 12252 9222
rect 12616 8730 12672 8732
rect 12696 8730 12752 8732
rect 12776 8730 12832 8732
rect 12856 8730 12912 8732
rect 12616 8678 12662 8730
rect 12662 8678 12672 8730
rect 12696 8678 12726 8730
rect 12726 8678 12738 8730
rect 12738 8678 12752 8730
rect 12776 8678 12790 8730
rect 12790 8678 12802 8730
rect 12802 8678 12832 8730
rect 12856 8678 12866 8730
rect 12866 8678 12912 8730
rect 12616 8676 12672 8678
rect 12696 8676 12752 8678
rect 12776 8676 12832 8678
rect 12856 8676 12912 8678
rect 11956 8186 12012 8188
rect 12036 8186 12092 8188
rect 12116 8186 12172 8188
rect 12196 8186 12252 8188
rect 11956 8134 12002 8186
rect 12002 8134 12012 8186
rect 12036 8134 12066 8186
rect 12066 8134 12078 8186
rect 12078 8134 12092 8186
rect 12116 8134 12130 8186
rect 12130 8134 12142 8186
rect 12142 8134 12172 8186
rect 12196 8134 12206 8186
rect 12206 8134 12252 8186
rect 11956 8132 12012 8134
rect 12036 8132 12092 8134
rect 12116 8132 12172 8134
rect 12196 8132 12252 8134
rect 12616 7642 12672 7644
rect 12696 7642 12752 7644
rect 12776 7642 12832 7644
rect 12856 7642 12912 7644
rect 12616 7590 12662 7642
rect 12662 7590 12672 7642
rect 12696 7590 12726 7642
rect 12726 7590 12738 7642
rect 12738 7590 12752 7642
rect 12776 7590 12790 7642
rect 12790 7590 12802 7642
rect 12802 7590 12832 7642
rect 12856 7590 12866 7642
rect 12866 7590 12912 7642
rect 12616 7588 12672 7590
rect 12696 7588 12752 7590
rect 12776 7588 12832 7590
rect 12856 7588 12912 7590
rect 11956 7098 12012 7100
rect 12036 7098 12092 7100
rect 12116 7098 12172 7100
rect 12196 7098 12252 7100
rect 11956 7046 12002 7098
rect 12002 7046 12012 7098
rect 12036 7046 12066 7098
rect 12066 7046 12078 7098
rect 12078 7046 12092 7098
rect 12116 7046 12130 7098
rect 12130 7046 12142 7098
rect 12142 7046 12172 7098
rect 12196 7046 12206 7098
rect 12206 7046 12252 7098
rect 11956 7044 12012 7046
rect 12036 7044 12092 7046
rect 12116 7044 12172 7046
rect 12196 7044 12252 7046
rect 12616 6554 12672 6556
rect 12696 6554 12752 6556
rect 12776 6554 12832 6556
rect 12856 6554 12912 6556
rect 12616 6502 12662 6554
rect 12662 6502 12672 6554
rect 12696 6502 12726 6554
rect 12726 6502 12738 6554
rect 12738 6502 12752 6554
rect 12776 6502 12790 6554
rect 12790 6502 12802 6554
rect 12802 6502 12832 6554
rect 12856 6502 12866 6554
rect 12866 6502 12912 6554
rect 12616 6500 12672 6502
rect 12696 6500 12752 6502
rect 12776 6500 12832 6502
rect 12856 6500 12912 6502
rect 11956 6010 12012 6012
rect 12036 6010 12092 6012
rect 12116 6010 12172 6012
rect 12196 6010 12252 6012
rect 11956 5958 12002 6010
rect 12002 5958 12012 6010
rect 12036 5958 12066 6010
rect 12066 5958 12078 6010
rect 12078 5958 12092 6010
rect 12116 5958 12130 6010
rect 12130 5958 12142 6010
rect 12142 5958 12172 6010
rect 12196 5958 12206 6010
rect 12206 5958 12252 6010
rect 11956 5956 12012 5958
rect 12036 5956 12092 5958
rect 12116 5956 12172 5958
rect 12196 5956 12252 5958
rect 12616 5466 12672 5468
rect 12696 5466 12752 5468
rect 12776 5466 12832 5468
rect 12856 5466 12912 5468
rect 12616 5414 12662 5466
rect 12662 5414 12672 5466
rect 12696 5414 12726 5466
rect 12726 5414 12738 5466
rect 12738 5414 12752 5466
rect 12776 5414 12790 5466
rect 12790 5414 12802 5466
rect 12802 5414 12832 5466
rect 12856 5414 12866 5466
rect 12866 5414 12912 5466
rect 12616 5412 12672 5414
rect 12696 5412 12752 5414
rect 12776 5412 12832 5414
rect 12856 5412 12912 5414
rect 11956 4922 12012 4924
rect 12036 4922 12092 4924
rect 12116 4922 12172 4924
rect 12196 4922 12252 4924
rect 11956 4870 12002 4922
rect 12002 4870 12012 4922
rect 12036 4870 12066 4922
rect 12066 4870 12078 4922
rect 12078 4870 12092 4922
rect 12116 4870 12130 4922
rect 12130 4870 12142 4922
rect 12142 4870 12172 4922
rect 12196 4870 12206 4922
rect 12206 4870 12252 4922
rect 11956 4868 12012 4870
rect 12036 4868 12092 4870
rect 12116 4868 12172 4870
rect 12196 4868 12252 4870
rect 11956 3834 12012 3836
rect 12036 3834 12092 3836
rect 12116 3834 12172 3836
rect 12196 3834 12252 3836
rect 11956 3782 12002 3834
rect 12002 3782 12012 3834
rect 12036 3782 12066 3834
rect 12066 3782 12078 3834
rect 12078 3782 12092 3834
rect 12116 3782 12130 3834
rect 12130 3782 12142 3834
rect 12142 3782 12172 3834
rect 12196 3782 12206 3834
rect 12206 3782 12252 3834
rect 11956 3780 12012 3782
rect 12036 3780 12092 3782
rect 12116 3780 12172 3782
rect 12196 3780 12252 3782
rect 12616 4378 12672 4380
rect 12696 4378 12752 4380
rect 12776 4378 12832 4380
rect 12856 4378 12912 4380
rect 12616 4326 12662 4378
rect 12662 4326 12672 4378
rect 12696 4326 12726 4378
rect 12726 4326 12738 4378
rect 12738 4326 12752 4378
rect 12776 4326 12790 4378
rect 12790 4326 12802 4378
rect 12802 4326 12832 4378
rect 12856 4326 12866 4378
rect 12866 4326 12912 4378
rect 12616 4324 12672 4326
rect 12696 4324 12752 4326
rect 12776 4324 12832 4326
rect 12856 4324 12912 4326
rect 12616 3290 12672 3292
rect 12696 3290 12752 3292
rect 12776 3290 12832 3292
rect 12856 3290 12912 3292
rect 12616 3238 12662 3290
rect 12662 3238 12672 3290
rect 12696 3238 12726 3290
rect 12726 3238 12738 3290
rect 12738 3238 12752 3290
rect 12776 3238 12790 3290
rect 12790 3238 12802 3290
rect 12802 3238 12832 3290
rect 12856 3238 12866 3290
rect 12866 3238 12912 3290
rect 12616 3236 12672 3238
rect 12696 3236 12752 3238
rect 12776 3236 12832 3238
rect 12856 3236 12912 3238
rect 11956 2746 12012 2748
rect 12036 2746 12092 2748
rect 12116 2746 12172 2748
rect 12196 2746 12252 2748
rect 11956 2694 12002 2746
rect 12002 2694 12012 2746
rect 12036 2694 12066 2746
rect 12066 2694 12078 2746
rect 12078 2694 12092 2746
rect 12116 2694 12130 2746
rect 12130 2694 12142 2746
rect 12142 2694 12172 2746
rect 12196 2694 12206 2746
rect 12206 2694 12252 2746
rect 11956 2692 12012 2694
rect 12036 2692 12092 2694
rect 12116 2692 12172 2694
rect 12196 2692 12252 2694
rect 14922 22752 14978 22808
rect 17616 68570 17672 68572
rect 17696 68570 17752 68572
rect 17776 68570 17832 68572
rect 17856 68570 17912 68572
rect 17616 68518 17662 68570
rect 17662 68518 17672 68570
rect 17696 68518 17726 68570
rect 17726 68518 17738 68570
rect 17738 68518 17752 68570
rect 17776 68518 17790 68570
rect 17790 68518 17802 68570
rect 17802 68518 17832 68570
rect 17856 68518 17866 68570
rect 17866 68518 17912 68570
rect 17616 68516 17672 68518
rect 17696 68516 17752 68518
rect 17776 68516 17832 68518
rect 17856 68516 17912 68518
rect 16956 68026 17012 68028
rect 17036 68026 17092 68028
rect 17116 68026 17172 68028
rect 17196 68026 17252 68028
rect 16956 67974 17002 68026
rect 17002 67974 17012 68026
rect 17036 67974 17066 68026
rect 17066 67974 17078 68026
rect 17078 67974 17092 68026
rect 17116 67974 17130 68026
rect 17130 67974 17142 68026
rect 17142 67974 17172 68026
rect 17196 67974 17206 68026
rect 17206 67974 17252 68026
rect 16956 67972 17012 67974
rect 17036 67972 17092 67974
rect 17116 67972 17172 67974
rect 17196 67972 17252 67974
rect 17616 67482 17672 67484
rect 17696 67482 17752 67484
rect 17776 67482 17832 67484
rect 17856 67482 17912 67484
rect 17616 67430 17662 67482
rect 17662 67430 17672 67482
rect 17696 67430 17726 67482
rect 17726 67430 17738 67482
rect 17738 67430 17752 67482
rect 17776 67430 17790 67482
rect 17790 67430 17802 67482
rect 17802 67430 17832 67482
rect 17856 67430 17866 67482
rect 17866 67430 17912 67482
rect 17616 67428 17672 67430
rect 17696 67428 17752 67430
rect 17776 67428 17832 67430
rect 17856 67428 17912 67430
rect 16956 66938 17012 66940
rect 17036 66938 17092 66940
rect 17116 66938 17172 66940
rect 17196 66938 17252 66940
rect 16956 66886 17002 66938
rect 17002 66886 17012 66938
rect 17036 66886 17066 66938
rect 17066 66886 17078 66938
rect 17078 66886 17092 66938
rect 17116 66886 17130 66938
rect 17130 66886 17142 66938
rect 17142 66886 17172 66938
rect 17196 66886 17206 66938
rect 17206 66886 17252 66938
rect 16956 66884 17012 66886
rect 17036 66884 17092 66886
rect 17116 66884 17172 66886
rect 17196 66884 17252 66886
rect 17616 66394 17672 66396
rect 17696 66394 17752 66396
rect 17776 66394 17832 66396
rect 17856 66394 17912 66396
rect 17616 66342 17662 66394
rect 17662 66342 17672 66394
rect 17696 66342 17726 66394
rect 17726 66342 17738 66394
rect 17738 66342 17752 66394
rect 17776 66342 17790 66394
rect 17790 66342 17802 66394
rect 17802 66342 17832 66394
rect 17856 66342 17866 66394
rect 17866 66342 17912 66394
rect 17616 66340 17672 66342
rect 17696 66340 17752 66342
rect 17776 66340 17832 66342
rect 17856 66340 17912 66342
rect 16956 65850 17012 65852
rect 17036 65850 17092 65852
rect 17116 65850 17172 65852
rect 17196 65850 17252 65852
rect 16956 65798 17002 65850
rect 17002 65798 17012 65850
rect 17036 65798 17066 65850
rect 17066 65798 17078 65850
rect 17078 65798 17092 65850
rect 17116 65798 17130 65850
rect 17130 65798 17142 65850
rect 17142 65798 17172 65850
rect 17196 65798 17206 65850
rect 17206 65798 17252 65850
rect 16956 65796 17012 65798
rect 17036 65796 17092 65798
rect 17116 65796 17172 65798
rect 17196 65796 17252 65798
rect 17616 65306 17672 65308
rect 17696 65306 17752 65308
rect 17776 65306 17832 65308
rect 17856 65306 17912 65308
rect 17616 65254 17662 65306
rect 17662 65254 17672 65306
rect 17696 65254 17726 65306
rect 17726 65254 17738 65306
rect 17738 65254 17752 65306
rect 17776 65254 17790 65306
rect 17790 65254 17802 65306
rect 17802 65254 17832 65306
rect 17856 65254 17866 65306
rect 17866 65254 17912 65306
rect 17616 65252 17672 65254
rect 17696 65252 17752 65254
rect 17776 65252 17832 65254
rect 17856 65252 17912 65254
rect 16956 64762 17012 64764
rect 17036 64762 17092 64764
rect 17116 64762 17172 64764
rect 17196 64762 17252 64764
rect 16956 64710 17002 64762
rect 17002 64710 17012 64762
rect 17036 64710 17066 64762
rect 17066 64710 17078 64762
rect 17078 64710 17092 64762
rect 17116 64710 17130 64762
rect 17130 64710 17142 64762
rect 17142 64710 17172 64762
rect 17196 64710 17206 64762
rect 17206 64710 17252 64762
rect 16956 64708 17012 64710
rect 17036 64708 17092 64710
rect 17116 64708 17172 64710
rect 17196 64708 17252 64710
rect 16956 63674 17012 63676
rect 17036 63674 17092 63676
rect 17116 63674 17172 63676
rect 17196 63674 17252 63676
rect 16956 63622 17002 63674
rect 17002 63622 17012 63674
rect 17036 63622 17066 63674
rect 17066 63622 17078 63674
rect 17078 63622 17092 63674
rect 17116 63622 17130 63674
rect 17130 63622 17142 63674
rect 17142 63622 17172 63674
rect 17196 63622 17206 63674
rect 17206 63622 17252 63674
rect 16956 63620 17012 63622
rect 17036 63620 17092 63622
rect 17116 63620 17172 63622
rect 17196 63620 17252 63622
rect 15198 35128 15254 35184
rect 16486 55256 16542 55312
rect 16956 62586 17012 62588
rect 17036 62586 17092 62588
rect 17116 62586 17172 62588
rect 17196 62586 17252 62588
rect 16956 62534 17002 62586
rect 17002 62534 17012 62586
rect 17036 62534 17066 62586
rect 17066 62534 17078 62586
rect 17078 62534 17092 62586
rect 17116 62534 17130 62586
rect 17130 62534 17142 62586
rect 17142 62534 17172 62586
rect 17196 62534 17206 62586
rect 17206 62534 17252 62586
rect 16956 62532 17012 62534
rect 17036 62532 17092 62534
rect 17116 62532 17172 62534
rect 17196 62532 17252 62534
rect 16956 61498 17012 61500
rect 17036 61498 17092 61500
rect 17116 61498 17172 61500
rect 17196 61498 17252 61500
rect 16956 61446 17002 61498
rect 17002 61446 17012 61498
rect 17036 61446 17066 61498
rect 17066 61446 17078 61498
rect 17078 61446 17092 61498
rect 17116 61446 17130 61498
rect 17130 61446 17142 61498
rect 17142 61446 17172 61498
rect 17196 61446 17206 61498
rect 17206 61446 17252 61498
rect 16956 61444 17012 61446
rect 17036 61444 17092 61446
rect 17116 61444 17172 61446
rect 17196 61444 17252 61446
rect 16956 60410 17012 60412
rect 17036 60410 17092 60412
rect 17116 60410 17172 60412
rect 17196 60410 17252 60412
rect 16956 60358 17002 60410
rect 17002 60358 17012 60410
rect 17036 60358 17066 60410
rect 17066 60358 17078 60410
rect 17078 60358 17092 60410
rect 17116 60358 17130 60410
rect 17130 60358 17142 60410
rect 17142 60358 17172 60410
rect 17196 60358 17206 60410
rect 17206 60358 17252 60410
rect 16956 60356 17012 60358
rect 17036 60356 17092 60358
rect 17116 60356 17172 60358
rect 17196 60356 17252 60358
rect 16956 59322 17012 59324
rect 17036 59322 17092 59324
rect 17116 59322 17172 59324
rect 17196 59322 17252 59324
rect 16956 59270 17002 59322
rect 17002 59270 17012 59322
rect 17036 59270 17066 59322
rect 17066 59270 17078 59322
rect 17078 59270 17092 59322
rect 17116 59270 17130 59322
rect 17130 59270 17142 59322
rect 17142 59270 17172 59322
rect 17196 59270 17206 59322
rect 17206 59270 17252 59322
rect 16956 59268 17012 59270
rect 17036 59268 17092 59270
rect 17116 59268 17172 59270
rect 17196 59268 17252 59270
rect 16956 58234 17012 58236
rect 17036 58234 17092 58236
rect 17116 58234 17172 58236
rect 17196 58234 17252 58236
rect 16956 58182 17002 58234
rect 17002 58182 17012 58234
rect 17036 58182 17066 58234
rect 17066 58182 17078 58234
rect 17078 58182 17092 58234
rect 17116 58182 17130 58234
rect 17130 58182 17142 58234
rect 17142 58182 17172 58234
rect 17196 58182 17206 58234
rect 17206 58182 17252 58234
rect 16956 58180 17012 58182
rect 17036 58180 17092 58182
rect 17116 58180 17172 58182
rect 17196 58180 17252 58182
rect 16956 57146 17012 57148
rect 17036 57146 17092 57148
rect 17116 57146 17172 57148
rect 17196 57146 17252 57148
rect 16956 57094 17002 57146
rect 17002 57094 17012 57146
rect 17036 57094 17066 57146
rect 17066 57094 17078 57146
rect 17078 57094 17092 57146
rect 17116 57094 17130 57146
rect 17130 57094 17142 57146
rect 17142 57094 17172 57146
rect 17196 57094 17206 57146
rect 17206 57094 17252 57146
rect 16956 57092 17012 57094
rect 17036 57092 17092 57094
rect 17116 57092 17172 57094
rect 17196 57092 17252 57094
rect 16956 56058 17012 56060
rect 17036 56058 17092 56060
rect 17116 56058 17172 56060
rect 17196 56058 17252 56060
rect 16956 56006 17002 56058
rect 17002 56006 17012 56058
rect 17036 56006 17066 56058
rect 17066 56006 17078 56058
rect 17078 56006 17092 56058
rect 17116 56006 17130 56058
rect 17130 56006 17142 56058
rect 17142 56006 17172 56058
rect 17196 56006 17206 56058
rect 17206 56006 17252 56058
rect 16956 56004 17012 56006
rect 17036 56004 17092 56006
rect 17116 56004 17172 56006
rect 17196 56004 17252 56006
rect 16956 54970 17012 54972
rect 17036 54970 17092 54972
rect 17116 54970 17172 54972
rect 17196 54970 17252 54972
rect 16956 54918 17002 54970
rect 17002 54918 17012 54970
rect 17036 54918 17066 54970
rect 17066 54918 17078 54970
rect 17078 54918 17092 54970
rect 17116 54918 17130 54970
rect 17130 54918 17142 54970
rect 17142 54918 17172 54970
rect 17196 54918 17206 54970
rect 17206 54918 17252 54970
rect 16956 54916 17012 54918
rect 17036 54916 17092 54918
rect 17116 54916 17172 54918
rect 17196 54916 17252 54918
rect 16956 53882 17012 53884
rect 17036 53882 17092 53884
rect 17116 53882 17172 53884
rect 17196 53882 17252 53884
rect 16956 53830 17002 53882
rect 17002 53830 17012 53882
rect 17036 53830 17066 53882
rect 17066 53830 17078 53882
rect 17078 53830 17092 53882
rect 17116 53830 17130 53882
rect 17130 53830 17142 53882
rect 17142 53830 17172 53882
rect 17196 53830 17206 53882
rect 17206 53830 17252 53882
rect 16956 53828 17012 53830
rect 17036 53828 17092 53830
rect 17116 53828 17172 53830
rect 17196 53828 17252 53830
rect 16956 52794 17012 52796
rect 17036 52794 17092 52796
rect 17116 52794 17172 52796
rect 17196 52794 17252 52796
rect 16956 52742 17002 52794
rect 17002 52742 17012 52794
rect 17036 52742 17066 52794
rect 17066 52742 17078 52794
rect 17078 52742 17092 52794
rect 17116 52742 17130 52794
rect 17130 52742 17142 52794
rect 17142 52742 17172 52794
rect 17196 52742 17206 52794
rect 17206 52742 17252 52794
rect 16956 52740 17012 52742
rect 17036 52740 17092 52742
rect 17116 52740 17172 52742
rect 17196 52740 17252 52742
rect 16956 51706 17012 51708
rect 17036 51706 17092 51708
rect 17116 51706 17172 51708
rect 17196 51706 17252 51708
rect 16956 51654 17002 51706
rect 17002 51654 17012 51706
rect 17036 51654 17066 51706
rect 17066 51654 17078 51706
rect 17078 51654 17092 51706
rect 17116 51654 17130 51706
rect 17130 51654 17142 51706
rect 17142 51654 17172 51706
rect 17196 51654 17206 51706
rect 17206 51654 17252 51706
rect 16956 51652 17012 51654
rect 17036 51652 17092 51654
rect 17116 51652 17172 51654
rect 17196 51652 17252 51654
rect 16956 50618 17012 50620
rect 17036 50618 17092 50620
rect 17116 50618 17172 50620
rect 17196 50618 17252 50620
rect 16956 50566 17002 50618
rect 17002 50566 17012 50618
rect 17036 50566 17066 50618
rect 17066 50566 17078 50618
rect 17078 50566 17092 50618
rect 17116 50566 17130 50618
rect 17130 50566 17142 50618
rect 17142 50566 17172 50618
rect 17196 50566 17206 50618
rect 17206 50566 17252 50618
rect 16956 50564 17012 50566
rect 17036 50564 17092 50566
rect 17116 50564 17172 50566
rect 17196 50564 17252 50566
rect 16956 49530 17012 49532
rect 17036 49530 17092 49532
rect 17116 49530 17172 49532
rect 17196 49530 17252 49532
rect 16956 49478 17002 49530
rect 17002 49478 17012 49530
rect 17036 49478 17066 49530
rect 17066 49478 17078 49530
rect 17078 49478 17092 49530
rect 17116 49478 17130 49530
rect 17130 49478 17142 49530
rect 17142 49478 17172 49530
rect 17196 49478 17206 49530
rect 17206 49478 17252 49530
rect 16956 49476 17012 49478
rect 17036 49476 17092 49478
rect 17116 49476 17172 49478
rect 17196 49476 17252 49478
rect 17616 64218 17672 64220
rect 17696 64218 17752 64220
rect 17776 64218 17832 64220
rect 17856 64218 17912 64220
rect 17616 64166 17662 64218
rect 17662 64166 17672 64218
rect 17696 64166 17726 64218
rect 17726 64166 17738 64218
rect 17738 64166 17752 64218
rect 17776 64166 17790 64218
rect 17790 64166 17802 64218
rect 17802 64166 17832 64218
rect 17856 64166 17866 64218
rect 17866 64166 17912 64218
rect 17616 64164 17672 64166
rect 17696 64164 17752 64166
rect 17776 64164 17832 64166
rect 17856 64164 17912 64166
rect 17616 63130 17672 63132
rect 17696 63130 17752 63132
rect 17776 63130 17832 63132
rect 17856 63130 17912 63132
rect 17616 63078 17662 63130
rect 17662 63078 17672 63130
rect 17696 63078 17726 63130
rect 17726 63078 17738 63130
rect 17738 63078 17752 63130
rect 17776 63078 17790 63130
rect 17790 63078 17802 63130
rect 17802 63078 17832 63130
rect 17856 63078 17866 63130
rect 17866 63078 17912 63130
rect 17616 63076 17672 63078
rect 17696 63076 17752 63078
rect 17776 63076 17832 63078
rect 17856 63076 17912 63078
rect 17616 62042 17672 62044
rect 17696 62042 17752 62044
rect 17776 62042 17832 62044
rect 17856 62042 17912 62044
rect 17616 61990 17662 62042
rect 17662 61990 17672 62042
rect 17696 61990 17726 62042
rect 17726 61990 17738 62042
rect 17738 61990 17752 62042
rect 17776 61990 17790 62042
rect 17790 61990 17802 62042
rect 17802 61990 17832 62042
rect 17856 61990 17866 62042
rect 17866 61990 17912 62042
rect 17616 61988 17672 61990
rect 17696 61988 17752 61990
rect 17776 61988 17832 61990
rect 17856 61988 17912 61990
rect 17616 60954 17672 60956
rect 17696 60954 17752 60956
rect 17776 60954 17832 60956
rect 17856 60954 17912 60956
rect 17616 60902 17662 60954
rect 17662 60902 17672 60954
rect 17696 60902 17726 60954
rect 17726 60902 17738 60954
rect 17738 60902 17752 60954
rect 17776 60902 17790 60954
rect 17790 60902 17802 60954
rect 17802 60902 17832 60954
rect 17856 60902 17866 60954
rect 17866 60902 17912 60954
rect 17616 60900 17672 60902
rect 17696 60900 17752 60902
rect 17776 60900 17832 60902
rect 17856 60900 17912 60902
rect 17616 59866 17672 59868
rect 17696 59866 17752 59868
rect 17776 59866 17832 59868
rect 17856 59866 17912 59868
rect 17616 59814 17662 59866
rect 17662 59814 17672 59866
rect 17696 59814 17726 59866
rect 17726 59814 17738 59866
rect 17738 59814 17752 59866
rect 17776 59814 17790 59866
rect 17790 59814 17802 59866
rect 17802 59814 17832 59866
rect 17856 59814 17866 59866
rect 17866 59814 17912 59866
rect 17616 59812 17672 59814
rect 17696 59812 17752 59814
rect 17776 59812 17832 59814
rect 17856 59812 17912 59814
rect 17616 58778 17672 58780
rect 17696 58778 17752 58780
rect 17776 58778 17832 58780
rect 17856 58778 17912 58780
rect 17616 58726 17662 58778
rect 17662 58726 17672 58778
rect 17696 58726 17726 58778
rect 17726 58726 17738 58778
rect 17738 58726 17752 58778
rect 17776 58726 17790 58778
rect 17790 58726 17802 58778
rect 17802 58726 17832 58778
rect 17856 58726 17866 58778
rect 17866 58726 17912 58778
rect 17616 58724 17672 58726
rect 17696 58724 17752 58726
rect 17776 58724 17832 58726
rect 17856 58724 17912 58726
rect 17616 57690 17672 57692
rect 17696 57690 17752 57692
rect 17776 57690 17832 57692
rect 17856 57690 17912 57692
rect 17616 57638 17662 57690
rect 17662 57638 17672 57690
rect 17696 57638 17726 57690
rect 17726 57638 17738 57690
rect 17738 57638 17752 57690
rect 17776 57638 17790 57690
rect 17790 57638 17802 57690
rect 17802 57638 17832 57690
rect 17856 57638 17866 57690
rect 17866 57638 17912 57690
rect 17616 57636 17672 57638
rect 17696 57636 17752 57638
rect 17776 57636 17832 57638
rect 17856 57636 17912 57638
rect 17616 56602 17672 56604
rect 17696 56602 17752 56604
rect 17776 56602 17832 56604
rect 17856 56602 17912 56604
rect 17616 56550 17662 56602
rect 17662 56550 17672 56602
rect 17696 56550 17726 56602
rect 17726 56550 17738 56602
rect 17738 56550 17752 56602
rect 17776 56550 17790 56602
rect 17790 56550 17802 56602
rect 17802 56550 17832 56602
rect 17856 56550 17866 56602
rect 17866 56550 17912 56602
rect 17616 56548 17672 56550
rect 17696 56548 17752 56550
rect 17776 56548 17832 56550
rect 17856 56548 17912 56550
rect 17616 55514 17672 55516
rect 17696 55514 17752 55516
rect 17776 55514 17832 55516
rect 17856 55514 17912 55516
rect 17616 55462 17662 55514
rect 17662 55462 17672 55514
rect 17696 55462 17726 55514
rect 17726 55462 17738 55514
rect 17738 55462 17752 55514
rect 17776 55462 17790 55514
rect 17790 55462 17802 55514
rect 17802 55462 17832 55514
rect 17856 55462 17866 55514
rect 17866 55462 17912 55514
rect 17616 55460 17672 55462
rect 17696 55460 17752 55462
rect 17776 55460 17832 55462
rect 17856 55460 17912 55462
rect 17616 54426 17672 54428
rect 17696 54426 17752 54428
rect 17776 54426 17832 54428
rect 17856 54426 17912 54428
rect 17616 54374 17662 54426
rect 17662 54374 17672 54426
rect 17696 54374 17726 54426
rect 17726 54374 17738 54426
rect 17738 54374 17752 54426
rect 17776 54374 17790 54426
rect 17790 54374 17802 54426
rect 17802 54374 17832 54426
rect 17856 54374 17866 54426
rect 17866 54374 17912 54426
rect 17616 54372 17672 54374
rect 17696 54372 17752 54374
rect 17776 54372 17832 54374
rect 17856 54372 17912 54374
rect 17616 53338 17672 53340
rect 17696 53338 17752 53340
rect 17776 53338 17832 53340
rect 17856 53338 17912 53340
rect 17616 53286 17662 53338
rect 17662 53286 17672 53338
rect 17696 53286 17726 53338
rect 17726 53286 17738 53338
rect 17738 53286 17752 53338
rect 17776 53286 17790 53338
rect 17790 53286 17802 53338
rect 17802 53286 17832 53338
rect 17856 53286 17866 53338
rect 17866 53286 17912 53338
rect 17616 53284 17672 53286
rect 17696 53284 17752 53286
rect 17776 53284 17832 53286
rect 17856 53284 17912 53286
rect 17616 52250 17672 52252
rect 17696 52250 17752 52252
rect 17776 52250 17832 52252
rect 17856 52250 17912 52252
rect 17616 52198 17662 52250
rect 17662 52198 17672 52250
rect 17696 52198 17726 52250
rect 17726 52198 17738 52250
rect 17738 52198 17752 52250
rect 17776 52198 17790 52250
rect 17790 52198 17802 52250
rect 17802 52198 17832 52250
rect 17856 52198 17866 52250
rect 17866 52198 17912 52250
rect 17616 52196 17672 52198
rect 17696 52196 17752 52198
rect 17776 52196 17832 52198
rect 17856 52196 17912 52198
rect 17616 51162 17672 51164
rect 17696 51162 17752 51164
rect 17776 51162 17832 51164
rect 17856 51162 17912 51164
rect 17616 51110 17662 51162
rect 17662 51110 17672 51162
rect 17696 51110 17726 51162
rect 17726 51110 17738 51162
rect 17738 51110 17752 51162
rect 17776 51110 17790 51162
rect 17790 51110 17802 51162
rect 17802 51110 17832 51162
rect 17856 51110 17866 51162
rect 17866 51110 17912 51162
rect 17616 51108 17672 51110
rect 17696 51108 17752 51110
rect 17776 51108 17832 51110
rect 17856 51108 17912 51110
rect 16956 48442 17012 48444
rect 17036 48442 17092 48444
rect 17116 48442 17172 48444
rect 17196 48442 17252 48444
rect 16956 48390 17002 48442
rect 17002 48390 17012 48442
rect 17036 48390 17066 48442
rect 17066 48390 17078 48442
rect 17078 48390 17092 48442
rect 17116 48390 17130 48442
rect 17130 48390 17142 48442
rect 17142 48390 17172 48442
rect 17196 48390 17206 48442
rect 17206 48390 17252 48442
rect 16956 48388 17012 48390
rect 17036 48388 17092 48390
rect 17116 48388 17172 48390
rect 17196 48388 17252 48390
rect 16956 47354 17012 47356
rect 17036 47354 17092 47356
rect 17116 47354 17172 47356
rect 17196 47354 17252 47356
rect 16956 47302 17002 47354
rect 17002 47302 17012 47354
rect 17036 47302 17066 47354
rect 17066 47302 17078 47354
rect 17078 47302 17092 47354
rect 17116 47302 17130 47354
rect 17130 47302 17142 47354
rect 17142 47302 17172 47354
rect 17196 47302 17206 47354
rect 17206 47302 17252 47354
rect 16956 47300 17012 47302
rect 17036 47300 17092 47302
rect 17116 47300 17172 47302
rect 17196 47300 17252 47302
rect 16956 46266 17012 46268
rect 17036 46266 17092 46268
rect 17116 46266 17172 46268
rect 17196 46266 17252 46268
rect 16956 46214 17002 46266
rect 17002 46214 17012 46266
rect 17036 46214 17066 46266
rect 17066 46214 17078 46266
rect 17078 46214 17092 46266
rect 17116 46214 17130 46266
rect 17130 46214 17142 46266
rect 17142 46214 17172 46266
rect 17196 46214 17206 46266
rect 17206 46214 17252 46266
rect 16956 46212 17012 46214
rect 17036 46212 17092 46214
rect 17116 46212 17172 46214
rect 17196 46212 17252 46214
rect 16956 45178 17012 45180
rect 17036 45178 17092 45180
rect 17116 45178 17172 45180
rect 17196 45178 17252 45180
rect 16956 45126 17002 45178
rect 17002 45126 17012 45178
rect 17036 45126 17066 45178
rect 17066 45126 17078 45178
rect 17078 45126 17092 45178
rect 17116 45126 17130 45178
rect 17130 45126 17142 45178
rect 17142 45126 17172 45178
rect 17196 45126 17206 45178
rect 17206 45126 17252 45178
rect 16956 45124 17012 45126
rect 17036 45124 17092 45126
rect 17116 45124 17172 45126
rect 17196 45124 17252 45126
rect 16956 44090 17012 44092
rect 17036 44090 17092 44092
rect 17116 44090 17172 44092
rect 17196 44090 17252 44092
rect 16956 44038 17002 44090
rect 17002 44038 17012 44090
rect 17036 44038 17066 44090
rect 17066 44038 17078 44090
rect 17078 44038 17092 44090
rect 17116 44038 17130 44090
rect 17130 44038 17142 44090
rect 17142 44038 17172 44090
rect 17196 44038 17206 44090
rect 17206 44038 17252 44090
rect 16956 44036 17012 44038
rect 17036 44036 17092 44038
rect 17116 44036 17172 44038
rect 17196 44036 17252 44038
rect 16956 43002 17012 43004
rect 17036 43002 17092 43004
rect 17116 43002 17172 43004
rect 17196 43002 17252 43004
rect 16956 42950 17002 43002
rect 17002 42950 17012 43002
rect 17036 42950 17066 43002
rect 17066 42950 17078 43002
rect 17078 42950 17092 43002
rect 17116 42950 17130 43002
rect 17130 42950 17142 43002
rect 17142 42950 17172 43002
rect 17196 42950 17206 43002
rect 17206 42950 17252 43002
rect 16956 42948 17012 42950
rect 17036 42948 17092 42950
rect 17116 42948 17172 42950
rect 17196 42948 17252 42950
rect 16956 41914 17012 41916
rect 17036 41914 17092 41916
rect 17116 41914 17172 41916
rect 17196 41914 17252 41916
rect 16956 41862 17002 41914
rect 17002 41862 17012 41914
rect 17036 41862 17066 41914
rect 17066 41862 17078 41914
rect 17078 41862 17092 41914
rect 17116 41862 17130 41914
rect 17130 41862 17142 41914
rect 17142 41862 17172 41914
rect 17196 41862 17206 41914
rect 17206 41862 17252 41914
rect 16956 41860 17012 41862
rect 17036 41860 17092 41862
rect 17116 41860 17172 41862
rect 17196 41860 17252 41862
rect 16956 40826 17012 40828
rect 17036 40826 17092 40828
rect 17116 40826 17172 40828
rect 17196 40826 17252 40828
rect 16956 40774 17002 40826
rect 17002 40774 17012 40826
rect 17036 40774 17066 40826
rect 17066 40774 17078 40826
rect 17078 40774 17092 40826
rect 17116 40774 17130 40826
rect 17130 40774 17142 40826
rect 17142 40774 17172 40826
rect 17196 40774 17206 40826
rect 17206 40774 17252 40826
rect 16956 40772 17012 40774
rect 17036 40772 17092 40774
rect 17116 40772 17172 40774
rect 17196 40772 17252 40774
rect 16956 39738 17012 39740
rect 17036 39738 17092 39740
rect 17116 39738 17172 39740
rect 17196 39738 17252 39740
rect 16956 39686 17002 39738
rect 17002 39686 17012 39738
rect 17036 39686 17066 39738
rect 17066 39686 17078 39738
rect 17078 39686 17092 39738
rect 17116 39686 17130 39738
rect 17130 39686 17142 39738
rect 17142 39686 17172 39738
rect 17196 39686 17206 39738
rect 17206 39686 17252 39738
rect 16956 39684 17012 39686
rect 17036 39684 17092 39686
rect 17116 39684 17172 39686
rect 17196 39684 17252 39686
rect 16956 38650 17012 38652
rect 17036 38650 17092 38652
rect 17116 38650 17172 38652
rect 17196 38650 17252 38652
rect 16956 38598 17002 38650
rect 17002 38598 17012 38650
rect 17036 38598 17066 38650
rect 17066 38598 17078 38650
rect 17078 38598 17092 38650
rect 17116 38598 17130 38650
rect 17130 38598 17142 38650
rect 17142 38598 17172 38650
rect 17196 38598 17206 38650
rect 17206 38598 17252 38650
rect 16956 38596 17012 38598
rect 17036 38596 17092 38598
rect 17116 38596 17172 38598
rect 17196 38596 17252 38598
rect 16956 37562 17012 37564
rect 17036 37562 17092 37564
rect 17116 37562 17172 37564
rect 17196 37562 17252 37564
rect 16956 37510 17002 37562
rect 17002 37510 17012 37562
rect 17036 37510 17066 37562
rect 17066 37510 17078 37562
rect 17078 37510 17092 37562
rect 17116 37510 17130 37562
rect 17130 37510 17142 37562
rect 17142 37510 17172 37562
rect 17196 37510 17206 37562
rect 17206 37510 17252 37562
rect 16956 37508 17012 37510
rect 17036 37508 17092 37510
rect 17116 37508 17172 37510
rect 17196 37508 17252 37510
rect 16956 36474 17012 36476
rect 17036 36474 17092 36476
rect 17116 36474 17172 36476
rect 17196 36474 17252 36476
rect 16956 36422 17002 36474
rect 17002 36422 17012 36474
rect 17036 36422 17066 36474
rect 17066 36422 17078 36474
rect 17078 36422 17092 36474
rect 17116 36422 17130 36474
rect 17130 36422 17142 36474
rect 17142 36422 17172 36474
rect 17196 36422 17206 36474
rect 17206 36422 17252 36474
rect 16956 36420 17012 36422
rect 17036 36420 17092 36422
rect 17116 36420 17172 36422
rect 17196 36420 17252 36422
rect 16956 35386 17012 35388
rect 17036 35386 17092 35388
rect 17116 35386 17172 35388
rect 17196 35386 17252 35388
rect 16956 35334 17002 35386
rect 17002 35334 17012 35386
rect 17036 35334 17066 35386
rect 17066 35334 17078 35386
rect 17078 35334 17092 35386
rect 17116 35334 17130 35386
rect 17130 35334 17142 35386
rect 17142 35334 17172 35386
rect 17196 35334 17206 35386
rect 17206 35334 17252 35386
rect 16956 35332 17012 35334
rect 17036 35332 17092 35334
rect 17116 35332 17172 35334
rect 17196 35332 17252 35334
rect 16956 34298 17012 34300
rect 17036 34298 17092 34300
rect 17116 34298 17172 34300
rect 17196 34298 17252 34300
rect 16956 34246 17002 34298
rect 17002 34246 17012 34298
rect 17036 34246 17066 34298
rect 17066 34246 17078 34298
rect 17078 34246 17092 34298
rect 17116 34246 17130 34298
rect 17130 34246 17142 34298
rect 17142 34246 17172 34298
rect 17196 34246 17206 34298
rect 17206 34246 17252 34298
rect 16956 34244 17012 34246
rect 17036 34244 17092 34246
rect 17116 34244 17172 34246
rect 17196 34244 17252 34246
rect 17616 50074 17672 50076
rect 17696 50074 17752 50076
rect 17776 50074 17832 50076
rect 17856 50074 17912 50076
rect 17616 50022 17662 50074
rect 17662 50022 17672 50074
rect 17696 50022 17726 50074
rect 17726 50022 17738 50074
rect 17738 50022 17752 50074
rect 17776 50022 17790 50074
rect 17790 50022 17802 50074
rect 17802 50022 17832 50074
rect 17856 50022 17866 50074
rect 17866 50022 17912 50074
rect 17616 50020 17672 50022
rect 17696 50020 17752 50022
rect 17776 50020 17832 50022
rect 17856 50020 17912 50022
rect 17616 48986 17672 48988
rect 17696 48986 17752 48988
rect 17776 48986 17832 48988
rect 17856 48986 17912 48988
rect 17616 48934 17662 48986
rect 17662 48934 17672 48986
rect 17696 48934 17726 48986
rect 17726 48934 17738 48986
rect 17738 48934 17752 48986
rect 17776 48934 17790 48986
rect 17790 48934 17802 48986
rect 17802 48934 17832 48986
rect 17856 48934 17866 48986
rect 17866 48934 17912 48986
rect 17616 48932 17672 48934
rect 17696 48932 17752 48934
rect 17776 48932 17832 48934
rect 17856 48932 17912 48934
rect 17616 47898 17672 47900
rect 17696 47898 17752 47900
rect 17776 47898 17832 47900
rect 17856 47898 17912 47900
rect 17616 47846 17662 47898
rect 17662 47846 17672 47898
rect 17696 47846 17726 47898
rect 17726 47846 17738 47898
rect 17738 47846 17752 47898
rect 17776 47846 17790 47898
rect 17790 47846 17802 47898
rect 17802 47846 17832 47898
rect 17856 47846 17866 47898
rect 17866 47846 17912 47898
rect 17616 47844 17672 47846
rect 17696 47844 17752 47846
rect 17776 47844 17832 47846
rect 17856 47844 17912 47846
rect 17616 46810 17672 46812
rect 17696 46810 17752 46812
rect 17776 46810 17832 46812
rect 17856 46810 17912 46812
rect 17616 46758 17662 46810
rect 17662 46758 17672 46810
rect 17696 46758 17726 46810
rect 17726 46758 17738 46810
rect 17738 46758 17752 46810
rect 17776 46758 17790 46810
rect 17790 46758 17802 46810
rect 17802 46758 17832 46810
rect 17856 46758 17866 46810
rect 17866 46758 17912 46810
rect 17616 46756 17672 46758
rect 17696 46756 17752 46758
rect 17776 46756 17832 46758
rect 17856 46756 17912 46758
rect 17616 45722 17672 45724
rect 17696 45722 17752 45724
rect 17776 45722 17832 45724
rect 17856 45722 17912 45724
rect 17616 45670 17662 45722
rect 17662 45670 17672 45722
rect 17696 45670 17726 45722
rect 17726 45670 17738 45722
rect 17738 45670 17752 45722
rect 17776 45670 17790 45722
rect 17790 45670 17802 45722
rect 17802 45670 17832 45722
rect 17856 45670 17866 45722
rect 17866 45670 17912 45722
rect 17616 45668 17672 45670
rect 17696 45668 17752 45670
rect 17776 45668 17832 45670
rect 17856 45668 17912 45670
rect 17616 44634 17672 44636
rect 17696 44634 17752 44636
rect 17776 44634 17832 44636
rect 17856 44634 17912 44636
rect 17616 44582 17662 44634
rect 17662 44582 17672 44634
rect 17696 44582 17726 44634
rect 17726 44582 17738 44634
rect 17738 44582 17752 44634
rect 17776 44582 17790 44634
rect 17790 44582 17802 44634
rect 17802 44582 17832 44634
rect 17856 44582 17866 44634
rect 17866 44582 17912 44634
rect 17616 44580 17672 44582
rect 17696 44580 17752 44582
rect 17776 44580 17832 44582
rect 17856 44580 17912 44582
rect 17616 43546 17672 43548
rect 17696 43546 17752 43548
rect 17776 43546 17832 43548
rect 17856 43546 17912 43548
rect 17616 43494 17662 43546
rect 17662 43494 17672 43546
rect 17696 43494 17726 43546
rect 17726 43494 17738 43546
rect 17738 43494 17752 43546
rect 17776 43494 17790 43546
rect 17790 43494 17802 43546
rect 17802 43494 17832 43546
rect 17856 43494 17866 43546
rect 17866 43494 17912 43546
rect 17616 43492 17672 43494
rect 17696 43492 17752 43494
rect 17776 43492 17832 43494
rect 17856 43492 17912 43494
rect 17616 42458 17672 42460
rect 17696 42458 17752 42460
rect 17776 42458 17832 42460
rect 17856 42458 17912 42460
rect 17616 42406 17662 42458
rect 17662 42406 17672 42458
rect 17696 42406 17726 42458
rect 17726 42406 17738 42458
rect 17738 42406 17752 42458
rect 17776 42406 17790 42458
rect 17790 42406 17802 42458
rect 17802 42406 17832 42458
rect 17856 42406 17866 42458
rect 17866 42406 17912 42458
rect 17616 42404 17672 42406
rect 17696 42404 17752 42406
rect 17776 42404 17832 42406
rect 17856 42404 17912 42406
rect 17616 41370 17672 41372
rect 17696 41370 17752 41372
rect 17776 41370 17832 41372
rect 17856 41370 17912 41372
rect 17616 41318 17662 41370
rect 17662 41318 17672 41370
rect 17696 41318 17726 41370
rect 17726 41318 17738 41370
rect 17738 41318 17752 41370
rect 17776 41318 17790 41370
rect 17790 41318 17802 41370
rect 17802 41318 17832 41370
rect 17856 41318 17866 41370
rect 17866 41318 17912 41370
rect 17616 41316 17672 41318
rect 17696 41316 17752 41318
rect 17776 41316 17832 41318
rect 17856 41316 17912 41318
rect 17616 40282 17672 40284
rect 17696 40282 17752 40284
rect 17776 40282 17832 40284
rect 17856 40282 17912 40284
rect 17616 40230 17662 40282
rect 17662 40230 17672 40282
rect 17696 40230 17726 40282
rect 17726 40230 17738 40282
rect 17738 40230 17752 40282
rect 17776 40230 17790 40282
rect 17790 40230 17802 40282
rect 17802 40230 17832 40282
rect 17856 40230 17866 40282
rect 17866 40230 17912 40282
rect 17616 40228 17672 40230
rect 17696 40228 17752 40230
rect 17776 40228 17832 40230
rect 17856 40228 17912 40230
rect 17616 39194 17672 39196
rect 17696 39194 17752 39196
rect 17776 39194 17832 39196
rect 17856 39194 17912 39196
rect 17616 39142 17662 39194
rect 17662 39142 17672 39194
rect 17696 39142 17726 39194
rect 17726 39142 17738 39194
rect 17738 39142 17752 39194
rect 17776 39142 17790 39194
rect 17790 39142 17802 39194
rect 17802 39142 17832 39194
rect 17856 39142 17866 39194
rect 17866 39142 17912 39194
rect 17616 39140 17672 39142
rect 17696 39140 17752 39142
rect 17776 39140 17832 39142
rect 17856 39140 17912 39142
rect 17616 38106 17672 38108
rect 17696 38106 17752 38108
rect 17776 38106 17832 38108
rect 17856 38106 17912 38108
rect 17616 38054 17662 38106
rect 17662 38054 17672 38106
rect 17696 38054 17726 38106
rect 17726 38054 17738 38106
rect 17738 38054 17752 38106
rect 17776 38054 17790 38106
rect 17790 38054 17802 38106
rect 17802 38054 17832 38106
rect 17856 38054 17866 38106
rect 17866 38054 17912 38106
rect 17616 38052 17672 38054
rect 17696 38052 17752 38054
rect 17776 38052 17832 38054
rect 17856 38052 17912 38054
rect 17616 37018 17672 37020
rect 17696 37018 17752 37020
rect 17776 37018 17832 37020
rect 17856 37018 17912 37020
rect 17616 36966 17662 37018
rect 17662 36966 17672 37018
rect 17696 36966 17726 37018
rect 17726 36966 17738 37018
rect 17738 36966 17752 37018
rect 17776 36966 17790 37018
rect 17790 36966 17802 37018
rect 17802 36966 17832 37018
rect 17856 36966 17866 37018
rect 17866 36966 17912 37018
rect 17616 36964 17672 36966
rect 17696 36964 17752 36966
rect 17776 36964 17832 36966
rect 17856 36964 17912 36966
rect 17616 35930 17672 35932
rect 17696 35930 17752 35932
rect 17776 35930 17832 35932
rect 17856 35930 17912 35932
rect 17616 35878 17662 35930
rect 17662 35878 17672 35930
rect 17696 35878 17726 35930
rect 17726 35878 17738 35930
rect 17738 35878 17752 35930
rect 17776 35878 17790 35930
rect 17790 35878 17802 35930
rect 17802 35878 17832 35930
rect 17856 35878 17866 35930
rect 17866 35878 17912 35930
rect 17616 35876 17672 35878
rect 17696 35876 17752 35878
rect 17776 35876 17832 35878
rect 17856 35876 17912 35878
rect 17616 34842 17672 34844
rect 17696 34842 17752 34844
rect 17776 34842 17832 34844
rect 17856 34842 17912 34844
rect 17616 34790 17662 34842
rect 17662 34790 17672 34842
rect 17696 34790 17726 34842
rect 17726 34790 17738 34842
rect 17738 34790 17752 34842
rect 17776 34790 17790 34842
rect 17790 34790 17802 34842
rect 17802 34790 17832 34842
rect 17856 34790 17866 34842
rect 17866 34790 17912 34842
rect 17616 34788 17672 34790
rect 17696 34788 17752 34790
rect 17776 34788 17832 34790
rect 17856 34788 17912 34790
rect 17616 33754 17672 33756
rect 17696 33754 17752 33756
rect 17776 33754 17832 33756
rect 17856 33754 17912 33756
rect 17616 33702 17662 33754
rect 17662 33702 17672 33754
rect 17696 33702 17726 33754
rect 17726 33702 17738 33754
rect 17738 33702 17752 33754
rect 17776 33702 17790 33754
rect 17790 33702 17802 33754
rect 17802 33702 17832 33754
rect 17856 33702 17866 33754
rect 17866 33702 17912 33754
rect 17616 33700 17672 33702
rect 17696 33700 17752 33702
rect 17776 33700 17832 33702
rect 17856 33700 17912 33702
rect 16956 33210 17012 33212
rect 17036 33210 17092 33212
rect 17116 33210 17172 33212
rect 17196 33210 17252 33212
rect 16956 33158 17002 33210
rect 17002 33158 17012 33210
rect 17036 33158 17066 33210
rect 17066 33158 17078 33210
rect 17078 33158 17092 33210
rect 17116 33158 17130 33210
rect 17130 33158 17142 33210
rect 17142 33158 17172 33210
rect 17196 33158 17206 33210
rect 17206 33158 17252 33210
rect 16956 33156 17012 33158
rect 17036 33156 17092 33158
rect 17116 33156 17172 33158
rect 17196 33156 17252 33158
rect 16956 32122 17012 32124
rect 17036 32122 17092 32124
rect 17116 32122 17172 32124
rect 17196 32122 17252 32124
rect 16956 32070 17002 32122
rect 17002 32070 17012 32122
rect 17036 32070 17066 32122
rect 17066 32070 17078 32122
rect 17078 32070 17092 32122
rect 17116 32070 17130 32122
rect 17130 32070 17142 32122
rect 17142 32070 17172 32122
rect 17196 32070 17206 32122
rect 17206 32070 17252 32122
rect 16956 32068 17012 32070
rect 17036 32068 17092 32070
rect 17116 32068 17172 32070
rect 17196 32068 17252 32070
rect 16578 26832 16634 26888
rect 16578 13368 16634 13424
rect 16956 31034 17012 31036
rect 17036 31034 17092 31036
rect 17116 31034 17172 31036
rect 17196 31034 17252 31036
rect 16956 30982 17002 31034
rect 17002 30982 17012 31034
rect 17036 30982 17066 31034
rect 17066 30982 17078 31034
rect 17078 30982 17092 31034
rect 17116 30982 17130 31034
rect 17130 30982 17142 31034
rect 17142 30982 17172 31034
rect 17196 30982 17206 31034
rect 17206 30982 17252 31034
rect 16956 30980 17012 30982
rect 17036 30980 17092 30982
rect 17116 30980 17172 30982
rect 17196 30980 17252 30982
rect 16956 29946 17012 29948
rect 17036 29946 17092 29948
rect 17116 29946 17172 29948
rect 17196 29946 17252 29948
rect 16956 29894 17002 29946
rect 17002 29894 17012 29946
rect 17036 29894 17066 29946
rect 17066 29894 17078 29946
rect 17078 29894 17092 29946
rect 17116 29894 17130 29946
rect 17130 29894 17142 29946
rect 17142 29894 17172 29946
rect 17196 29894 17206 29946
rect 17206 29894 17252 29946
rect 16956 29892 17012 29894
rect 17036 29892 17092 29894
rect 17116 29892 17172 29894
rect 17196 29892 17252 29894
rect 16956 28858 17012 28860
rect 17036 28858 17092 28860
rect 17116 28858 17172 28860
rect 17196 28858 17252 28860
rect 16956 28806 17002 28858
rect 17002 28806 17012 28858
rect 17036 28806 17066 28858
rect 17066 28806 17078 28858
rect 17078 28806 17092 28858
rect 17116 28806 17130 28858
rect 17130 28806 17142 28858
rect 17142 28806 17172 28858
rect 17196 28806 17206 28858
rect 17206 28806 17252 28858
rect 16956 28804 17012 28806
rect 17036 28804 17092 28806
rect 17116 28804 17172 28806
rect 17196 28804 17252 28806
rect 16956 27770 17012 27772
rect 17036 27770 17092 27772
rect 17116 27770 17172 27772
rect 17196 27770 17252 27772
rect 16956 27718 17002 27770
rect 17002 27718 17012 27770
rect 17036 27718 17066 27770
rect 17066 27718 17078 27770
rect 17078 27718 17092 27770
rect 17116 27718 17130 27770
rect 17130 27718 17142 27770
rect 17142 27718 17172 27770
rect 17196 27718 17206 27770
rect 17206 27718 17252 27770
rect 16956 27716 17012 27718
rect 17036 27716 17092 27718
rect 17116 27716 17172 27718
rect 17196 27716 17252 27718
rect 17314 26968 17370 27024
rect 16956 26682 17012 26684
rect 17036 26682 17092 26684
rect 17116 26682 17172 26684
rect 17196 26682 17252 26684
rect 16956 26630 17002 26682
rect 17002 26630 17012 26682
rect 17036 26630 17066 26682
rect 17066 26630 17078 26682
rect 17078 26630 17092 26682
rect 17116 26630 17130 26682
rect 17130 26630 17142 26682
rect 17142 26630 17172 26682
rect 17196 26630 17206 26682
rect 17206 26630 17252 26682
rect 16956 26628 17012 26630
rect 17036 26628 17092 26630
rect 17116 26628 17172 26630
rect 17196 26628 17252 26630
rect 16956 25594 17012 25596
rect 17036 25594 17092 25596
rect 17116 25594 17172 25596
rect 17196 25594 17252 25596
rect 16956 25542 17002 25594
rect 17002 25542 17012 25594
rect 17036 25542 17066 25594
rect 17066 25542 17078 25594
rect 17078 25542 17092 25594
rect 17116 25542 17130 25594
rect 17130 25542 17142 25594
rect 17142 25542 17172 25594
rect 17196 25542 17206 25594
rect 17206 25542 17252 25594
rect 16956 25540 17012 25542
rect 17036 25540 17092 25542
rect 17116 25540 17172 25542
rect 17196 25540 17252 25542
rect 17616 32666 17672 32668
rect 17696 32666 17752 32668
rect 17776 32666 17832 32668
rect 17856 32666 17912 32668
rect 17616 32614 17662 32666
rect 17662 32614 17672 32666
rect 17696 32614 17726 32666
rect 17726 32614 17738 32666
rect 17738 32614 17752 32666
rect 17776 32614 17790 32666
rect 17790 32614 17802 32666
rect 17802 32614 17832 32666
rect 17856 32614 17866 32666
rect 17866 32614 17912 32666
rect 17616 32612 17672 32614
rect 17696 32612 17752 32614
rect 17776 32612 17832 32614
rect 17856 32612 17912 32614
rect 17616 31578 17672 31580
rect 17696 31578 17752 31580
rect 17776 31578 17832 31580
rect 17856 31578 17912 31580
rect 17616 31526 17662 31578
rect 17662 31526 17672 31578
rect 17696 31526 17726 31578
rect 17726 31526 17738 31578
rect 17738 31526 17752 31578
rect 17776 31526 17790 31578
rect 17790 31526 17802 31578
rect 17802 31526 17832 31578
rect 17856 31526 17866 31578
rect 17866 31526 17912 31578
rect 17616 31524 17672 31526
rect 17696 31524 17752 31526
rect 17776 31524 17832 31526
rect 17856 31524 17912 31526
rect 17616 30490 17672 30492
rect 17696 30490 17752 30492
rect 17776 30490 17832 30492
rect 17856 30490 17912 30492
rect 17616 30438 17662 30490
rect 17662 30438 17672 30490
rect 17696 30438 17726 30490
rect 17726 30438 17738 30490
rect 17738 30438 17752 30490
rect 17776 30438 17790 30490
rect 17790 30438 17802 30490
rect 17802 30438 17832 30490
rect 17856 30438 17866 30490
rect 17866 30438 17912 30490
rect 17616 30436 17672 30438
rect 17696 30436 17752 30438
rect 17776 30436 17832 30438
rect 17856 30436 17912 30438
rect 17616 29402 17672 29404
rect 17696 29402 17752 29404
rect 17776 29402 17832 29404
rect 17856 29402 17912 29404
rect 17616 29350 17662 29402
rect 17662 29350 17672 29402
rect 17696 29350 17726 29402
rect 17726 29350 17738 29402
rect 17738 29350 17752 29402
rect 17776 29350 17790 29402
rect 17790 29350 17802 29402
rect 17802 29350 17832 29402
rect 17856 29350 17866 29402
rect 17866 29350 17912 29402
rect 17616 29348 17672 29350
rect 17696 29348 17752 29350
rect 17776 29348 17832 29350
rect 17856 29348 17912 29350
rect 17616 28314 17672 28316
rect 17696 28314 17752 28316
rect 17776 28314 17832 28316
rect 17856 28314 17912 28316
rect 17616 28262 17662 28314
rect 17662 28262 17672 28314
rect 17696 28262 17726 28314
rect 17726 28262 17738 28314
rect 17738 28262 17752 28314
rect 17776 28262 17790 28314
rect 17790 28262 17802 28314
rect 17802 28262 17832 28314
rect 17856 28262 17866 28314
rect 17866 28262 17912 28314
rect 17616 28260 17672 28262
rect 17696 28260 17752 28262
rect 17776 28260 17832 28262
rect 17856 28260 17912 28262
rect 17616 27226 17672 27228
rect 17696 27226 17752 27228
rect 17776 27226 17832 27228
rect 17856 27226 17912 27228
rect 17616 27174 17662 27226
rect 17662 27174 17672 27226
rect 17696 27174 17726 27226
rect 17726 27174 17738 27226
rect 17738 27174 17752 27226
rect 17776 27174 17790 27226
rect 17790 27174 17802 27226
rect 17802 27174 17832 27226
rect 17856 27174 17866 27226
rect 17866 27174 17912 27226
rect 17616 27172 17672 27174
rect 17696 27172 17752 27174
rect 17776 27172 17832 27174
rect 17856 27172 17912 27174
rect 17616 26138 17672 26140
rect 17696 26138 17752 26140
rect 17776 26138 17832 26140
rect 17856 26138 17912 26140
rect 17616 26086 17662 26138
rect 17662 26086 17672 26138
rect 17696 26086 17726 26138
rect 17726 26086 17738 26138
rect 17738 26086 17752 26138
rect 17776 26086 17790 26138
rect 17790 26086 17802 26138
rect 17802 26086 17832 26138
rect 17856 26086 17866 26138
rect 17866 26086 17912 26138
rect 17616 26084 17672 26086
rect 17696 26084 17752 26086
rect 17776 26084 17832 26086
rect 17856 26084 17912 26086
rect 16956 24506 17012 24508
rect 17036 24506 17092 24508
rect 17116 24506 17172 24508
rect 17196 24506 17252 24508
rect 16956 24454 17002 24506
rect 17002 24454 17012 24506
rect 17036 24454 17066 24506
rect 17066 24454 17078 24506
rect 17078 24454 17092 24506
rect 17116 24454 17130 24506
rect 17130 24454 17142 24506
rect 17142 24454 17172 24506
rect 17196 24454 17206 24506
rect 17206 24454 17252 24506
rect 16956 24452 17012 24454
rect 17036 24452 17092 24454
rect 17116 24452 17172 24454
rect 17196 24452 17252 24454
rect 16956 23418 17012 23420
rect 17036 23418 17092 23420
rect 17116 23418 17172 23420
rect 17196 23418 17252 23420
rect 16956 23366 17002 23418
rect 17002 23366 17012 23418
rect 17036 23366 17066 23418
rect 17066 23366 17078 23418
rect 17078 23366 17092 23418
rect 17116 23366 17130 23418
rect 17130 23366 17142 23418
rect 17142 23366 17172 23418
rect 17196 23366 17206 23418
rect 17206 23366 17252 23418
rect 16956 23364 17012 23366
rect 17036 23364 17092 23366
rect 17116 23364 17172 23366
rect 17196 23364 17252 23366
rect 16956 22330 17012 22332
rect 17036 22330 17092 22332
rect 17116 22330 17172 22332
rect 17196 22330 17252 22332
rect 16956 22278 17002 22330
rect 17002 22278 17012 22330
rect 17036 22278 17066 22330
rect 17066 22278 17078 22330
rect 17078 22278 17092 22330
rect 17116 22278 17130 22330
rect 17130 22278 17142 22330
rect 17142 22278 17172 22330
rect 17196 22278 17206 22330
rect 17206 22278 17252 22330
rect 16956 22276 17012 22278
rect 17036 22276 17092 22278
rect 17116 22276 17172 22278
rect 17196 22276 17252 22278
rect 16956 21242 17012 21244
rect 17036 21242 17092 21244
rect 17116 21242 17172 21244
rect 17196 21242 17252 21244
rect 16956 21190 17002 21242
rect 17002 21190 17012 21242
rect 17036 21190 17066 21242
rect 17066 21190 17078 21242
rect 17078 21190 17092 21242
rect 17116 21190 17130 21242
rect 17130 21190 17142 21242
rect 17142 21190 17172 21242
rect 17196 21190 17206 21242
rect 17206 21190 17252 21242
rect 16956 21188 17012 21190
rect 17036 21188 17092 21190
rect 17116 21188 17172 21190
rect 17196 21188 17252 21190
rect 16956 20154 17012 20156
rect 17036 20154 17092 20156
rect 17116 20154 17172 20156
rect 17196 20154 17252 20156
rect 16956 20102 17002 20154
rect 17002 20102 17012 20154
rect 17036 20102 17066 20154
rect 17066 20102 17078 20154
rect 17078 20102 17092 20154
rect 17116 20102 17130 20154
rect 17130 20102 17142 20154
rect 17142 20102 17172 20154
rect 17196 20102 17206 20154
rect 17206 20102 17252 20154
rect 16956 20100 17012 20102
rect 17036 20100 17092 20102
rect 17116 20100 17172 20102
rect 17196 20100 17252 20102
rect 16956 19066 17012 19068
rect 17036 19066 17092 19068
rect 17116 19066 17172 19068
rect 17196 19066 17252 19068
rect 16956 19014 17002 19066
rect 17002 19014 17012 19066
rect 17036 19014 17066 19066
rect 17066 19014 17078 19066
rect 17078 19014 17092 19066
rect 17116 19014 17130 19066
rect 17130 19014 17142 19066
rect 17142 19014 17172 19066
rect 17196 19014 17206 19066
rect 17206 19014 17252 19066
rect 16956 19012 17012 19014
rect 17036 19012 17092 19014
rect 17116 19012 17172 19014
rect 17196 19012 17252 19014
rect 16956 17978 17012 17980
rect 17036 17978 17092 17980
rect 17116 17978 17172 17980
rect 17196 17978 17252 17980
rect 16956 17926 17002 17978
rect 17002 17926 17012 17978
rect 17036 17926 17066 17978
rect 17066 17926 17078 17978
rect 17078 17926 17092 17978
rect 17116 17926 17130 17978
rect 17130 17926 17142 17978
rect 17142 17926 17172 17978
rect 17196 17926 17206 17978
rect 17206 17926 17252 17978
rect 16956 17924 17012 17926
rect 17036 17924 17092 17926
rect 17116 17924 17172 17926
rect 17196 17924 17252 17926
rect 16956 16890 17012 16892
rect 17036 16890 17092 16892
rect 17116 16890 17172 16892
rect 17196 16890 17252 16892
rect 16956 16838 17002 16890
rect 17002 16838 17012 16890
rect 17036 16838 17066 16890
rect 17066 16838 17078 16890
rect 17078 16838 17092 16890
rect 17116 16838 17130 16890
rect 17130 16838 17142 16890
rect 17142 16838 17172 16890
rect 17196 16838 17206 16890
rect 17206 16838 17252 16890
rect 16956 16836 17012 16838
rect 17036 16836 17092 16838
rect 17116 16836 17172 16838
rect 17196 16836 17252 16838
rect 16956 15802 17012 15804
rect 17036 15802 17092 15804
rect 17116 15802 17172 15804
rect 17196 15802 17252 15804
rect 16956 15750 17002 15802
rect 17002 15750 17012 15802
rect 17036 15750 17066 15802
rect 17066 15750 17078 15802
rect 17078 15750 17092 15802
rect 17116 15750 17130 15802
rect 17130 15750 17142 15802
rect 17142 15750 17172 15802
rect 17196 15750 17206 15802
rect 17206 15750 17252 15802
rect 16956 15748 17012 15750
rect 17036 15748 17092 15750
rect 17116 15748 17172 15750
rect 17196 15748 17252 15750
rect 16956 14714 17012 14716
rect 17036 14714 17092 14716
rect 17116 14714 17172 14716
rect 17196 14714 17252 14716
rect 16956 14662 17002 14714
rect 17002 14662 17012 14714
rect 17036 14662 17066 14714
rect 17066 14662 17078 14714
rect 17078 14662 17092 14714
rect 17116 14662 17130 14714
rect 17130 14662 17142 14714
rect 17142 14662 17172 14714
rect 17196 14662 17206 14714
rect 17206 14662 17252 14714
rect 16956 14660 17012 14662
rect 17036 14660 17092 14662
rect 17116 14660 17172 14662
rect 17196 14660 17252 14662
rect 16956 13626 17012 13628
rect 17036 13626 17092 13628
rect 17116 13626 17172 13628
rect 17196 13626 17252 13628
rect 16956 13574 17002 13626
rect 17002 13574 17012 13626
rect 17036 13574 17066 13626
rect 17066 13574 17078 13626
rect 17078 13574 17092 13626
rect 17116 13574 17130 13626
rect 17130 13574 17142 13626
rect 17142 13574 17172 13626
rect 17196 13574 17206 13626
rect 17206 13574 17252 13626
rect 16956 13572 17012 13574
rect 17036 13572 17092 13574
rect 17116 13572 17172 13574
rect 17196 13572 17252 13574
rect 16956 12538 17012 12540
rect 17036 12538 17092 12540
rect 17116 12538 17172 12540
rect 17196 12538 17252 12540
rect 16956 12486 17002 12538
rect 17002 12486 17012 12538
rect 17036 12486 17066 12538
rect 17066 12486 17078 12538
rect 17078 12486 17092 12538
rect 17116 12486 17130 12538
rect 17130 12486 17142 12538
rect 17142 12486 17172 12538
rect 17196 12486 17206 12538
rect 17206 12486 17252 12538
rect 16956 12484 17012 12486
rect 17036 12484 17092 12486
rect 17116 12484 17172 12486
rect 17196 12484 17252 12486
rect 16956 11450 17012 11452
rect 17036 11450 17092 11452
rect 17116 11450 17172 11452
rect 17196 11450 17252 11452
rect 16956 11398 17002 11450
rect 17002 11398 17012 11450
rect 17036 11398 17066 11450
rect 17066 11398 17078 11450
rect 17078 11398 17092 11450
rect 17116 11398 17130 11450
rect 17130 11398 17142 11450
rect 17142 11398 17172 11450
rect 17196 11398 17206 11450
rect 17206 11398 17252 11450
rect 16956 11396 17012 11398
rect 17036 11396 17092 11398
rect 17116 11396 17172 11398
rect 17196 11396 17252 11398
rect 16956 10362 17012 10364
rect 17036 10362 17092 10364
rect 17116 10362 17172 10364
rect 17196 10362 17252 10364
rect 16956 10310 17002 10362
rect 17002 10310 17012 10362
rect 17036 10310 17066 10362
rect 17066 10310 17078 10362
rect 17078 10310 17092 10362
rect 17116 10310 17130 10362
rect 17130 10310 17142 10362
rect 17142 10310 17172 10362
rect 17196 10310 17206 10362
rect 17206 10310 17252 10362
rect 16956 10308 17012 10310
rect 17036 10308 17092 10310
rect 17116 10308 17172 10310
rect 17196 10308 17252 10310
rect 16956 9274 17012 9276
rect 17036 9274 17092 9276
rect 17116 9274 17172 9276
rect 17196 9274 17252 9276
rect 16956 9222 17002 9274
rect 17002 9222 17012 9274
rect 17036 9222 17066 9274
rect 17066 9222 17078 9274
rect 17078 9222 17092 9274
rect 17116 9222 17130 9274
rect 17130 9222 17142 9274
rect 17142 9222 17172 9274
rect 17196 9222 17206 9274
rect 17206 9222 17252 9274
rect 16956 9220 17012 9222
rect 17036 9220 17092 9222
rect 17116 9220 17172 9222
rect 17196 9220 17252 9222
rect 16956 8186 17012 8188
rect 17036 8186 17092 8188
rect 17116 8186 17172 8188
rect 17196 8186 17252 8188
rect 16956 8134 17002 8186
rect 17002 8134 17012 8186
rect 17036 8134 17066 8186
rect 17066 8134 17078 8186
rect 17078 8134 17092 8186
rect 17116 8134 17130 8186
rect 17130 8134 17142 8186
rect 17142 8134 17172 8186
rect 17196 8134 17206 8186
rect 17206 8134 17252 8186
rect 16956 8132 17012 8134
rect 17036 8132 17092 8134
rect 17116 8132 17172 8134
rect 17196 8132 17252 8134
rect 16956 7098 17012 7100
rect 17036 7098 17092 7100
rect 17116 7098 17172 7100
rect 17196 7098 17252 7100
rect 16956 7046 17002 7098
rect 17002 7046 17012 7098
rect 17036 7046 17066 7098
rect 17066 7046 17078 7098
rect 17078 7046 17092 7098
rect 17116 7046 17130 7098
rect 17130 7046 17142 7098
rect 17142 7046 17172 7098
rect 17196 7046 17206 7098
rect 17206 7046 17252 7098
rect 16956 7044 17012 7046
rect 17036 7044 17092 7046
rect 17116 7044 17172 7046
rect 17196 7044 17252 7046
rect 16956 6010 17012 6012
rect 17036 6010 17092 6012
rect 17116 6010 17172 6012
rect 17196 6010 17252 6012
rect 16956 5958 17002 6010
rect 17002 5958 17012 6010
rect 17036 5958 17066 6010
rect 17066 5958 17078 6010
rect 17078 5958 17092 6010
rect 17116 5958 17130 6010
rect 17130 5958 17142 6010
rect 17142 5958 17172 6010
rect 17196 5958 17206 6010
rect 17206 5958 17252 6010
rect 16956 5956 17012 5958
rect 17036 5956 17092 5958
rect 17116 5956 17172 5958
rect 17196 5956 17252 5958
rect 16956 4922 17012 4924
rect 17036 4922 17092 4924
rect 17116 4922 17172 4924
rect 17196 4922 17252 4924
rect 16956 4870 17002 4922
rect 17002 4870 17012 4922
rect 17036 4870 17066 4922
rect 17066 4870 17078 4922
rect 17078 4870 17092 4922
rect 17116 4870 17130 4922
rect 17130 4870 17142 4922
rect 17142 4870 17172 4922
rect 17196 4870 17206 4922
rect 17206 4870 17252 4922
rect 16956 4868 17012 4870
rect 17036 4868 17092 4870
rect 17116 4868 17172 4870
rect 17196 4868 17252 4870
rect 16956 3834 17012 3836
rect 17036 3834 17092 3836
rect 17116 3834 17172 3836
rect 17196 3834 17252 3836
rect 16956 3782 17002 3834
rect 17002 3782 17012 3834
rect 17036 3782 17066 3834
rect 17066 3782 17078 3834
rect 17078 3782 17092 3834
rect 17116 3782 17130 3834
rect 17130 3782 17142 3834
rect 17142 3782 17172 3834
rect 17196 3782 17206 3834
rect 17206 3782 17252 3834
rect 16956 3780 17012 3782
rect 17036 3780 17092 3782
rect 17116 3780 17172 3782
rect 17196 3780 17252 3782
rect 17616 25050 17672 25052
rect 17696 25050 17752 25052
rect 17776 25050 17832 25052
rect 17856 25050 17912 25052
rect 17616 24998 17662 25050
rect 17662 24998 17672 25050
rect 17696 24998 17726 25050
rect 17726 24998 17738 25050
rect 17738 24998 17752 25050
rect 17776 24998 17790 25050
rect 17790 24998 17802 25050
rect 17802 24998 17832 25050
rect 17856 24998 17866 25050
rect 17866 24998 17912 25050
rect 17616 24996 17672 24998
rect 17696 24996 17752 24998
rect 17776 24996 17832 24998
rect 17856 24996 17912 24998
rect 17616 23962 17672 23964
rect 17696 23962 17752 23964
rect 17776 23962 17832 23964
rect 17856 23962 17912 23964
rect 17616 23910 17662 23962
rect 17662 23910 17672 23962
rect 17696 23910 17726 23962
rect 17726 23910 17738 23962
rect 17738 23910 17752 23962
rect 17776 23910 17790 23962
rect 17790 23910 17802 23962
rect 17802 23910 17832 23962
rect 17856 23910 17866 23962
rect 17866 23910 17912 23962
rect 17616 23908 17672 23910
rect 17696 23908 17752 23910
rect 17776 23908 17832 23910
rect 17856 23908 17912 23910
rect 17616 22874 17672 22876
rect 17696 22874 17752 22876
rect 17776 22874 17832 22876
rect 17856 22874 17912 22876
rect 17616 22822 17662 22874
rect 17662 22822 17672 22874
rect 17696 22822 17726 22874
rect 17726 22822 17738 22874
rect 17738 22822 17752 22874
rect 17776 22822 17790 22874
rect 17790 22822 17802 22874
rect 17802 22822 17832 22874
rect 17856 22822 17866 22874
rect 17866 22822 17912 22874
rect 17616 22820 17672 22822
rect 17696 22820 17752 22822
rect 17776 22820 17832 22822
rect 17856 22820 17912 22822
rect 17616 21786 17672 21788
rect 17696 21786 17752 21788
rect 17776 21786 17832 21788
rect 17856 21786 17912 21788
rect 17616 21734 17662 21786
rect 17662 21734 17672 21786
rect 17696 21734 17726 21786
rect 17726 21734 17738 21786
rect 17738 21734 17752 21786
rect 17776 21734 17790 21786
rect 17790 21734 17802 21786
rect 17802 21734 17832 21786
rect 17856 21734 17866 21786
rect 17866 21734 17912 21786
rect 17616 21732 17672 21734
rect 17696 21732 17752 21734
rect 17776 21732 17832 21734
rect 17856 21732 17912 21734
rect 17616 20698 17672 20700
rect 17696 20698 17752 20700
rect 17776 20698 17832 20700
rect 17856 20698 17912 20700
rect 17616 20646 17662 20698
rect 17662 20646 17672 20698
rect 17696 20646 17726 20698
rect 17726 20646 17738 20698
rect 17738 20646 17752 20698
rect 17776 20646 17790 20698
rect 17790 20646 17802 20698
rect 17802 20646 17832 20698
rect 17856 20646 17866 20698
rect 17866 20646 17912 20698
rect 17616 20644 17672 20646
rect 17696 20644 17752 20646
rect 17776 20644 17832 20646
rect 17856 20644 17912 20646
rect 17616 19610 17672 19612
rect 17696 19610 17752 19612
rect 17776 19610 17832 19612
rect 17856 19610 17912 19612
rect 17616 19558 17662 19610
rect 17662 19558 17672 19610
rect 17696 19558 17726 19610
rect 17726 19558 17738 19610
rect 17738 19558 17752 19610
rect 17776 19558 17790 19610
rect 17790 19558 17802 19610
rect 17802 19558 17832 19610
rect 17856 19558 17866 19610
rect 17866 19558 17912 19610
rect 17616 19556 17672 19558
rect 17696 19556 17752 19558
rect 17776 19556 17832 19558
rect 17856 19556 17912 19558
rect 17616 18522 17672 18524
rect 17696 18522 17752 18524
rect 17776 18522 17832 18524
rect 17856 18522 17912 18524
rect 17616 18470 17662 18522
rect 17662 18470 17672 18522
rect 17696 18470 17726 18522
rect 17726 18470 17738 18522
rect 17738 18470 17752 18522
rect 17776 18470 17790 18522
rect 17790 18470 17802 18522
rect 17802 18470 17832 18522
rect 17856 18470 17866 18522
rect 17866 18470 17912 18522
rect 17616 18468 17672 18470
rect 17696 18468 17752 18470
rect 17776 18468 17832 18470
rect 17856 18468 17912 18470
rect 17616 17434 17672 17436
rect 17696 17434 17752 17436
rect 17776 17434 17832 17436
rect 17856 17434 17912 17436
rect 17616 17382 17662 17434
rect 17662 17382 17672 17434
rect 17696 17382 17726 17434
rect 17726 17382 17738 17434
rect 17738 17382 17752 17434
rect 17776 17382 17790 17434
rect 17790 17382 17802 17434
rect 17802 17382 17832 17434
rect 17856 17382 17866 17434
rect 17866 17382 17912 17434
rect 17616 17380 17672 17382
rect 17696 17380 17752 17382
rect 17776 17380 17832 17382
rect 17856 17380 17912 17382
rect 17616 16346 17672 16348
rect 17696 16346 17752 16348
rect 17776 16346 17832 16348
rect 17856 16346 17912 16348
rect 17616 16294 17662 16346
rect 17662 16294 17672 16346
rect 17696 16294 17726 16346
rect 17726 16294 17738 16346
rect 17738 16294 17752 16346
rect 17776 16294 17790 16346
rect 17790 16294 17802 16346
rect 17802 16294 17832 16346
rect 17856 16294 17866 16346
rect 17866 16294 17912 16346
rect 17616 16292 17672 16294
rect 17696 16292 17752 16294
rect 17776 16292 17832 16294
rect 17856 16292 17912 16294
rect 17616 15258 17672 15260
rect 17696 15258 17752 15260
rect 17776 15258 17832 15260
rect 17856 15258 17912 15260
rect 17616 15206 17662 15258
rect 17662 15206 17672 15258
rect 17696 15206 17726 15258
rect 17726 15206 17738 15258
rect 17738 15206 17752 15258
rect 17776 15206 17790 15258
rect 17790 15206 17802 15258
rect 17802 15206 17832 15258
rect 17856 15206 17866 15258
rect 17866 15206 17912 15258
rect 17616 15204 17672 15206
rect 17696 15204 17752 15206
rect 17776 15204 17832 15206
rect 17856 15204 17912 15206
rect 17616 14170 17672 14172
rect 17696 14170 17752 14172
rect 17776 14170 17832 14172
rect 17856 14170 17912 14172
rect 17616 14118 17662 14170
rect 17662 14118 17672 14170
rect 17696 14118 17726 14170
rect 17726 14118 17738 14170
rect 17738 14118 17752 14170
rect 17776 14118 17790 14170
rect 17790 14118 17802 14170
rect 17802 14118 17832 14170
rect 17856 14118 17866 14170
rect 17866 14118 17912 14170
rect 17616 14116 17672 14118
rect 17696 14116 17752 14118
rect 17776 14116 17832 14118
rect 17856 14116 17912 14118
rect 17616 13082 17672 13084
rect 17696 13082 17752 13084
rect 17776 13082 17832 13084
rect 17856 13082 17912 13084
rect 17616 13030 17662 13082
rect 17662 13030 17672 13082
rect 17696 13030 17726 13082
rect 17726 13030 17738 13082
rect 17738 13030 17752 13082
rect 17776 13030 17790 13082
rect 17790 13030 17802 13082
rect 17802 13030 17832 13082
rect 17856 13030 17866 13082
rect 17866 13030 17912 13082
rect 17616 13028 17672 13030
rect 17696 13028 17752 13030
rect 17776 13028 17832 13030
rect 17856 13028 17912 13030
rect 17616 11994 17672 11996
rect 17696 11994 17752 11996
rect 17776 11994 17832 11996
rect 17856 11994 17912 11996
rect 17616 11942 17662 11994
rect 17662 11942 17672 11994
rect 17696 11942 17726 11994
rect 17726 11942 17738 11994
rect 17738 11942 17752 11994
rect 17776 11942 17790 11994
rect 17790 11942 17802 11994
rect 17802 11942 17832 11994
rect 17856 11942 17866 11994
rect 17866 11942 17912 11994
rect 17616 11940 17672 11942
rect 17696 11940 17752 11942
rect 17776 11940 17832 11942
rect 17856 11940 17912 11942
rect 17616 10906 17672 10908
rect 17696 10906 17752 10908
rect 17776 10906 17832 10908
rect 17856 10906 17912 10908
rect 17616 10854 17662 10906
rect 17662 10854 17672 10906
rect 17696 10854 17726 10906
rect 17726 10854 17738 10906
rect 17738 10854 17752 10906
rect 17776 10854 17790 10906
rect 17790 10854 17802 10906
rect 17802 10854 17832 10906
rect 17856 10854 17866 10906
rect 17866 10854 17912 10906
rect 17616 10852 17672 10854
rect 17696 10852 17752 10854
rect 17776 10852 17832 10854
rect 17856 10852 17912 10854
rect 17616 9818 17672 9820
rect 17696 9818 17752 9820
rect 17776 9818 17832 9820
rect 17856 9818 17912 9820
rect 17616 9766 17662 9818
rect 17662 9766 17672 9818
rect 17696 9766 17726 9818
rect 17726 9766 17738 9818
rect 17738 9766 17752 9818
rect 17776 9766 17790 9818
rect 17790 9766 17802 9818
rect 17802 9766 17832 9818
rect 17856 9766 17866 9818
rect 17866 9766 17912 9818
rect 17616 9764 17672 9766
rect 17696 9764 17752 9766
rect 17776 9764 17832 9766
rect 17856 9764 17912 9766
rect 17616 8730 17672 8732
rect 17696 8730 17752 8732
rect 17776 8730 17832 8732
rect 17856 8730 17912 8732
rect 17616 8678 17662 8730
rect 17662 8678 17672 8730
rect 17696 8678 17726 8730
rect 17726 8678 17738 8730
rect 17738 8678 17752 8730
rect 17776 8678 17790 8730
rect 17790 8678 17802 8730
rect 17802 8678 17832 8730
rect 17856 8678 17866 8730
rect 17866 8678 17912 8730
rect 17616 8676 17672 8678
rect 17696 8676 17752 8678
rect 17776 8676 17832 8678
rect 17856 8676 17912 8678
rect 17616 7642 17672 7644
rect 17696 7642 17752 7644
rect 17776 7642 17832 7644
rect 17856 7642 17912 7644
rect 17616 7590 17662 7642
rect 17662 7590 17672 7642
rect 17696 7590 17726 7642
rect 17726 7590 17738 7642
rect 17738 7590 17752 7642
rect 17776 7590 17790 7642
rect 17790 7590 17802 7642
rect 17802 7590 17832 7642
rect 17856 7590 17866 7642
rect 17866 7590 17912 7642
rect 17616 7588 17672 7590
rect 17696 7588 17752 7590
rect 17776 7588 17832 7590
rect 17856 7588 17912 7590
rect 17616 6554 17672 6556
rect 17696 6554 17752 6556
rect 17776 6554 17832 6556
rect 17856 6554 17912 6556
rect 17616 6502 17662 6554
rect 17662 6502 17672 6554
rect 17696 6502 17726 6554
rect 17726 6502 17738 6554
rect 17738 6502 17752 6554
rect 17776 6502 17790 6554
rect 17790 6502 17802 6554
rect 17802 6502 17832 6554
rect 17856 6502 17866 6554
rect 17866 6502 17912 6554
rect 17616 6500 17672 6502
rect 17696 6500 17752 6502
rect 17776 6500 17832 6502
rect 17856 6500 17912 6502
rect 17616 5466 17672 5468
rect 17696 5466 17752 5468
rect 17776 5466 17832 5468
rect 17856 5466 17912 5468
rect 17616 5414 17662 5466
rect 17662 5414 17672 5466
rect 17696 5414 17726 5466
rect 17726 5414 17738 5466
rect 17738 5414 17752 5466
rect 17776 5414 17790 5466
rect 17790 5414 17802 5466
rect 17802 5414 17832 5466
rect 17856 5414 17866 5466
rect 17866 5414 17912 5466
rect 17616 5412 17672 5414
rect 17696 5412 17752 5414
rect 17776 5412 17832 5414
rect 17856 5412 17912 5414
rect 21956 68026 22012 68028
rect 22036 68026 22092 68028
rect 22116 68026 22172 68028
rect 22196 68026 22252 68028
rect 21956 67974 22002 68026
rect 22002 67974 22012 68026
rect 22036 67974 22066 68026
rect 22066 67974 22078 68026
rect 22078 67974 22092 68026
rect 22116 67974 22130 68026
rect 22130 67974 22142 68026
rect 22142 67974 22172 68026
rect 22196 67974 22206 68026
rect 22206 67974 22252 68026
rect 21956 67972 22012 67974
rect 22036 67972 22092 67974
rect 22116 67972 22172 67974
rect 22196 67972 22252 67974
rect 21956 66938 22012 66940
rect 22036 66938 22092 66940
rect 22116 66938 22172 66940
rect 22196 66938 22252 66940
rect 21956 66886 22002 66938
rect 22002 66886 22012 66938
rect 22036 66886 22066 66938
rect 22066 66886 22078 66938
rect 22078 66886 22092 66938
rect 22116 66886 22130 66938
rect 22130 66886 22142 66938
rect 22142 66886 22172 66938
rect 22196 66886 22206 66938
rect 22206 66886 22252 66938
rect 21956 66884 22012 66886
rect 22036 66884 22092 66886
rect 22116 66884 22172 66886
rect 22196 66884 22252 66886
rect 21956 65850 22012 65852
rect 22036 65850 22092 65852
rect 22116 65850 22172 65852
rect 22196 65850 22252 65852
rect 21956 65798 22002 65850
rect 22002 65798 22012 65850
rect 22036 65798 22066 65850
rect 22066 65798 22078 65850
rect 22078 65798 22092 65850
rect 22116 65798 22130 65850
rect 22130 65798 22142 65850
rect 22142 65798 22172 65850
rect 22196 65798 22206 65850
rect 22206 65798 22252 65850
rect 21956 65796 22012 65798
rect 22036 65796 22092 65798
rect 22116 65796 22172 65798
rect 22196 65796 22252 65798
rect 20166 38936 20222 38992
rect 20350 63552 20406 63608
rect 21956 64762 22012 64764
rect 22036 64762 22092 64764
rect 22116 64762 22172 64764
rect 22196 64762 22252 64764
rect 21956 64710 22002 64762
rect 22002 64710 22012 64762
rect 22036 64710 22066 64762
rect 22066 64710 22078 64762
rect 22078 64710 22092 64762
rect 22116 64710 22130 64762
rect 22130 64710 22142 64762
rect 22142 64710 22172 64762
rect 22196 64710 22206 64762
rect 22206 64710 22252 64762
rect 21956 64708 22012 64710
rect 22036 64708 22092 64710
rect 22116 64708 22172 64710
rect 22196 64708 22252 64710
rect 20626 51992 20682 52048
rect 20350 38836 20352 38856
rect 20352 38836 20404 38856
rect 20404 38836 20406 38856
rect 20350 38800 20406 38836
rect 21956 63674 22012 63676
rect 22036 63674 22092 63676
rect 22116 63674 22172 63676
rect 22196 63674 22252 63676
rect 21956 63622 22002 63674
rect 22002 63622 22012 63674
rect 22036 63622 22066 63674
rect 22066 63622 22078 63674
rect 22078 63622 22092 63674
rect 22116 63622 22130 63674
rect 22130 63622 22142 63674
rect 22142 63622 22172 63674
rect 22196 63622 22206 63674
rect 22206 63622 22252 63674
rect 21956 63620 22012 63622
rect 22036 63620 22092 63622
rect 22116 63620 22172 63622
rect 22196 63620 22252 63622
rect 21730 63552 21786 63608
rect 26956 69114 27012 69116
rect 27036 69114 27092 69116
rect 27116 69114 27172 69116
rect 27196 69114 27252 69116
rect 26956 69062 27002 69114
rect 27002 69062 27012 69114
rect 27036 69062 27066 69114
rect 27066 69062 27078 69114
rect 27078 69062 27092 69114
rect 27116 69062 27130 69114
rect 27130 69062 27142 69114
rect 27142 69062 27172 69114
rect 27196 69062 27206 69114
rect 27206 69062 27252 69114
rect 26956 69060 27012 69062
rect 27036 69060 27092 69062
rect 27116 69060 27172 69062
rect 27196 69060 27252 69062
rect 31956 69114 32012 69116
rect 32036 69114 32092 69116
rect 32116 69114 32172 69116
rect 32196 69114 32252 69116
rect 31956 69062 32002 69114
rect 32002 69062 32012 69114
rect 32036 69062 32066 69114
rect 32066 69062 32078 69114
rect 32078 69062 32092 69114
rect 32116 69062 32130 69114
rect 32130 69062 32142 69114
rect 32142 69062 32172 69114
rect 32196 69062 32206 69114
rect 32206 69062 32252 69114
rect 31956 69060 32012 69062
rect 32036 69060 32092 69062
rect 32116 69060 32172 69062
rect 32196 69060 32252 69062
rect 22616 68570 22672 68572
rect 22696 68570 22752 68572
rect 22776 68570 22832 68572
rect 22856 68570 22912 68572
rect 22616 68518 22662 68570
rect 22662 68518 22672 68570
rect 22696 68518 22726 68570
rect 22726 68518 22738 68570
rect 22738 68518 22752 68570
rect 22776 68518 22790 68570
rect 22790 68518 22802 68570
rect 22802 68518 22832 68570
rect 22856 68518 22866 68570
rect 22866 68518 22912 68570
rect 22616 68516 22672 68518
rect 22696 68516 22752 68518
rect 22776 68516 22832 68518
rect 22856 68516 22912 68518
rect 27616 68570 27672 68572
rect 27696 68570 27752 68572
rect 27776 68570 27832 68572
rect 27856 68570 27912 68572
rect 27616 68518 27662 68570
rect 27662 68518 27672 68570
rect 27696 68518 27726 68570
rect 27726 68518 27738 68570
rect 27738 68518 27752 68570
rect 27776 68518 27790 68570
rect 27790 68518 27802 68570
rect 27802 68518 27832 68570
rect 27856 68518 27866 68570
rect 27866 68518 27912 68570
rect 27616 68516 27672 68518
rect 27696 68516 27752 68518
rect 27776 68516 27832 68518
rect 27856 68516 27912 68518
rect 22616 67482 22672 67484
rect 22696 67482 22752 67484
rect 22776 67482 22832 67484
rect 22856 67482 22912 67484
rect 22616 67430 22662 67482
rect 22662 67430 22672 67482
rect 22696 67430 22726 67482
rect 22726 67430 22738 67482
rect 22738 67430 22752 67482
rect 22776 67430 22790 67482
rect 22790 67430 22802 67482
rect 22802 67430 22832 67482
rect 22856 67430 22866 67482
rect 22866 67430 22912 67482
rect 22616 67428 22672 67430
rect 22696 67428 22752 67430
rect 22776 67428 22832 67430
rect 22856 67428 22912 67430
rect 22616 66394 22672 66396
rect 22696 66394 22752 66396
rect 22776 66394 22832 66396
rect 22856 66394 22912 66396
rect 22616 66342 22662 66394
rect 22662 66342 22672 66394
rect 22696 66342 22726 66394
rect 22726 66342 22738 66394
rect 22738 66342 22752 66394
rect 22776 66342 22790 66394
rect 22790 66342 22802 66394
rect 22802 66342 22832 66394
rect 22856 66342 22866 66394
rect 22866 66342 22912 66394
rect 22616 66340 22672 66342
rect 22696 66340 22752 66342
rect 22776 66340 22832 66342
rect 22856 66340 22912 66342
rect 22616 65306 22672 65308
rect 22696 65306 22752 65308
rect 22776 65306 22832 65308
rect 22856 65306 22912 65308
rect 22616 65254 22662 65306
rect 22662 65254 22672 65306
rect 22696 65254 22726 65306
rect 22726 65254 22738 65306
rect 22738 65254 22752 65306
rect 22776 65254 22790 65306
rect 22790 65254 22802 65306
rect 22802 65254 22832 65306
rect 22856 65254 22866 65306
rect 22866 65254 22912 65306
rect 22616 65252 22672 65254
rect 22696 65252 22752 65254
rect 22776 65252 22832 65254
rect 22856 65252 22912 65254
rect 22616 64218 22672 64220
rect 22696 64218 22752 64220
rect 22776 64218 22832 64220
rect 22856 64218 22912 64220
rect 22616 64166 22662 64218
rect 22662 64166 22672 64218
rect 22696 64166 22726 64218
rect 22726 64166 22738 64218
rect 22738 64166 22752 64218
rect 22776 64166 22790 64218
rect 22790 64166 22802 64218
rect 22802 64166 22832 64218
rect 22856 64166 22866 64218
rect 22866 64166 22912 64218
rect 22616 64164 22672 64166
rect 22696 64164 22752 64166
rect 22776 64164 22832 64166
rect 22856 64164 22912 64166
rect 21956 62586 22012 62588
rect 22036 62586 22092 62588
rect 22116 62586 22172 62588
rect 22196 62586 22252 62588
rect 21956 62534 22002 62586
rect 22002 62534 22012 62586
rect 22036 62534 22066 62586
rect 22066 62534 22078 62586
rect 22078 62534 22092 62586
rect 22116 62534 22130 62586
rect 22130 62534 22142 62586
rect 22142 62534 22172 62586
rect 22196 62534 22206 62586
rect 22206 62534 22252 62586
rect 21956 62532 22012 62534
rect 22036 62532 22092 62534
rect 22116 62532 22172 62534
rect 22196 62532 22252 62534
rect 21956 61498 22012 61500
rect 22036 61498 22092 61500
rect 22116 61498 22172 61500
rect 22196 61498 22252 61500
rect 21956 61446 22002 61498
rect 22002 61446 22012 61498
rect 22036 61446 22066 61498
rect 22066 61446 22078 61498
rect 22078 61446 22092 61498
rect 22116 61446 22130 61498
rect 22130 61446 22142 61498
rect 22142 61446 22172 61498
rect 22196 61446 22206 61498
rect 22206 61446 22252 61498
rect 21956 61444 22012 61446
rect 22036 61444 22092 61446
rect 22116 61444 22172 61446
rect 22196 61444 22252 61446
rect 21956 60410 22012 60412
rect 22036 60410 22092 60412
rect 22116 60410 22172 60412
rect 22196 60410 22252 60412
rect 21956 60358 22002 60410
rect 22002 60358 22012 60410
rect 22036 60358 22066 60410
rect 22066 60358 22078 60410
rect 22078 60358 22092 60410
rect 22116 60358 22130 60410
rect 22130 60358 22142 60410
rect 22142 60358 22172 60410
rect 22196 60358 22206 60410
rect 22206 60358 22252 60410
rect 21956 60356 22012 60358
rect 22036 60356 22092 60358
rect 22116 60356 22172 60358
rect 22196 60356 22252 60358
rect 22098 59472 22154 59528
rect 21956 59322 22012 59324
rect 22036 59322 22092 59324
rect 22116 59322 22172 59324
rect 22196 59322 22252 59324
rect 21956 59270 22002 59322
rect 22002 59270 22012 59322
rect 22036 59270 22066 59322
rect 22066 59270 22078 59322
rect 22078 59270 22092 59322
rect 22116 59270 22130 59322
rect 22130 59270 22142 59322
rect 22142 59270 22172 59322
rect 22196 59270 22206 59322
rect 22206 59270 22252 59322
rect 21956 59268 22012 59270
rect 22036 59268 22092 59270
rect 22116 59268 22172 59270
rect 22196 59268 22252 59270
rect 22616 63130 22672 63132
rect 22696 63130 22752 63132
rect 22776 63130 22832 63132
rect 22856 63130 22912 63132
rect 22616 63078 22662 63130
rect 22662 63078 22672 63130
rect 22696 63078 22726 63130
rect 22726 63078 22738 63130
rect 22738 63078 22752 63130
rect 22776 63078 22790 63130
rect 22790 63078 22802 63130
rect 22802 63078 22832 63130
rect 22856 63078 22866 63130
rect 22866 63078 22912 63130
rect 22616 63076 22672 63078
rect 22696 63076 22752 63078
rect 22776 63076 22832 63078
rect 22856 63076 22912 63078
rect 22616 62042 22672 62044
rect 22696 62042 22752 62044
rect 22776 62042 22832 62044
rect 22856 62042 22912 62044
rect 22616 61990 22662 62042
rect 22662 61990 22672 62042
rect 22696 61990 22726 62042
rect 22726 61990 22738 62042
rect 22738 61990 22752 62042
rect 22776 61990 22790 62042
rect 22790 61990 22802 62042
rect 22802 61990 22832 62042
rect 22856 61990 22866 62042
rect 22866 61990 22912 62042
rect 22616 61988 22672 61990
rect 22696 61988 22752 61990
rect 22776 61988 22832 61990
rect 22856 61988 22912 61990
rect 22616 60954 22672 60956
rect 22696 60954 22752 60956
rect 22776 60954 22832 60956
rect 22856 60954 22912 60956
rect 22616 60902 22662 60954
rect 22662 60902 22672 60954
rect 22696 60902 22726 60954
rect 22726 60902 22738 60954
rect 22738 60902 22752 60954
rect 22776 60902 22790 60954
rect 22790 60902 22802 60954
rect 22802 60902 22832 60954
rect 22856 60902 22866 60954
rect 22866 60902 22912 60954
rect 22616 60900 22672 60902
rect 22696 60900 22752 60902
rect 22776 60900 22832 60902
rect 22856 60900 22912 60902
rect 21956 58234 22012 58236
rect 22036 58234 22092 58236
rect 22116 58234 22172 58236
rect 22196 58234 22252 58236
rect 21956 58182 22002 58234
rect 22002 58182 22012 58234
rect 22036 58182 22066 58234
rect 22066 58182 22078 58234
rect 22078 58182 22092 58234
rect 22116 58182 22130 58234
rect 22130 58182 22142 58234
rect 22142 58182 22172 58234
rect 22196 58182 22206 58234
rect 22206 58182 22252 58234
rect 21956 58180 22012 58182
rect 22036 58180 22092 58182
rect 22116 58180 22172 58182
rect 22196 58180 22252 58182
rect 21956 57146 22012 57148
rect 22036 57146 22092 57148
rect 22116 57146 22172 57148
rect 22196 57146 22252 57148
rect 21956 57094 22002 57146
rect 22002 57094 22012 57146
rect 22036 57094 22066 57146
rect 22066 57094 22078 57146
rect 22078 57094 22092 57146
rect 22116 57094 22130 57146
rect 22130 57094 22142 57146
rect 22142 57094 22172 57146
rect 22196 57094 22206 57146
rect 22206 57094 22252 57146
rect 21956 57092 22012 57094
rect 22036 57092 22092 57094
rect 22116 57092 22172 57094
rect 22196 57092 22252 57094
rect 21956 56058 22012 56060
rect 22036 56058 22092 56060
rect 22116 56058 22172 56060
rect 22196 56058 22252 56060
rect 21956 56006 22002 56058
rect 22002 56006 22012 56058
rect 22036 56006 22066 56058
rect 22066 56006 22078 56058
rect 22078 56006 22092 56058
rect 22116 56006 22130 56058
rect 22130 56006 22142 56058
rect 22142 56006 22172 56058
rect 22196 56006 22206 56058
rect 22206 56006 22252 56058
rect 21956 56004 22012 56006
rect 22036 56004 22092 56006
rect 22116 56004 22172 56006
rect 22196 56004 22252 56006
rect 21956 54970 22012 54972
rect 22036 54970 22092 54972
rect 22116 54970 22172 54972
rect 22196 54970 22252 54972
rect 21956 54918 22002 54970
rect 22002 54918 22012 54970
rect 22036 54918 22066 54970
rect 22066 54918 22078 54970
rect 22078 54918 22092 54970
rect 22116 54918 22130 54970
rect 22130 54918 22142 54970
rect 22142 54918 22172 54970
rect 22196 54918 22206 54970
rect 22206 54918 22252 54970
rect 21956 54916 22012 54918
rect 22036 54916 22092 54918
rect 22116 54916 22172 54918
rect 22196 54916 22252 54918
rect 21454 52028 21456 52048
rect 21456 52028 21508 52048
rect 21508 52028 21510 52048
rect 21454 51992 21510 52028
rect 21956 53882 22012 53884
rect 22036 53882 22092 53884
rect 22116 53882 22172 53884
rect 22196 53882 22252 53884
rect 21956 53830 22002 53882
rect 22002 53830 22012 53882
rect 22036 53830 22066 53882
rect 22066 53830 22078 53882
rect 22078 53830 22092 53882
rect 22116 53830 22130 53882
rect 22130 53830 22142 53882
rect 22142 53830 22172 53882
rect 22196 53830 22206 53882
rect 22206 53830 22252 53882
rect 21956 53828 22012 53830
rect 22036 53828 22092 53830
rect 22116 53828 22172 53830
rect 22196 53828 22252 53830
rect 21956 52794 22012 52796
rect 22036 52794 22092 52796
rect 22116 52794 22172 52796
rect 22196 52794 22252 52796
rect 21956 52742 22002 52794
rect 22002 52742 22012 52794
rect 22036 52742 22066 52794
rect 22066 52742 22078 52794
rect 22078 52742 22092 52794
rect 22116 52742 22130 52794
rect 22130 52742 22142 52794
rect 22142 52742 22172 52794
rect 22196 52742 22206 52794
rect 22206 52742 22252 52794
rect 21956 52740 22012 52742
rect 22036 52740 22092 52742
rect 22116 52740 22172 52742
rect 22196 52740 22252 52742
rect 21956 51706 22012 51708
rect 22036 51706 22092 51708
rect 22116 51706 22172 51708
rect 22196 51706 22252 51708
rect 21956 51654 22002 51706
rect 22002 51654 22012 51706
rect 22036 51654 22066 51706
rect 22066 51654 22078 51706
rect 22078 51654 22092 51706
rect 22116 51654 22130 51706
rect 22130 51654 22142 51706
rect 22142 51654 22172 51706
rect 22196 51654 22206 51706
rect 22206 51654 22252 51706
rect 21956 51652 22012 51654
rect 22036 51652 22092 51654
rect 22116 51652 22172 51654
rect 22196 51652 22252 51654
rect 21956 50618 22012 50620
rect 22036 50618 22092 50620
rect 22116 50618 22172 50620
rect 22196 50618 22252 50620
rect 21956 50566 22002 50618
rect 22002 50566 22012 50618
rect 22036 50566 22066 50618
rect 22066 50566 22078 50618
rect 22078 50566 22092 50618
rect 22116 50566 22130 50618
rect 22130 50566 22142 50618
rect 22142 50566 22172 50618
rect 22196 50566 22206 50618
rect 22206 50566 22252 50618
rect 21956 50564 22012 50566
rect 22036 50564 22092 50566
rect 22116 50564 22172 50566
rect 22196 50564 22252 50566
rect 21956 49530 22012 49532
rect 22036 49530 22092 49532
rect 22116 49530 22172 49532
rect 22196 49530 22252 49532
rect 21956 49478 22002 49530
rect 22002 49478 22012 49530
rect 22036 49478 22066 49530
rect 22066 49478 22078 49530
rect 22078 49478 22092 49530
rect 22116 49478 22130 49530
rect 22130 49478 22142 49530
rect 22142 49478 22172 49530
rect 22196 49478 22206 49530
rect 22206 49478 22252 49530
rect 21956 49476 22012 49478
rect 22036 49476 22092 49478
rect 22116 49476 22172 49478
rect 22196 49476 22252 49478
rect 21956 48442 22012 48444
rect 22036 48442 22092 48444
rect 22116 48442 22172 48444
rect 22196 48442 22252 48444
rect 21956 48390 22002 48442
rect 22002 48390 22012 48442
rect 22036 48390 22066 48442
rect 22066 48390 22078 48442
rect 22078 48390 22092 48442
rect 22116 48390 22130 48442
rect 22130 48390 22142 48442
rect 22142 48390 22172 48442
rect 22196 48390 22206 48442
rect 22206 48390 22252 48442
rect 21956 48388 22012 48390
rect 22036 48388 22092 48390
rect 22116 48388 22172 48390
rect 22196 48388 22252 48390
rect 21956 47354 22012 47356
rect 22036 47354 22092 47356
rect 22116 47354 22172 47356
rect 22196 47354 22252 47356
rect 21956 47302 22002 47354
rect 22002 47302 22012 47354
rect 22036 47302 22066 47354
rect 22066 47302 22078 47354
rect 22078 47302 22092 47354
rect 22116 47302 22130 47354
rect 22130 47302 22142 47354
rect 22142 47302 22172 47354
rect 22196 47302 22206 47354
rect 22206 47302 22252 47354
rect 21956 47300 22012 47302
rect 22036 47300 22092 47302
rect 22116 47300 22172 47302
rect 22196 47300 22252 47302
rect 21956 46266 22012 46268
rect 22036 46266 22092 46268
rect 22116 46266 22172 46268
rect 22196 46266 22252 46268
rect 21956 46214 22002 46266
rect 22002 46214 22012 46266
rect 22036 46214 22066 46266
rect 22066 46214 22078 46266
rect 22078 46214 22092 46266
rect 22116 46214 22130 46266
rect 22130 46214 22142 46266
rect 22142 46214 22172 46266
rect 22196 46214 22206 46266
rect 22206 46214 22252 46266
rect 21956 46212 22012 46214
rect 22036 46212 22092 46214
rect 22116 46212 22172 46214
rect 22196 46212 22252 46214
rect 21956 45178 22012 45180
rect 22036 45178 22092 45180
rect 22116 45178 22172 45180
rect 22196 45178 22252 45180
rect 21956 45126 22002 45178
rect 22002 45126 22012 45178
rect 22036 45126 22066 45178
rect 22066 45126 22078 45178
rect 22078 45126 22092 45178
rect 22116 45126 22130 45178
rect 22130 45126 22142 45178
rect 22142 45126 22172 45178
rect 22196 45126 22206 45178
rect 22206 45126 22252 45178
rect 21956 45124 22012 45126
rect 22036 45124 22092 45126
rect 22116 45124 22172 45126
rect 22196 45124 22252 45126
rect 21956 44090 22012 44092
rect 22036 44090 22092 44092
rect 22116 44090 22172 44092
rect 22196 44090 22252 44092
rect 21956 44038 22002 44090
rect 22002 44038 22012 44090
rect 22036 44038 22066 44090
rect 22066 44038 22078 44090
rect 22078 44038 22092 44090
rect 22116 44038 22130 44090
rect 22130 44038 22142 44090
rect 22142 44038 22172 44090
rect 22196 44038 22206 44090
rect 22206 44038 22252 44090
rect 21956 44036 22012 44038
rect 22036 44036 22092 44038
rect 22116 44036 22172 44038
rect 22196 44036 22252 44038
rect 21956 43002 22012 43004
rect 22036 43002 22092 43004
rect 22116 43002 22172 43004
rect 22196 43002 22252 43004
rect 21956 42950 22002 43002
rect 22002 42950 22012 43002
rect 22036 42950 22066 43002
rect 22066 42950 22078 43002
rect 22078 42950 22092 43002
rect 22116 42950 22130 43002
rect 22130 42950 22142 43002
rect 22142 42950 22172 43002
rect 22196 42950 22206 43002
rect 22206 42950 22252 43002
rect 21956 42948 22012 42950
rect 22036 42948 22092 42950
rect 22116 42948 22172 42950
rect 22196 42948 22252 42950
rect 22098 42744 22154 42800
rect 22616 59866 22672 59868
rect 22696 59866 22752 59868
rect 22776 59866 22832 59868
rect 22856 59866 22912 59868
rect 22616 59814 22662 59866
rect 22662 59814 22672 59866
rect 22696 59814 22726 59866
rect 22726 59814 22738 59866
rect 22738 59814 22752 59866
rect 22776 59814 22790 59866
rect 22790 59814 22802 59866
rect 22802 59814 22832 59866
rect 22856 59814 22866 59866
rect 22866 59814 22912 59866
rect 22616 59812 22672 59814
rect 22696 59812 22752 59814
rect 22776 59812 22832 59814
rect 22856 59812 22912 59814
rect 22616 58778 22672 58780
rect 22696 58778 22752 58780
rect 22776 58778 22832 58780
rect 22856 58778 22912 58780
rect 22616 58726 22662 58778
rect 22662 58726 22672 58778
rect 22696 58726 22726 58778
rect 22726 58726 22738 58778
rect 22738 58726 22752 58778
rect 22776 58726 22790 58778
rect 22790 58726 22802 58778
rect 22802 58726 22832 58778
rect 22856 58726 22866 58778
rect 22866 58726 22912 58778
rect 22616 58724 22672 58726
rect 22696 58724 22752 58726
rect 22776 58724 22832 58726
rect 22856 58724 22912 58726
rect 22616 57690 22672 57692
rect 22696 57690 22752 57692
rect 22776 57690 22832 57692
rect 22856 57690 22912 57692
rect 22616 57638 22662 57690
rect 22662 57638 22672 57690
rect 22696 57638 22726 57690
rect 22726 57638 22738 57690
rect 22738 57638 22752 57690
rect 22776 57638 22790 57690
rect 22790 57638 22802 57690
rect 22802 57638 22832 57690
rect 22856 57638 22866 57690
rect 22866 57638 22912 57690
rect 22616 57636 22672 57638
rect 22696 57636 22752 57638
rect 22776 57636 22832 57638
rect 22856 57636 22912 57638
rect 22616 56602 22672 56604
rect 22696 56602 22752 56604
rect 22776 56602 22832 56604
rect 22856 56602 22912 56604
rect 22616 56550 22662 56602
rect 22662 56550 22672 56602
rect 22696 56550 22726 56602
rect 22726 56550 22738 56602
rect 22738 56550 22752 56602
rect 22776 56550 22790 56602
rect 22790 56550 22802 56602
rect 22802 56550 22832 56602
rect 22856 56550 22866 56602
rect 22866 56550 22912 56602
rect 22616 56548 22672 56550
rect 22696 56548 22752 56550
rect 22776 56548 22832 56550
rect 22856 56548 22912 56550
rect 22616 55514 22672 55516
rect 22696 55514 22752 55516
rect 22776 55514 22832 55516
rect 22856 55514 22912 55516
rect 22616 55462 22662 55514
rect 22662 55462 22672 55514
rect 22696 55462 22726 55514
rect 22726 55462 22738 55514
rect 22738 55462 22752 55514
rect 22776 55462 22790 55514
rect 22790 55462 22802 55514
rect 22802 55462 22832 55514
rect 22856 55462 22866 55514
rect 22866 55462 22912 55514
rect 22616 55460 22672 55462
rect 22696 55460 22752 55462
rect 22776 55460 22832 55462
rect 22856 55460 22912 55462
rect 22616 54426 22672 54428
rect 22696 54426 22752 54428
rect 22776 54426 22832 54428
rect 22856 54426 22912 54428
rect 22616 54374 22662 54426
rect 22662 54374 22672 54426
rect 22696 54374 22726 54426
rect 22726 54374 22738 54426
rect 22738 54374 22752 54426
rect 22776 54374 22790 54426
rect 22790 54374 22802 54426
rect 22802 54374 22832 54426
rect 22856 54374 22866 54426
rect 22866 54374 22912 54426
rect 22616 54372 22672 54374
rect 22696 54372 22752 54374
rect 22776 54372 22832 54374
rect 22856 54372 22912 54374
rect 22616 53338 22672 53340
rect 22696 53338 22752 53340
rect 22776 53338 22832 53340
rect 22856 53338 22912 53340
rect 22616 53286 22662 53338
rect 22662 53286 22672 53338
rect 22696 53286 22726 53338
rect 22726 53286 22738 53338
rect 22738 53286 22752 53338
rect 22776 53286 22790 53338
rect 22790 53286 22802 53338
rect 22802 53286 22832 53338
rect 22856 53286 22866 53338
rect 22866 53286 22912 53338
rect 22616 53284 22672 53286
rect 22696 53284 22752 53286
rect 22776 53284 22832 53286
rect 22856 53284 22912 53286
rect 22616 52250 22672 52252
rect 22696 52250 22752 52252
rect 22776 52250 22832 52252
rect 22856 52250 22912 52252
rect 22616 52198 22662 52250
rect 22662 52198 22672 52250
rect 22696 52198 22726 52250
rect 22726 52198 22738 52250
rect 22738 52198 22752 52250
rect 22776 52198 22790 52250
rect 22790 52198 22802 52250
rect 22802 52198 22832 52250
rect 22856 52198 22866 52250
rect 22866 52198 22912 52250
rect 22616 52196 22672 52198
rect 22696 52196 22752 52198
rect 22776 52196 22832 52198
rect 22856 52196 22912 52198
rect 22616 51162 22672 51164
rect 22696 51162 22752 51164
rect 22776 51162 22832 51164
rect 22856 51162 22912 51164
rect 22616 51110 22662 51162
rect 22662 51110 22672 51162
rect 22696 51110 22726 51162
rect 22726 51110 22738 51162
rect 22738 51110 22752 51162
rect 22776 51110 22790 51162
rect 22790 51110 22802 51162
rect 22802 51110 22832 51162
rect 22856 51110 22866 51162
rect 22866 51110 22912 51162
rect 22616 51108 22672 51110
rect 22696 51108 22752 51110
rect 22776 51108 22832 51110
rect 22856 51108 22912 51110
rect 22616 50074 22672 50076
rect 22696 50074 22752 50076
rect 22776 50074 22832 50076
rect 22856 50074 22912 50076
rect 22616 50022 22662 50074
rect 22662 50022 22672 50074
rect 22696 50022 22726 50074
rect 22726 50022 22738 50074
rect 22738 50022 22752 50074
rect 22776 50022 22790 50074
rect 22790 50022 22802 50074
rect 22802 50022 22832 50074
rect 22856 50022 22866 50074
rect 22866 50022 22912 50074
rect 22616 50020 22672 50022
rect 22696 50020 22752 50022
rect 22776 50020 22832 50022
rect 22856 50020 22912 50022
rect 22616 48986 22672 48988
rect 22696 48986 22752 48988
rect 22776 48986 22832 48988
rect 22856 48986 22912 48988
rect 22616 48934 22662 48986
rect 22662 48934 22672 48986
rect 22696 48934 22726 48986
rect 22726 48934 22738 48986
rect 22738 48934 22752 48986
rect 22776 48934 22790 48986
rect 22790 48934 22802 48986
rect 22802 48934 22832 48986
rect 22856 48934 22866 48986
rect 22866 48934 22912 48986
rect 22616 48932 22672 48934
rect 22696 48932 22752 48934
rect 22776 48932 22832 48934
rect 22856 48932 22912 48934
rect 22616 47898 22672 47900
rect 22696 47898 22752 47900
rect 22776 47898 22832 47900
rect 22856 47898 22912 47900
rect 22616 47846 22662 47898
rect 22662 47846 22672 47898
rect 22696 47846 22726 47898
rect 22726 47846 22738 47898
rect 22738 47846 22752 47898
rect 22776 47846 22790 47898
rect 22790 47846 22802 47898
rect 22802 47846 22832 47898
rect 22856 47846 22866 47898
rect 22866 47846 22912 47898
rect 22616 47844 22672 47846
rect 22696 47844 22752 47846
rect 22776 47844 22832 47846
rect 22856 47844 22912 47846
rect 22616 46810 22672 46812
rect 22696 46810 22752 46812
rect 22776 46810 22832 46812
rect 22856 46810 22912 46812
rect 22616 46758 22662 46810
rect 22662 46758 22672 46810
rect 22696 46758 22726 46810
rect 22726 46758 22738 46810
rect 22738 46758 22752 46810
rect 22776 46758 22790 46810
rect 22790 46758 22802 46810
rect 22802 46758 22832 46810
rect 22856 46758 22866 46810
rect 22866 46758 22912 46810
rect 22616 46756 22672 46758
rect 22696 46756 22752 46758
rect 22776 46756 22832 46758
rect 22856 46756 22912 46758
rect 22616 45722 22672 45724
rect 22696 45722 22752 45724
rect 22776 45722 22832 45724
rect 22856 45722 22912 45724
rect 22616 45670 22662 45722
rect 22662 45670 22672 45722
rect 22696 45670 22726 45722
rect 22726 45670 22738 45722
rect 22738 45670 22752 45722
rect 22776 45670 22790 45722
rect 22790 45670 22802 45722
rect 22802 45670 22832 45722
rect 22856 45670 22866 45722
rect 22866 45670 22912 45722
rect 22616 45668 22672 45670
rect 22696 45668 22752 45670
rect 22776 45668 22832 45670
rect 22856 45668 22912 45670
rect 22616 44634 22672 44636
rect 22696 44634 22752 44636
rect 22776 44634 22832 44636
rect 22856 44634 22912 44636
rect 22616 44582 22662 44634
rect 22662 44582 22672 44634
rect 22696 44582 22726 44634
rect 22726 44582 22738 44634
rect 22738 44582 22752 44634
rect 22776 44582 22790 44634
rect 22790 44582 22802 44634
rect 22802 44582 22832 44634
rect 22856 44582 22866 44634
rect 22866 44582 22912 44634
rect 22616 44580 22672 44582
rect 22696 44580 22752 44582
rect 22776 44580 22832 44582
rect 22856 44580 22912 44582
rect 22616 43546 22672 43548
rect 22696 43546 22752 43548
rect 22776 43546 22832 43548
rect 22856 43546 22912 43548
rect 22616 43494 22662 43546
rect 22662 43494 22672 43546
rect 22696 43494 22726 43546
rect 22726 43494 22738 43546
rect 22738 43494 22752 43546
rect 22776 43494 22790 43546
rect 22790 43494 22802 43546
rect 22802 43494 22832 43546
rect 22856 43494 22866 43546
rect 22866 43494 22912 43546
rect 22616 43492 22672 43494
rect 22696 43492 22752 43494
rect 22776 43492 22832 43494
rect 22856 43492 22912 43494
rect 22466 42744 22522 42800
rect 21956 41914 22012 41916
rect 22036 41914 22092 41916
rect 22116 41914 22172 41916
rect 22196 41914 22252 41916
rect 21956 41862 22002 41914
rect 22002 41862 22012 41914
rect 22036 41862 22066 41914
rect 22066 41862 22078 41914
rect 22078 41862 22092 41914
rect 22116 41862 22130 41914
rect 22130 41862 22142 41914
rect 22142 41862 22172 41914
rect 22196 41862 22206 41914
rect 22206 41862 22252 41914
rect 21956 41860 22012 41862
rect 22036 41860 22092 41862
rect 22116 41860 22172 41862
rect 22196 41860 22252 41862
rect 21956 40826 22012 40828
rect 22036 40826 22092 40828
rect 22116 40826 22172 40828
rect 22196 40826 22252 40828
rect 21956 40774 22002 40826
rect 22002 40774 22012 40826
rect 22036 40774 22066 40826
rect 22066 40774 22078 40826
rect 22078 40774 22092 40826
rect 22116 40774 22130 40826
rect 22130 40774 22142 40826
rect 22142 40774 22172 40826
rect 22196 40774 22206 40826
rect 22206 40774 22252 40826
rect 21956 40772 22012 40774
rect 22036 40772 22092 40774
rect 22116 40772 22172 40774
rect 22196 40772 22252 40774
rect 21956 39738 22012 39740
rect 22036 39738 22092 39740
rect 22116 39738 22172 39740
rect 22196 39738 22252 39740
rect 21956 39686 22002 39738
rect 22002 39686 22012 39738
rect 22036 39686 22066 39738
rect 22066 39686 22078 39738
rect 22078 39686 22092 39738
rect 22116 39686 22130 39738
rect 22130 39686 22142 39738
rect 22142 39686 22172 39738
rect 22196 39686 22206 39738
rect 22206 39686 22252 39738
rect 21956 39684 22012 39686
rect 22036 39684 22092 39686
rect 22116 39684 22172 39686
rect 22196 39684 22252 39686
rect 22190 39344 22246 39400
rect 21956 38650 22012 38652
rect 22036 38650 22092 38652
rect 22116 38650 22172 38652
rect 22196 38650 22252 38652
rect 21956 38598 22002 38650
rect 22002 38598 22012 38650
rect 22036 38598 22066 38650
rect 22066 38598 22078 38650
rect 22078 38598 22092 38650
rect 22116 38598 22130 38650
rect 22130 38598 22142 38650
rect 22142 38598 22172 38650
rect 22196 38598 22206 38650
rect 22206 38598 22252 38650
rect 21956 38596 22012 38598
rect 22036 38596 22092 38598
rect 22116 38596 22172 38598
rect 22196 38596 22252 38598
rect 21956 37562 22012 37564
rect 22036 37562 22092 37564
rect 22116 37562 22172 37564
rect 22196 37562 22252 37564
rect 21956 37510 22002 37562
rect 22002 37510 22012 37562
rect 22036 37510 22066 37562
rect 22066 37510 22078 37562
rect 22078 37510 22092 37562
rect 22116 37510 22130 37562
rect 22130 37510 22142 37562
rect 22142 37510 22172 37562
rect 22196 37510 22206 37562
rect 22206 37510 22252 37562
rect 21956 37508 22012 37510
rect 22036 37508 22092 37510
rect 22116 37508 22172 37510
rect 22196 37508 22252 37510
rect 21956 36474 22012 36476
rect 22036 36474 22092 36476
rect 22116 36474 22172 36476
rect 22196 36474 22252 36476
rect 21956 36422 22002 36474
rect 22002 36422 22012 36474
rect 22036 36422 22066 36474
rect 22066 36422 22078 36474
rect 22078 36422 22092 36474
rect 22116 36422 22130 36474
rect 22130 36422 22142 36474
rect 22142 36422 22172 36474
rect 22196 36422 22206 36474
rect 22206 36422 22252 36474
rect 21956 36420 22012 36422
rect 22036 36420 22092 36422
rect 22116 36420 22172 36422
rect 22196 36420 22252 36422
rect 21956 35386 22012 35388
rect 22036 35386 22092 35388
rect 22116 35386 22172 35388
rect 22196 35386 22252 35388
rect 21956 35334 22002 35386
rect 22002 35334 22012 35386
rect 22036 35334 22066 35386
rect 22066 35334 22078 35386
rect 22078 35334 22092 35386
rect 22116 35334 22130 35386
rect 22130 35334 22142 35386
rect 22142 35334 22172 35386
rect 22196 35334 22206 35386
rect 22206 35334 22252 35386
rect 21956 35332 22012 35334
rect 22036 35332 22092 35334
rect 22116 35332 22172 35334
rect 22196 35332 22252 35334
rect 21956 34298 22012 34300
rect 22036 34298 22092 34300
rect 22116 34298 22172 34300
rect 22196 34298 22252 34300
rect 21956 34246 22002 34298
rect 22002 34246 22012 34298
rect 22036 34246 22066 34298
rect 22066 34246 22078 34298
rect 22078 34246 22092 34298
rect 22116 34246 22130 34298
rect 22130 34246 22142 34298
rect 22142 34246 22172 34298
rect 22196 34246 22206 34298
rect 22206 34246 22252 34298
rect 21956 34244 22012 34246
rect 22036 34244 22092 34246
rect 22116 34244 22172 34246
rect 22196 34244 22252 34246
rect 21956 33210 22012 33212
rect 22036 33210 22092 33212
rect 22116 33210 22172 33212
rect 22196 33210 22252 33212
rect 21956 33158 22002 33210
rect 22002 33158 22012 33210
rect 22036 33158 22066 33210
rect 22066 33158 22078 33210
rect 22078 33158 22092 33210
rect 22116 33158 22130 33210
rect 22130 33158 22142 33210
rect 22142 33158 22172 33210
rect 22196 33158 22206 33210
rect 22206 33158 22252 33210
rect 21956 33156 22012 33158
rect 22036 33156 22092 33158
rect 22116 33156 22172 33158
rect 22196 33156 22252 33158
rect 21956 32122 22012 32124
rect 22036 32122 22092 32124
rect 22116 32122 22172 32124
rect 22196 32122 22252 32124
rect 21956 32070 22002 32122
rect 22002 32070 22012 32122
rect 22036 32070 22066 32122
rect 22066 32070 22078 32122
rect 22078 32070 22092 32122
rect 22116 32070 22130 32122
rect 22130 32070 22142 32122
rect 22142 32070 22172 32122
rect 22196 32070 22206 32122
rect 22206 32070 22252 32122
rect 21956 32068 22012 32070
rect 22036 32068 22092 32070
rect 22116 32068 22172 32070
rect 22196 32068 22252 32070
rect 21956 31034 22012 31036
rect 22036 31034 22092 31036
rect 22116 31034 22172 31036
rect 22196 31034 22252 31036
rect 21956 30982 22002 31034
rect 22002 30982 22012 31034
rect 22036 30982 22066 31034
rect 22066 30982 22078 31034
rect 22078 30982 22092 31034
rect 22116 30982 22130 31034
rect 22130 30982 22142 31034
rect 22142 30982 22172 31034
rect 22196 30982 22206 31034
rect 22206 30982 22252 31034
rect 21956 30980 22012 30982
rect 22036 30980 22092 30982
rect 22116 30980 22172 30982
rect 22196 30980 22252 30982
rect 21956 29946 22012 29948
rect 22036 29946 22092 29948
rect 22116 29946 22172 29948
rect 22196 29946 22252 29948
rect 21956 29894 22002 29946
rect 22002 29894 22012 29946
rect 22036 29894 22066 29946
rect 22066 29894 22078 29946
rect 22078 29894 22092 29946
rect 22116 29894 22130 29946
rect 22130 29894 22142 29946
rect 22142 29894 22172 29946
rect 22196 29894 22206 29946
rect 22206 29894 22252 29946
rect 21956 29892 22012 29894
rect 22036 29892 22092 29894
rect 22116 29892 22172 29894
rect 22196 29892 22252 29894
rect 21956 28858 22012 28860
rect 22036 28858 22092 28860
rect 22116 28858 22172 28860
rect 22196 28858 22252 28860
rect 21956 28806 22002 28858
rect 22002 28806 22012 28858
rect 22036 28806 22066 28858
rect 22066 28806 22078 28858
rect 22078 28806 22092 28858
rect 22116 28806 22130 28858
rect 22130 28806 22142 28858
rect 22142 28806 22172 28858
rect 22196 28806 22206 28858
rect 22206 28806 22252 28858
rect 21956 28804 22012 28806
rect 22036 28804 22092 28806
rect 22116 28804 22172 28806
rect 22196 28804 22252 28806
rect 21956 27770 22012 27772
rect 22036 27770 22092 27772
rect 22116 27770 22172 27772
rect 22196 27770 22252 27772
rect 21956 27718 22002 27770
rect 22002 27718 22012 27770
rect 22036 27718 22066 27770
rect 22066 27718 22078 27770
rect 22078 27718 22092 27770
rect 22116 27718 22130 27770
rect 22130 27718 22142 27770
rect 22142 27718 22172 27770
rect 22196 27718 22206 27770
rect 22206 27718 22252 27770
rect 21956 27716 22012 27718
rect 22036 27716 22092 27718
rect 22116 27716 22172 27718
rect 22196 27716 22252 27718
rect 21956 26682 22012 26684
rect 22036 26682 22092 26684
rect 22116 26682 22172 26684
rect 22196 26682 22252 26684
rect 21956 26630 22002 26682
rect 22002 26630 22012 26682
rect 22036 26630 22066 26682
rect 22066 26630 22078 26682
rect 22078 26630 22092 26682
rect 22116 26630 22130 26682
rect 22130 26630 22142 26682
rect 22142 26630 22172 26682
rect 22196 26630 22206 26682
rect 22206 26630 22252 26682
rect 21956 26628 22012 26630
rect 22036 26628 22092 26630
rect 22116 26628 22172 26630
rect 22196 26628 22252 26630
rect 21956 25594 22012 25596
rect 22036 25594 22092 25596
rect 22116 25594 22172 25596
rect 22196 25594 22252 25596
rect 21956 25542 22002 25594
rect 22002 25542 22012 25594
rect 22036 25542 22066 25594
rect 22066 25542 22078 25594
rect 22078 25542 22092 25594
rect 22116 25542 22130 25594
rect 22130 25542 22142 25594
rect 22142 25542 22172 25594
rect 22196 25542 22206 25594
rect 22206 25542 22252 25594
rect 21956 25540 22012 25542
rect 22036 25540 22092 25542
rect 22116 25540 22172 25542
rect 22196 25540 22252 25542
rect 21956 24506 22012 24508
rect 22036 24506 22092 24508
rect 22116 24506 22172 24508
rect 22196 24506 22252 24508
rect 21956 24454 22002 24506
rect 22002 24454 22012 24506
rect 22036 24454 22066 24506
rect 22066 24454 22078 24506
rect 22078 24454 22092 24506
rect 22116 24454 22130 24506
rect 22130 24454 22142 24506
rect 22142 24454 22172 24506
rect 22196 24454 22206 24506
rect 22206 24454 22252 24506
rect 21956 24452 22012 24454
rect 22036 24452 22092 24454
rect 22116 24452 22172 24454
rect 22196 24452 22252 24454
rect 21956 23418 22012 23420
rect 22036 23418 22092 23420
rect 22116 23418 22172 23420
rect 22196 23418 22252 23420
rect 21956 23366 22002 23418
rect 22002 23366 22012 23418
rect 22036 23366 22066 23418
rect 22066 23366 22078 23418
rect 22078 23366 22092 23418
rect 22116 23366 22130 23418
rect 22130 23366 22142 23418
rect 22142 23366 22172 23418
rect 22196 23366 22206 23418
rect 22206 23366 22252 23418
rect 21956 23364 22012 23366
rect 22036 23364 22092 23366
rect 22116 23364 22172 23366
rect 22196 23364 22252 23366
rect 21956 22330 22012 22332
rect 22036 22330 22092 22332
rect 22116 22330 22172 22332
rect 22196 22330 22252 22332
rect 21956 22278 22002 22330
rect 22002 22278 22012 22330
rect 22036 22278 22066 22330
rect 22066 22278 22078 22330
rect 22078 22278 22092 22330
rect 22116 22278 22130 22330
rect 22130 22278 22142 22330
rect 22142 22278 22172 22330
rect 22196 22278 22206 22330
rect 22206 22278 22252 22330
rect 21956 22276 22012 22278
rect 22036 22276 22092 22278
rect 22116 22276 22172 22278
rect 22196 22276 22252 22278
rect 21956 21242 22012 21244
rect 22036 21242 22092 21244
rect 22116 21242 22172 21244
rect 22196 21242 22252 21244
rect 21956 21190 22002 21242
rect 22002 21190 22012 21242
rect 22036 21190 22066 21242
rect 22066 21190 22078 21242
rect 22078 21190 22092 21242
rect 22116 21190 22130 21242
rect 22130 21190 22142 21242
rect 22142 21190 22172 21242
rect 22196 21190 22206 21242
rect 22206 21190 22252 21242
rect 21956 21188 22012 21190
rect 22036 21188 22092 21190
rect 22116 21188 22172 21190
rect 22196 21188 22252 21190
rect 22616 42458 22672 42460
rect 22696 42458 22752 42460
rect 22776 42458 22832 42460
rect 22856 42458 22912 42460
rect 22616 42406 22662 42458
rect 22662 42406 22672 42458
rect 22696 42406 22726 42458
rect 22726 42406 22738 42458
rect 22738 42406 22752 42458
rect 22776 42406 22790 42458
rect 22790 42406 22802 42458
rect 22802 42406 22832 42458
rect 22856 42406 22866 42458
rect 22866 42406 22912 42458
rect 22616 42404 22672 42406
rect 22696 42404 22752 42406
rect 22776 42404 22832 42406
rect 22856 42404 22912 42406
rect 22616 41370 22672 41372
rect 22696 41370 22752 41372
rect 22776 41370 22832 41372
rect 22856 41370 22912 41372
rect 22616 41318 22662 41370
rect 22662 41318 22672 41370
rect 22696 41318 22726 41370
rect 22726 41318 22738 41370
rect 22738 41318 22752 41370
rect 22776 41318 22790 41370
rect 22790 41318 22802 41370
rect 22802 41318 22832 41370
rect 22856 41318 22866 41370
rect 22866 41318 22912 41370
rect 22616 41316 22672 41318
rect 22696 41316 22752 41318
rect 22776 41316 22832 41318
rect 22856 41316 22912 41318
rect 22616 40282 22672 40284
rect 22696 40282 22752 40284
rect 22776 40282 22832 40284
rect 22856 40282 22912 40284
rect 22616 40230 22662 40282
rect 22662 40230 22672 40282
rect 22696 40230 22726 40282
rect 22726 40230 22738 40282
rect 22738 40230 22752 40282
rect 22776 40230 22790 40282
rect 22790 40230 22802 40282
rect 22802 40230 22832 40282
rect 22856 40230 22866 40282
rect 22866 40230 22912 40282
rect 22616 40228 22672 40230
rect 22696 40228 22752 40230
rect 22776 40228 22832 40230
rect 22856 40228 22912 40230
rect 26956 68026 27012 68028
rect 27036 68026 27092 68028
rect 27116 68026 27172 68028
rect 27196 68026 27252 68028
rect 26956 67974 27002 68026
rect 27002 67974 27012 68026
rect 27036 67974 27066 68026
rect 27066 67974 27078 68026
rect 27078 67974 27092 68026
rect 27116 67974 27130 68026
rect 27130 67974 27142 68026
rect 27142 67974 27172 68026
rect 27196 67974 27206 68026
rect 27206 67974 27252 68026
rect 26956 67972 27012 67974
rect 27036 67972 27092 67974
rect 27116 67972 27172 67974
rect 27196 67972 27252 67974
rect 23570 40568 23626 40624
rect 27616 67482 27672 67484
rect 27696 67482 27752 67484
rect 27776 67482 27832 67484
rect 27856 67482 27912 67484
rect 27616 67430 27662 67482
rect 27662 67430 27672 67482
rect 27696 67430 27726 67482
rect 27726 67430 27738 67482
rect 27738 67430 27752 67482
rect 27776 67430 27790 67482
rect 27790 67430 27802 67482
rect 27802 67430 27832 67482
rect 27856 67430 27866 67482
rect 27866 67430 27912 67482
rect 27616 67428 27672 67430
rect 27696 67428 27752 67430
rect 27776 67428 27832 67430
rect 27856 67428 27912 67430
rect 26956 66938 27012 66940
rect 27036 66938 27092 66940
rect 27116 66938 27172 66940
rect 27196 66938 27252 66940
rect 26956 66886 27002 66938
rect 27002 66886 27012 66938
rect 27036 66886 27066 66938
rect 27066 66886 27078 66938
rect 27078 66886 27092 66938
rect 27116 66886 27130 66938
rect 27130 66886 27142 66938
rect 27142 66886 27172 66938
rect 27196 66886 27206 66938
rect 27206 66886 27252 66938
rect 26956 66884 27012 66886
rect 27036 66884 27092 66886
rect 27116 66884 27172 66886
rect 27196 66884 27252 66886
rect 22616 39194 22672 39196
rect 22696 39194 22752 39196
rect 22776 39194 22832 39196
rect 22856 39194 22912 39196
rect 22616 39142 22662 39194
rect 22662 39142 22672 39194
rect 22696 39142 22726 39194
rect 22726 39142 22738 39194
rect 22738 39142 22752 39194
rect 22776 39142 22790 39194
rect 22790 39142 22802 39194
rect 22802 39142 22832 39194
rect 22856 39142 22866 39194
rect 22866 39142 22912 39194
rect 22616 39140 22672 39142
rect 22696 39140 22752 39142
rect 22776 39140 22832 39142
rect 22856 39140 22912 39142
rect 22616 38106 22672 38108
rect 22696 38106 22752 38108
rect 22776 38106 22832 38108
rect 22856 38106 22912 38108
rect 22616 38054 22662 38106
rect 22662 38054 22672 38106
rect 22696 38054 22726 38106
rect 22726 38054 22738 38106
rect 22738 38054 22752 38106
rect 22776 38054 22790 38106
rect 22790 38054 22802 38106
rect 22802 38054 22832 38106
rect 22856 38054 22866 38106
rect 22866 38054 22912 38106
rect 22616 38052 22672 38054
rect 22696 38052 22752 38054
rect 22776 38052 22832 38054
rect 22856 38052 22912 38054
rect 22616 37018 22672 37020
rect 22696 37018 22752 37020
rect 22776 37018 22832 37020
rect 22856 37018 22912 37020
rect 22616 36966 22662 37018
rect 22662 36966 22672 37018
rect 22696 36966 22726 37018
rect 22726 36966 22738 37018
rect 22738 36966 22752 37018
rect 22776 36966 22790 37018
rect 22790 36966 22802 37018
rect 22802 36966 22832 37018
rect 22856 36966 22866 37018
rect 22866 36966 22912 37018
rect 22616 36964 22672 36966
rect 22696 36964 22752 36966
rect 22776 36964 22832 36966
rect 22856 36964 22912 36966
rect 22616 35930 22672 35932
rect 22696 35930 22752 35932
rect 22776 35930 22832 35932
rect 22856 35930 22912 35932
rect 22616 35878 22662 35930
rect 22662 35878 22672 35930
rect 22696 35878 22726 35930
rect 22726 35878 22738 35930
rect 22738 35878 22752 35930
rect 22776 35878 22790 35930
rect 22790 35878 22802 35930
rect 22802 35878 22832 35930
rect 22856 35878 22866 35930
rect 22866 35878 22912 35930
rect 22616 35876 22672 35878
rect 22696 35876 22752 35878
rect 22776 35876 22832 35878
rect 22856 35876 22912 35878
rect 22616 34842 22672 34844
rect 22696 34842 22752 34844
rect 22776 34842 22832 34844
rect 22856 34842 22912 34844
rect 22616 34790 22662 34842
rect 22662 34790 22672 34842
rect 22696 34790 22726 34842
rect 22726 34790 22738 34842
rect 22738 34790 22752 34842
rect 22776 34790 22790 34842
rect 22790 34790 22802 34842
rect 22802 34790 22832 34842
rect 22856 34790 22866 34842
rect 22866 34790 22912 34842
rect 22616 34788 22672 34790
rect 22696 34788 22752 34790
rect 22776 34788 22832 34790
rect 22856 34788 22912 34790
rect 22616 33754 22672 33756
rect 22696 33754 22752 33756
rect 22776 33754 22832 33756
rect 22856 33754 22912 33756
rect 22616 33702 22662 33754
rect 22662 33702 22672 33754
rect 22696 33702 22726 33754
rect 22726 33702 22738 33754
rect 22738 33702 22752 33754
rect 22776 33702 22790 33754
rect 22790 33702 22802 33754
rect 22802 33702 22832 33754
rect 22856 33702 22866 33754
rect 22866 33702 22912 33754
rect 22616 33700 22672 33702
rect 22696 33700 22752 33702
rect 22776 33700 22832 33702
rect 22856 33700 22912 33702
rect 22616 32666 22672 32668
rect 22696 32666 22752 32668
rect 22776 32666 22832 32668
rect 22856 32666 22912 32668
rect 22616 32614 22662 32666
rect 22662 32614 22672 32666
rect 22696 32614 22726 32666
rect 22726 32614 22738 32666
rect 22738 32614 22752 32666
rect 22776 32614 22790 32666
rect 22790 32614 22802 32666
rect 22802 32614 22832 32666
rect 22856 32614 22866 32666
rect 22866 32614 22912 32666
rect 22616 32612 22672 32614
rect 22696 32612 22752 32614
rect 22776 32612 22832 32614
rect 22856 32612 22912 32614
rect 22616 31578 22672 31580
rect 22696 31578 22752 31580
rect 22776 31578 22832 31580
rect 22856 31578 22912 31580
rect 22616 31526 22662 31578
rect 22662 31526 22672 31578
rect 22696 31526 22726 31578
rect 22726 31526 22738 31578
rect 22738 31526 22752 31578
rect 22776 31526 22790 31578
rect 22790 31526 22802 31578
rect 22802 31526 22832 31578
rect 22856 31526 22866 31578
rect 22866 31526 22912 31578
rect 22616 31524 22672 31526
rect 22696 31524 22752 31526
rect 22776 31524 22832 31526
rect 22856 31524 22912 31526
rect 22616 30490 22672 30492
rect 22696 30490 22752 30492
rect 22776 30490 22832 30492
rect 22856 30490 22912 30492
rect 22616 30438 22662 30490
rect 22662 30438 22672 30490
rect 22696 30438 22726 30490
rect 22726 30438 22738 30490
rect 22738 30438 22752 30490
rect 22776 30438 22790 30490
rect 22790 30438 22802 30490
rect 22802 30438 22832 30490
rect 22856 30438 22866 30490
rect 22866 30438 22912 30490
rect 22616 30436 22672 30438
rect 22696 30436 22752 30438
rect 22776 30436 22832 30438
rect 22856 30436 22912 30438
rect 22616 29402 22672 29404
rect 22696 29402 22752 29404
rect 22776 29402 22832 29404
rect 22856 29402 22912 29404
rect 22616 29350 22662 29402
rect 22662 29350 22672 29402
rect 22696 29350 22726 29402
rect 22726 29350 22738 29402
rect 22738 29350 22752 29402
rect 22776 29350 22790 29402
rect 22790 29350 22802 29402
rect 22802 29350 22832 29402
rect 22856 29350 22866 29402
rect 22866 29350 22912 29402
rect 22616 29348 22672 29350
rect 22696 29348 22752 29350
rect 22776 29348 22832 29350
rect 22856 29348 22912 29350
rect 22616 28314 22672 28316
rect 22696 28314 22752 28316
rect 22776 28314 22832 28316
rect 22856 28314 22912 28316
rect 22616 28262 22662 28314
rect 22662 28262 22672 28314
rect 22696 28262 22726 28314
rect 22726 28262 22738 28314
rect 22738 28262 22752 28314
rect 22776 28262 22790 28314
rect 22790 28262 22802 28314
rect 22802 28262 22832 28314
rect 22856 28262 22866 28314
rect 22866 28262 22912 28314
rect 22616 28260 22672 28262
rect 22696 28260 22752 28262
rect 22776 28260 22832 28262
rect 22856 28260 22912 28262
rect 22616 27226 22672 27228
rect 22696 27226 22752 27228
rect 22776 27226 22832 27228
rect 22856 27226 22912 27228
rect 22616 27174 22662 27226
rect 22662 27174 22672 27226
rect 22696 27174 22726 27226
rect 22726 27174 22738 27226
rect 22738 27174 22752 27226
rect 22776 27174 22790 27226
rect 22790 27174 22802 27226
rect 22802 27174 22832 27226
rect 22856 27174 22866 27226
rect 22866 27174 22912 27226
rect 22616 27172 22672 27174
rect 22696 27172 22752 27174
rect 22776 27172 22832 27174
rect 22856 27172 22912 27174
rect 22616 26138 22672 26140
rect 22696 26138 22752 26140
rect 22776 26138 22832 26140
rect 22856 26138 22912 26140
rect 22616 26086 22662 26138
rect 22662 26086 22672 26138
rect 22696 26086 22726 26138
rect 22726 26086 22738 26138
rect 22738 26086 22752 26138
rect 22776 26086 22790 26138
rect 22790 26086 22802 26138
rect 22802 26086 22832 26138
rect 22856 26086 22866 26138
rect 22866 26086 22912 26138
rect 22616 26084 22672 26086
rect 22696 26084 22752 26086
rect 22776 26084 22832 26086
rect 22856 26084 22912 26086
rect 22616 25050 22672 25052
rect 22696 25050 22752 25052
rect 22776 25050 22832 25052
rect 22856 25050 22912 25052
rect 22616 24998 22662 25050
rect 22662 24998 22672 25050
rect 22696 24998 22726 25050
rect 22726 24998 22738 25050
rect 22738 24998 22752 25050
rect 22776 24998 22790 25050
rect 22790 24998 22802 25050
rect 22802 24998 22832 25050
rect 22856 24998 22866 25050
rect 22866 24998 22912 25050
rect 22616 24996 22672 24998
rect 22696 24996 22752 24998
rect 22776 24996 22832 24998
rect 22856 24996 22912 24998
rect 22616 23962 22672 23964
rect 22696 23962 22752 23964
rect 22776 23962 22832 23964
rect 22856 23962 22912 23964
rect 22616 23910 22662 23962
rect 22662 23910 22672 23962
rect 22696 23910 22726 23962
rect 22726 23910 22738 23962
rect 22738 23910 22752 23962
rect 22776 23910 22790 23962
rect 22790 23910 22802 23962
rect 22802 23910 22832 23962
rect 22856 23910 22866 23962
rect 22866 23910 22912 23962
rect 22616 23908 22672 23910
rect 22696 23908 22752 23910
rect 22776 23908 22832 23910
rect 22856 23908 22912 23910
rect 22616 22874 22672 22876
rect 22696 22874 22752 22876
rect 22776 22874 22832 22876
rect 22856 22874 22912 22876
rect 22616 22822 22662 22874
rect 22662 22822 22672 22874
rect 22696 22822 22726 22874
rect 22726 22822 22738 22874
rect 22738 22822 22752 22874
rect 22776 22822 22790 22874
rect 22790 22822 22802 22874
rect 22802 22822 22832 22874
rect 22856 22822 22866 22874
rect 22866 22822 22912 22874
rect 22616 22820 22672 22822
rect 22696 22820 22752 22822
rect 22776 22820 22832 22822
rect 22856 22820 22912 22822
rect 22616 21786 22672 21788
rect 22696 21786 22752 21788
rect 22776 21786 22832 21788
rect 22856 21786 22912 21788
rect 22616 21734 22662 21786
rect 22662 21734 22672 21786
rect 22696 21734 22726 21786
rect 22726 21734 22738 21786
rect 22738 21734 22752 21786
rect 22776 21734 22790 21786
rect 22790 21734 22802 21786
rect 22802 21734 22832 21786
rect 22856 21734 22866 21786
rect 22866 21734 22912 21786
rect 22616 21732 22672 21734
rect 22696 21732 22752 21734
rect 22776 21732 22832 21734
rect 22856 21732 22912 21734
rect 21956 20154 22012 20156
rect 22036 20154 22092 20156
rect 22116 20154 22172 20156
rect 22196 20154 22252 20156
rect 21956 20102 22002 20154
rect 22002 20102 22012 20154
rect 22036 20102 22066 20154
rect 22066 20102 22078 20154
rect 22078 20102 22092 20154
rect 22116 20102 22130 20154
rect 22130 20102 22142 20154
rect 22142 20102 22172 20154
rect 22196 20102 22206 20154
rect 22206 20102 22252 20154
rect 21956 20100 22012 20102
rect 22036 20100 22092 20102
rect 22116 20100 22172 20102
rect 22196 20100 22252 20102
rect 21956 19066 22012 19068
rect 22036 19066 22092 19068
rect 22116 19066 22172 19068
rect 22196 19066 22252 19068
rect 21956 19014 22002 19066
rect 22002 19014 22012 19066
rect 22036 19014 22066 19066
rect 22066 19014 22078 19066
rect 22078 19014 22092 19066
rect 22116 19014 22130 19066
rect 22130 19014 22142 19066
rect 22142 19014 22172 19066
rect 22196 19014 22206 19066
rect 22206 19014 22252 19066
rect 21956 19012 22012 19014
rect 22036 19012 22092 19014
rect 22116 19012 22172 19014
rect 22196 19012 22252 19014
rect 21956 17978 22012 17980
rect 22036 17978 22092 17980
rect 22116 17978 22172 17980
rect 22196 17978 22252 17980
rect 21956 17926 22002 17978
rect 22002 17926 22012 17978
rect 22036 17926 22066 17978
rect 22066 17926 22078 17978
rect 22078 17926 22092 17978
rect 22116 17926 22130 17978
rect 22130 17926 22142 17978
rect 22142 17926 22172 17978
rect 22196 17926 22206 17978
rect 22206 17926 22252 17978
rect 21956 17924 22012 17926
rect 22036 17924 22092 17926
rect 22116 17924 22172 17926
rect 22196 17924 22252 17926
rect 21956 16890 22012 16892
rect 22036 16890 22092 16892
rect 22116 16890 22172 16892
rect 22196 16890 22252 16892
rect 21956 16838 22002 16890
rect 22002 16838 22012 16890
rect 22036 16838 22066 16890
rect 22066 16838 22078 16890
rect 22078 16838 22092 16890
rect 22116 16838 22130 16890
rect 22130 16838 22142 16890
rect 22142 16838 22172 16890
rect 22196 16838 22206 16890
rect 22206 16838 22252 16890
rect 21956 16836 22012 16838
rect 22036 16836 22092 16838
rect 22116 16836 22172 16838
rect 22196 16836 22252 16838
rect 21956 15802 22012 15804
rect 22036 15802 22092 15804
rect 22116 15802 22172 15804
rect 22196 15802 22252 15804
rect 21956 15750 22002 15802
rect 22002 15750 22012 15802
rect 22036 15750 22066 15802
rect 22066 15750 22078 15802
rect 22078 15750 22092 15802
rect 22116 15750 22130 15802
rect 22130 15750 22142 15802
rect 22142 15750 22172 15802
rect 22196 15750 22206 15802
rect 22206 15750 22252 15802
rect 21956 15748 22012 15750
rect 22036 15748 22092 15750
rect 22116 15748 22172 15750
rect 22196 15748 22252 15750
rect 22374 15000 22430 15056
rect 21956 14714 22012 14716
rect 22036 14714 22092 14716
rect 22116 14714 22172 14716
rect 22196 14714 22252 14716
rect 21956 14662 22002 14714
rect 22002 14662 22012 14714
rect 22036 14662 22066 14714
rect 22066 14662 22078 14714
rect 22078 14662 22092 14714
rect 22116 14662 22130 14714
rect 22130 14662 22142 14714
rect 22142 14662 22172 14714
rect 22196 14662 22206 14714
rect 22206 14662 22252 14714
rect 21956 14660 22012 14662
rect 22036 14660 22092 14662
rect 22116 14660 22172 14662
rect 22196 14660 22252 14662
rect 21956 13626 22012 13628
rect 22036 13626 22092 13628
rect 22116 13626 22172 13628
rect 22196 13626 22252 13628
rect 21956 13574 22002 13626
rect 22002 13574 22012 13626
rect 22036 13574 22066 13626
rect 22066 13574 22078 13626
rect 22078 13574 22092 13626
rect 22116 13574 22130 13626
rect 22130 13574 22142 13626
rect 22142 13574 22172 13626
rect 22196 13574 22206 13626
rect 22206 13574 22252 13626
rect 21956 13572 22012 13574
rect 22036 13572 22092 13574
rect 22116 13572 22172 13574
rect 22196 13572 22252 13574
rect 21956 12538 22012 12540
rect 22036 12538 22092 12540
rect 22116 12538 22172 12540
rect 22196 12538 22252 12540
rect 21956 12486 22002 12538
rect 22002 12486 22012 12538
rect 22036 12486 22066 12538
rect 22066 12486 22078 12538
rect 22078 12486 22092 12538
rect 22116 12486 22130 12538
rect 22130 12486 22142 12538
rect 22142 12486 22172 12538
rect 22196 12486 22206 12538
rect 22206 12486 22252 12538
rect 21956 12484 22012 12486
rect 22036 12484 22092 12486
rect 22116 12484 22172 12486
rect 22196 12484 22252 12486
rect 17616 4378 17672 4380
rect 17696 4378 17752 4380
rect 17776 4378 17832 4380
rect 17856 4378 17912 4380
rect 17616 4326 17662 4378
rect 17662 4326 17672 4378
rect 17696 4326 17726 4378
rect 17726 4326 17738 4378
rect 17738 4326 17752 4378
rect 17776 4326 17790 4378
rect 17790 4326 17802 4378
rect 17802 4326 17832 4378
rect 17856 4326 17866 4378
rect 17866 4326 17912 4378
rect 17616 4324 17672 4326
rect 17696 4324 17752 4326
rect 17776 4324 17832 4326
rect 17856 4324 17912 4326
rect 17616 3290 17672 3292
rect 17696 3290 17752 3292
rect 17776 3290 17832 3292
rect 17856 3290 17912 3292
rect 17616 3238 17662 3290
rect 17662 3238 17672 3290
rect 17696 3238 17726 3290
rect 17726 3238 17738 3290
rect 17738 3238 17752 3290
rect 17776 3238 17790 3290
rect 17790 3238 17802 3290
rect 17802 3238 17832 3290
rect 17856 3238 17866 3290
rect 17866 3238 17912 3290
rect 17616 3236 17672 3238
rect 17696 3236 17752 3238
rect 17776 3236 17832 3238
rect 17856 3236 17912 3238
rect 21956 11450 22012 11452
rect 22036 11450 22092 11452
rect 22116 11450 22172 11452
rect 22196 11450 22252 11452
rect 21956 11398 22002 11450
rect 22002 11398 22012 11450
rect 22036 11398 22066 11450
rect 22066 11398 22078 11450
rect 22078 11398 22092 11450
rect 22116 11398 22130 11450
rect 22130 11398 22142 11450
rect 22142 11398 22172 11450
rect 22196 11398 22206 11450
rect 22206 11398 22252 11450
rect 21956 11396 22012 11398
rect 22036 11396 22092 11398
rect 22116 11396 22172 11398
rect 22196 11396 22252 11398
rect 21956 10362 22012 10364
rect 22036 10362 22092 10364
rect 22116 10362 22172 10364
rect 22196 10362 22252 10364
rect 21956 10310 22002 10362
rect 22002 10310 22012 10362
rect 22036 10310 22066 10362
rect 22066 10310 22078 10362
rect 22078 10310 22092 10362
rect 22116 10310 22130 10362
rect 22130 10310 22142 10362
rect 22142 10310 22172 10362
rect 22196 10310 22206 10362
rect 22206 10310 22252 10362
rect 21956 10308 22012 10310
rect 22036 10308 22092 10310
rect 22116 10308 22172 10310
rect 22196 10308 22252 10310
rect 21956 9274 22012 9276
rect 22036 9274 22092 9276
rect 22116 9274 22172 9276
rect 22196 9274 22252 9276
rect 21956 9222 22002 9274
rect 22002 9222 22012 9274
rect 22036 9222 22066 9274
rect 22066 9222 22078 9274
rect 22078 9222 22092 9274
rect 22116 9222 22130 9274
rect 22130 9222 22142 9274
rect 22142 9222 22172 9274
rect 22196 9222 22206 9274
rect 22206 9222 22252 9274
rect 21956 9220 22012 9222
rect 22036 9220 22092 9222
rect 22116 9220 22172 9222
rect 22196 9220 22252 9222
rect 21956 8186 22012 8188
rect 22036 8186 22092 8188
rect 22116 8186 22172 8188
rect 22196 8186 22252 8188
rect 21956 8134 22002 8186
rect 22002 8134 22012 8186
rect 22036 8134 22066 8186
rect 22066 8134 22078 8186
rect 22078 8134 22092 8186
rect 22116 8134 22130 8186
rect 22130 8134 22142 8186
rect 22142 8134 22172 8186
rect 22196 8134 22206 8186
rect 22206 8134 22252 8186
rect 21956 8132 22012 8134
rect 22036 8132 22092 8134
rect 22116 8132 22172 8134
rect 22196 8132 22252 8134
rect 22616 20698 22672 20700
rect 22696 20698 22752 20700
rect 22776 20698 22832 20700
rect 22856 20698 22912 20700
rect 22616 20646 22662 20698
rect 22662 20646 22672 20698
rect 22696 20646 22726 20698
rect 22726 20646 22738 20698
rect 22738 20646 22752 20698
rect 22776 20646 22790 20698
rect 22790 20646 22802 20698
rect 22802 20646 22832 20698
rect 22856 20646 22866 20698
rect 22866 20646 22912 20698
rect 22616 20644 22672 20646
rect 22696 20644 22752 20646
rect 22776 20644 22832 20646
rect 22856 20644 22912 20646
rect 23386 38700 23388 38720
rect 23388 38700 23440 38720
rect 23440 38700 23442 38720
rect 23386 38664 23442 38700
rect 23386 31048 23442 31104
rect 22616 19610 22672 19612
rect 22696 19610 22752 19612
rect 22776 19610 22832 19612
rect 22856 19610 22912 19612
rect 22616 19558 22662 19610
rect 22662 19558 22672 19610
rect 22696 19558 22726 19610
rect 22726 19558 22738 19610
rect 22738 19558 22752 19610
rect 22776 19558 22790 19610
rect 22790 19558 22802 19610
rect 22802 19558 22832 19610
rect 22856 19558 22866 19610
rect 22866 19558 22912 19610
rect 22616 19556 22672 19558
rect 22696 19556 22752 19558
rect 22776 19556 22832 19558
rect 22856 19556 22912 19558
rect 22616 18522 22672 18524
rect 22696 18522 22752 18524
rect 22776 18522 22832 18524
rect 22856 18522 22912 18524
rect 22616 18470 22662 18522
rect 22662 18470 22672 18522
rect 22696 18470 22726 18522
rect 22726 18470 22738 18522
rect 22738 18470 22752 18522
rect 22776 18470 22790 18522
rect 22790 18470 22802 18522
rect 22802 18470 22832 18522
rect 22856 18470 22866 18522
rect 22866 18470 22912 18522
rect 22616 18468 22672 18470
rect 22696 18468 22752 18470
rect 22776 18468 22832 18470
rect 22856 18468 22912 18470
rect 22616 17434 22672 17436
rect 22696 17434 22752 17436
rect 22776 17434 22832 17436
rect 22856 17434 22912 17436
rect 22616 17382 22662 17434
rect 22662 17382 22672 17434
rect 22696 17382 22726 17434
rect 22726 17382 22738 17434
rect 22738 17382 22752 17434
rect 22776 17382 22790 17434
rect 22790 17382 22802 17434
rect 22802 17382 22832 17434
rect 22856 17382 22866 17434
rect 22866 17382 22912 17434
rect 22616 17380 22672 17382
rect 22696 17380 22752 17382
rect 22776 17380 22832 17382
rect 22856 17380 22912 17382
rect 22616 16346 22672 16348
rect 22696 16346 22752 16348
rect 22776 16346 22832 16348
rect 22856 16346 22912 16348
rect 22616 16294 22662 16346
rect 22662 16294 22672 16346
rect 22696 16294 22726 16346
rect 22726 16294 22738 16346
rect 22738 16294 22752 16346
rect 22776 16294 22790 16346
rect 22790 16294 22802 16346
rect 22802 16294 22832 16346
rect 22856 16294 22866 16346
rect 22866 16294 22912 16346
rect 22616 16292 22672 16294
rect 22696 16292 22752 16294
rect 22776 16292 22832 16294
rect 22856 16292 22912 16294
rect 22616 15258 22672 15260
rect 22696 15258 22752 15260
rect 22776 15258 22832 15260
rect 22856 15258 22912 15260
rect 22616 15206 22662 15258
rect 22662 15206 22672 15258
rect 22696 15206 22726 15258
rect 22726 15206 22738 15258
rect 22738 15206 22752 15258
rect 22776 15206 22790 15258
rect 22790 15206 22802 15258
rect 22802 15206 22832 15258
rect 22856 15206 22866 15258
rect 22866 15206 22912 15258
rect 22616 15204 22672 15206
rect 22696 15204 22752 15206
rect 22776 15204 22832 15206
rect 22856 15204 22912 15206
rect 22616 14170 22672 14172
rect 22696 14170 22752 14172
rect 22776 14170 22832 14172
rect 22856 14170 22912 14172
rect 22616 14118 22662 14170
rect 22662 14118 22672 14170
rect 22696 14118 22726 14170
rect 22726 14118 22738 14170
rect 22738 14118 22752 14170
rect 22776 14118 22790 14170
rect 22790 14118 22802 14170
rect 22802 14118 22832 14170
rect 22856 14118 22866 14170
rect 22866 14118 22912 14170
rect 22616 14116 22672 14118
rect 22696 14116 22752 14118
rect 22776 14116 22832 14118
rect 22856 14116 22912 14118
rect 22616 13082 22672 13084
rect 22696 13082 22752 13084
rect 22776 13082 22832 13084
rect 22856 13082 22912 13084
rect 22616 13030 22662 13082
rect 22662 13030 22672 13082
rect 22696 13030 22726 13082
rect 22726 13030 22738 13082
rect 22738 13030 22752 13082
rect 22776 13030 22790 13082
rect 22790 13030 22802 13082
rect 22802 13030 22832 13082
rect 22856 13030 22866 13082
rect 22866 13030 22912 13082
rect 22616 13028 22672 13030
rect 22696 13028 22752 13030
rect 22776 13028 22832 13030
rect 22856 13028 22912 13030
rect 23846 39344 23902 39400
rect 23754 36624 23810 36680
rect 24306 38836 24308 38856
rect 24308 38836 24360 38856
rect 24360 38836 24362 38856
rect 24306 38800 24362 38836
rect 24582 38936 24638 38992
rect 24766 38412 24822 38448
rect 24766 38392 24768 38412
rect 24768 38392 24820 38412
rect 24820 38392 24822 38412
rect 24950 26288 25006 26344
rect 25226 37984 25282 38040
rect 27616 66394 27672 66396
rect 27696 66394 27752 66396
rect 27776 66394 27832 66396
rect 27856 66394 27912 66396
rect 27616 66342 27662 66394
rect 27662 66342 27672 66394
rect 27696 66342 27726 66394
rect 27726 66342 27738 66394
rect 27738 66342 27752 66394
rect 27776 66342 27790 66394
rect 27790 66342 27802 66394
rect 27802 66342 27832 66394
rect 27856 66342 27866 66394
rect 27866 66342 27912 66394
rect 27616 66340 27672 66342
rect 27696 66340 27752 66342
rect 27776 66340 27832 66342
rect 27856 66340 27912 66342
rect 26956 65850 27012 65852
rect 27036 65850 27092 65852
rect 27116 65850 27172 65852
rect 27196 65850 27252 65852
rect 26956 65798 27002 65850
rect 27002 65798 27012 65850
rect 27036 65798 27066 65850
rect 27066 65798 27078 65850
rect 27078 65798 27092 65850
rect 27116 65798 27130 65850
rect 27130 65798 27142 65850
rect 27142 65798 27172 65850
rect 27196 65798 27206 65850
rect 27206 65798 27252 65850
rect 26956 65796 27012 65798
rect 27036 65796 27092 65798
rect 27116 65796 27172 65798
rect 27196 65796 27252 65798
rect 27616 65306 27672 65308
rect 27696 65306 27752 65308
rect 27776 65306 27832 65308
rect 27856 65306 27912 65308
rect 27616 65254 27662 65306
rect 27662 65254 27672 65306
rect 27696 65254 27726 65306
rect 27726 65254 27738 65306
rect 27738 65254 27752 65306
rect 27776 65254 27790 65306
rect 27790 65254 27802 65306
rect 27802 65254 27832 65306
rect 27856 65254 27866 65306
rect 27866 65254 27912 65306
rect 27616 65252 27672 65254
rect 27696 65252 27752 65254
rect 27776 65252 27832 65254
rect 27856 65252 27912 65254
rect 26956 64762 27012 64764
rect 27036 64762 27092 64764
rect 27116 64762 27172 64764
rect 27196 64762 27252 64764
rect 26956 64710 27002 64762
rect 27002 64710 27012 64762
rect 27036 64710 27066 64762
rect 27066 64710 27078 64762
rect 27078 64710 27092 64762
rect 27116 64710 27130 64762
rect 27130 64710 27142 64762
rect 27142 64710 27172 64762
rect 27196 64710 27206 64762
rect 27206 64710 27252 64762
rect 26956 64708 27012 64710
rect 27036 64708 27092 64710
rect 27116 64708 27172 64710
rect 27196 64708 27252 64710
rect 27616 64218 27672 64220
rect 27696 64218 27752 64220
rect 27776 64218 27832 64220
rect 27856 64218 27912 64220
rect 27616 64166 27662 64218
rect 27662 64166 27672 64218
rect 27696 64166 27726 64218
rect 27726 64166 27738 64218
rect 27738 64166 27752 64218
rect 27776 64166 27790 64218
rect 27790 64166 27802 64218
rect 27802 64166 27832 64218
rect 27856 64166 27866 64218
rect 27866 64166 27912 64218
rect 27616 64164 27672 64166
rect 27696 64164 27752 64166
rect 27776 64164 27832 64166
rect 27856 64164 27912 64166
rect 26956 63674 27012 63676
rect 27036 63674 27092 63676
rect 27116 63674 27172 63676
rect 27196 63674 27252 63676
rect 26956 63622 27002 63674
rect 27002 63622 27012 63674
rect 27036 63622 27066 63674
rect 27066 63622 27078 63674
rect 27078 63622 27092 63674
rect 27116 63622 27130 63674
rect 27130 63622 27142 63674
rect 27142 63622 27172 63674
rect 27196 63622 27206 63674
rect 27206 63622 27252 63674
rect 26956 63620 27012 63622
rect 27036 63620 27092 63622
rect 27116 63620 27172 63622
rect 27196 63620 27252 63622
rect 27616 63130 27672 63132
rect 27696 63130 27752 63132
rect 27776 63130 27832 63132
rect 27856 63130 27912 63132
rect 27616 63078 27662 63130
rect 27662 63078 27672 63130
rect 27696 63078 27726 63130
rect 27726 63078 27738 63130
rect 27738 63078 27752 63130
rect 27776 63078 27790 63130
rect 27790 63078 27802 63130
rect 27802 63078 27832 63130
rect 27856 63078 27866 63130
rect 27866 63078 27912 63130
rect 27616 63076 27672 63078
rect 27696 63076 27752 63078
rect 27776 63076 27832 63078
rect 27856 63076 27912 63078
rect 26956 62586 27012 62588
rect 27036 62586 27092 62588
rect 27116 62586 27172 62588
rect 27196 62586 27252 62588
rect 26956 62534 27002 62586
rect 27002 62534 27012 62586
rect 27036 62534 27066 62586
rect 27066 62534 27078 62586
rect 27078 62534 27092 62586
rect 27116 62534 27130 62586
rect 27130 62534 27142 62586
rect 27142 62534 27172 62586
rect 27196 62534 27206 62586
rect 27206 62534 27252 62586
rect 26956 62532 27012 62534
rect 27036 62532 27092 62534
rect 27116 62532 27172 62534
rect 27196 62532 27252 62534
rect 26956 61498 27012 61500
rect 27036 61498 27092 61500
rect 27116 61498 27172 61500
rect 27196 61498 27252 61500
rect 26956 61446 27002 61498
rect 27002 61446 27012 61498
rect 27036 61446 27066 61498
rect 27066 61446 27078 61498
rect 27078 61446 27092 61498
rect 27116 61446 27130 61498
rect 27130 61446 27142 61498
rect 27142 61446 27172 61498
rect 27196 61446 27206 61498
rect 27206 61446 27252 61498
rect 26956 61444 27012 61446
rect 27036 61444 27092 61446
rect 27116 61444 27172 61446
rect 27196 61444 27252 61446
rect 26956 60410 27012 60412
rect 27036 60410 27092 60412
rect 27116 60410 27172 60412
rect 27196 60410 27252 60412
rect 26956 60358 27002 60410
rect 27002 60358 27012 60410
rect 27036 60358 27066 60410
rect 27066 60358 27078 60410
rect 27078 60358 27092 60410
rect 27116 60358 27130 60410
rect 27130 60358 27142 60410
rect 27142 60358 27172 60410
rect 27196 60358 27206 60410
rect 27206 60358 27252 60410
rect 26956 60356 27012 60358
rect 27036 60356 27092 60358
rect 27116 60356 27172 60358
rect 27196 60356 27252 60358
rect 26956 59322 27012 59324
rect 27036 59322 27092 59324
rect 27116 59322 27172 59324
rect 27196 59322 27252 59324
rect 26956 59270 27002 59322
rect 27002 59270 27012 59322
rect 27036 59270 27066 59322
rect 27066 59270 27078 59322
rect 27078 59270 27092 59322
rect 27116 59270 27130 59322
rect 27130 59270 27142 59322
rect 27142 59270 27172 59322
rect 27196 59270 27206 59322
rect 27206 59270 27252 59322
rect 26956 59268 27012 59270
rect 27036 59268 27092 59270
rect 27116 59268 27172 59270
rect 27196 59268 27252 59270
rect 27616 62042 27672 62044
rect 27696 62042 27752 62044
rect 27776 62042 27832 62044
rect 27856 62042 27912 62044
rect 27616 61990 27662 62042
rect 27662 61990 27672 62042
rect 27696 61990 27726 62042
rect 27726 61990 27738 62042
rect 27738 61990 27752 62042
rect 27776 61990 27790 62042
rect 27790 61990 27802 62042
rect 27802 61990 27832 62042
rect 27856 61990 27866 62042
rect 27866 61990 27912 62042
rect 27616 61988 27672 61990
rect 27696 61988 27752 61990
rect 27776 61988 27832 61990
rect 27856 61988 27912 61990
rect 27616 60954 27672 60956
rect 27696 60954 27752 60956
rect 27776 60954 27832 60956
rect 27856 60954 27912 60956
rect 27616 60902 27662 60954
rect 27662 60902 27672 60954
rect 27696 60902 27726 60954
rect 27726 60902 27738 60954
rect 27738 60902 27752 60954
rect 27776 60902 27790 60954
rect 27790 60902 27802 60954
rect 27802 60902 27832 60954
rect 27856 60902 27866 60954
rect 27866 60902 27912 60954
rect 27616 60900 27672 60902
rect 27696 60900 27752 60902
rect 27776 60900 27832 60902
rect 27856 60900 27912 60902
rect 26956 58234 27012 58236
rect 27036 58234 27092 58236
rect 27116 58234 27172 58236
rect 27196 58234 27252 58236
rect 26956 58182 27002 58234
rect 27002 58182 27012 58234
rect 27036 58182 27066 58234
rect 27066 58182 27078 58234
rect 27078 58182 27092 58234
rect 27116 58182 27130 58234
rect 27130 58182 27142 58234
rect 27142 58182 27172 58234
rect 27196 58182 27206 58234
rect 27206 58182 27252 58234
rect 26956 58180 27012 58182
rect 27036 58180 27092 58182
rect 27116 58180 27172 58182
rect 27196 58180 27252 58182
rect 26956 57146 27012 57148
rect 27036 57146 27092 57148
rect 27116 57146 27172 57148
rect 27196 57146 27252 57148
rect 26956 57094 27002 57146
rect 27002 57094 27012 57146
rect 27036 57094 27066 57146
rect 27066 57094 27078 57146
rect 27078 57094 27092 57146
rect 27116 57094 27130 57146
rect 27130 57094 27142 57146
rect 27142 57094 27172 57146
rect 27196 57094 27206 57146
rect 27206 57094 27252 57146
rect 26956 57092 27012 57094
rect 27036 57092 27092 57094
rect 27116 57092 27172 57094
rect 27196 57092 27252 57094
rect 26956 56058 27012 56060
rect 27036 56058 27092 56060
rect 27116 56058 27172 56060
rect 27196 56058 27252 56060
rect 26956 56006 27002 56058
rect 27002 56006 27012 56058
rect 27036 56006 27066 56058
rect 27066 56006 27078 56058
rect 27078 56006 27092 56058
rect 27116 56006 27130 56058
rect 27130 56006 27142 56058
rect 27142 56006 27172 56058
rect 27196 56006 27206 56058
rect 27206 56006 27252 56058
rect 26956 56004 27012 56006
rect 27036 56004 27092 56006
rect 27116 56004 27172 56006
rect 27196 56004 27252 56006
rect 26956 54970 27012 54972
rect 27036 54970 27092 54972
rect 27116 54970 27172 54972
rect 27196 54970 27252 54972
rect 26956 54918 27002 54970
rect 27002 54918 27012 54970
rect 27036 54918 27066 54970
rect 27066 54918 27078 54970
rect 27078 54918 27092 54970
rect 27116 54918 27130 54970
rect 27130 54918 27142 54970
rect 27142 54918 27172 54970
rect 27196 54918 27206 54970
rect 27206 54918 27252 54970
rect 26956 54916 27012 54918
rect 27036 54916 27092 54918
rect 27116 54916 27172 54918
rect 27196 54916 27252 54918
rect 26956 53882 27012 53884
rect 27036 53882 27092 53884
rect 27116 53882 27172 53884
rect 27196 53882 27252 53884
rect 26956 53830 27002 53882
rect 27002 53830 27012 53882
rect 27036 53830 27066 53882
rect 27066 53830 27078 53882
rect 27078 53830 27092 53882
rect 27116 53830 27130 53882
rect 27130 53830 27142 53882
rect 27142 53830 27172 53882
rect 27196 53830 27206 53882
rect 27206 53830 27252 53882
rect 26956 53828 27012 53830
rect 27036 53828 27092 53830
rect 27116 53828 27172 53830
rect 27196 53828 27252 53830
rect 22616 11994 22672 11996
rect 22696 11994 22752 11996
rect 22776 11994 22832 11996
rect 22856 11994 22912 11996
rect 22616 11942 22662 11994
rect 22662 11942 22672 11994
rect 22696 11942 22726 11994
rect 22726 11942 22738 11994
rect 22738 11942 22752 11994
rect 22776 11942 22790 11994
rect 22790 11942 22802 11994
rect 22802 11942 22832 11994
rect 22856 11942 22866 11994
rect 22866 11942 22912 11994
rect 22616 11940 22672 11942
rect 22696 11940 22752 11942
rect 22776 11940 22832 11942
rect 22856 11940 22912 11942
rect 22616 10906 22672 10908
rect 22696 10906 22752 10908
rect 22776 10906 22832 10908
rect 22856 10906 22912 10908
rect 22616 10854 22662 10906
rect 22662 10854 22672 10906
rect 22696 10854 22726 10906
rect 22726 10854 22738 10906
rect 22738 10854 22752 10906
rect 22776 10854 22790 10906
rect 22790 10854 22802 10906
rect 22802 10854 22832 10906
rect 22856 10854 22866 10906
rect 22866 10854 22912 10906
rect 22616 10852 22672 10854
rect 22696 10852 22752 10854
rect 22776 10852 22832 10854
rect 22856 10852 22912 10854
rect 22616 9818 22672 9820
rect 22696 9818 22752 9820
rect 22776 9818 22832 9820
rect 22856 9818 22912 9820
rect 22616 9766 22662 9818
rect 22662 9766 22672 9818
rect 22696 9766 22726 9818
rect 22726 9766 22738 9818
rect 22738 9766 22752 9818
rect 22776 9766 22790 9818
rect 22790 9766 22802 9818
rect 22802 9766 22832 9818
rect 22856 9766 22866 9818
rect 22866 9766 22912 9818
rect 22616 9764 22672 9766
rect 22696 9764 22752 9766
rect 22776 9764 22832 9766
rect 22856 9764 22912 9766
rect 22616 8730 22672 8732
rect 22696 8730 22752 8732
rect 22776 8730 22832 8732
rect 22856 8730 22912 8732
rect 22616 8678 22662 8730
rect 22662 8678 22672 8730
rect 22696 8678 22726 8730
rect 22726 8678 22738 8730
rect 22738 8678 22752 8730
rect 22776 8678 22790 8730
rect 22790 8678 22802 8730
rect 22802 8678 22832 8730
rect 22856 8678 22866 8730
rect 22866 8678 22912 8730
rect 22616 8676 22672 8678
rect 22696 8676 22752 8678
rect 22776 8676 22832 8678
rect 22856 8676 22912 8678
rect 21956 7098 22012 7100
rect 22036 7098 22092 7100
rect 22116 7098 22172 7100
rect 22196 7098 22252 7100
rect 21956 7046 22002 7098
rect 22002 7046 22012 7098
rect 22036 7046 22066 7098
rect 22066 7046 22078 7098
rect 22078 7046 22092 7098
rect 22116 7046 22130 7098
rect 22130 7046 22142 7098
rect 22142 7046 22172 7098
rect 22196 7046 22206 7098
rect 22206 7046 22252 7098
rect 21956 7044 22012 7046
rect 22036 7044 22092 7046
rect 22116 7044 22172 7046
rect 22196 7044 22252 7046
rect 21956 6010 22012 6012
rect 22036 6010 22092 6012
rect 22116 6010 22172 6012
rect 22196 6010 22252 6012
rect 21956 5958 22002 6010
rect 22002 5958 22012 6010
rect 22036 5958 22066 6010
rect 22066 5958 22078 6010
rect 22078 5958 22092 6010
rect 22116 5958 22130 6010
rect 22130 5958 22142 6010
rect 22142 5958 22172 6010
rect 22196 5958 22206 6010
rect 22206 5958 22252 6010
rect 21956 5956 22012 5958
rect 22036 5956 22092 5958
rect 22116 5956 22172 5958
rect 22196 5956 22252 5958
rect 22616 7642 22672 7644
rect 22696 7642 22752 7644
rect 22776 7642 22832 7644
rect 22856 7642 22912 7644
rect 22616 7590 22662 7642
rect 22662 7590 22672 7642
rect 22696 7590 22726 7642
rect 22726 7590 22738 7642
rect 22738 7590 22752 7642
rect 22776 7590 22790 7642
rect 22790 7590 22802 7642
rect 22802 7590 22832 7642
rect 22856 7590 22866 7642
rect 22866 7590 22912 7642
rect 22616 7588 22672 7590
rect 22696 7588 22752 7590
rect 22776 7588 22832 7590
rect 22856 7588 22912 7590
rect 22616 6554 22672 6556
rect 22696 6554 22752 6556
rect 22776 6554 22832 6556
rect 22856 6554 22912 6556
rect 22616 6502 22662 6554
rect 22662 6502 22672 6554
rect 22696 6502 22726 6554
rect 22726 6502 22738 6554
rect 22738 6502 22752 6554
rect 22776 6502 22790 6554
rect 22790 6502 22802 6554
rect 22802 6502 22832 6554
rect 22856 6502 22866 6554
rect 22866 6502 22912 6554
rect 22616 6500 22672 6502
rect 22696 6500 22752 6502
rect 22776 6500 22832 6502
rect 22856 6500 22912 6502
rect 22616 5466 22672 5468
rect 22696 5466 22752 5468
rect 22776 5466 22832 5468
rect 22856 5466 22912 5468
rect 22616 5414 22662 5466
rect 22662 5414 22672 5466
rect 22696 5414 22726 5466
rect 22726 5414 22738 5466
rect 22738 5414 22752 5466
rect 22776 5414 22790 5466
rect 22790 5414 22802 5466
rect 22802 5414 22832 5466
rect 22856 5414 22866 5466
rect 22866 5414 22912 5466
rect 22616 5412 22672 5414
rect 22696 5412 22752 5414
rect 22776 5412 22832 5414
rect 22856 5412 22912 5414
rect 21956 4922 22012 4924
rect 22036 4922 22092 4924
rect 22116 4922 22172 4924
rect 22196 4922 22252 4924
rect 21956 4870 22002 4922
rect 22002 4870 22012 4922
rect 22036 4870 22066 4922
rect 22066 4870 22078 4922
rect 22078 4870 22092 4922
rect 22116 4870 22130 4922
rect 22130 4870 22142 4922
rect 22142 4870 22172 4922
rect 22196 4870 22206 4922
rect 22206 4870 22252 4922
rect 21956 4868 22012 4870
rect 22036 4868 22092 4870
rect 22116 4868 22172 4870
rect 22196 4868 22252 4870
rect 22616 4378 22672 4380
rect 22696 4378 22752 4380
rect 22776 4378 22832 4380
rect 22856 4378 22912 4380
rect 22616 4326 22662 4378
rect 22662 4326 22672 4378
rect 22696 4326 22726 4378
rect 22726 4326 22738 4378
rect 22738 4326 22752 4378
rect 22776 4326 22790 4378
rect 22790 4326 22802 4378
rect 22802 4326 22832 4378
rect 22856 4326 22866 4378
rect 22866 4326 22912 4378
rect 22616 4324 22672 4326
rect 22696 4324 22752 4326
rect 22776 4324 22832 4326
rect 22856 4324 22912 4326
rect 21956 3834 22012 3836
rect 22036 3834 22092 3836
rect 22116 3834 22172 3836
rect 22196 3834 22252 3836
rect 21956 3782 22002 3834
rect 22002 3782 22012 3834
rect 22036 3782 22066 3834
rect 22066 3782 22078 3834
rect 22078 3782 22092 3834
rect 22116 3782 22130 3834
rect 22130 3782 22142 3834
rect 22142 3782 22172 3834
rect 22196 3782 22206 3834
rect 22206 3782 22252 3834
rect 21956 3780 22012 3782
rect 22036 3780 22092 3782
rect 22116 3780 22172 3782
rect 22196 3780 22252 3782
rect 22616 3290 22672 3292
rect 22696 3290 22752 3292
rect 22776 3290 22832 3292
rect 22856 3290 22912 3292
rect 22616 3238 22662 3290
rect 22662 3238 22672 3290
rect 22696 3238 22726 3290
rect 22726 3238 22738 3290
rect 22738 3238 22752 3290
rect 22776 3238 22790 3290
rect 22790 3238 22802 3290
rect 22802 3238 22832 3290
rect 22856 3238 22866 3290
rect 22866 3238 22912 3290
rect 22616 3236 22672 3238
rect 22696 3236 22752 3238
rect 22776 3236 22832 3238
rect 22856 3236 22912 3238
rect 16956 2746 17012 2748
rect 17036 2746 17092 2748
rect 17116 2746 17172 2748
rect 17196 2746 17252 2748
rect 16956 2694 17002 2746
rect 17002 2694 17012 2746
rect 17036 2694 17066 2746
rect 17066 2694 17078 2746
rect 17078 2694 17092 2746
rect 17116 2694 17130 2746
rect 17130 2694 17142 2746
rect 17142 2694 17172 2746
rect 17196 2694 17206 2746
rect 17206 2694 17252 2746
rect 16956 2692 17012 2694
rect 17036 2692 17092 2694
rect 17116 2692 17172 2694
rect 17196 2692 17252 2694
rect 21956 2746 22012 2748
rect 22036 2746 22092 2748
rect 22116 2746 22172 2748
rect 22196 2746 22252 2748
rect 21956 2694 22002 2746
rect 22002 2694 22012 2746
rect 22036 2694 22066 2746
rect 22066 2694 22078 2746
rect 22078 2694 22092 2746
rect 22116 2694 22130 2746
rect 22130 2694 22142 2746
rect 22142 2694 22172 2746
rect 22196 2694 22206 2746
rect 22206 2694 22252 2746
rect 21956 2692 22012 2694
rect 22036 2692 22092 2694
rect 22116 2692 22172 2694
rect 22196 2692 22252 2694
rect 24858 12144 24914 12200
rect 26956 52794 27012 52796
rect 27036 52794 27092 52796
rect 27116 52794 27172 52796
rect 27196 52794 27252 52796
rect 26956 52742 27002 52794
rect 27002 52742 27012 52794
rect 27036 52742 27066 52794
rect 27066 52742 27078 52794
rect 27078 52742 27092 52794
rect 27116 52742 27130 52794
rect 27130 52742 27142 52794
rect 27142 52742 27172 52794
rect 27196 52742 27206 52794
rect 27206 52742 27252 52794
rect 26956 52740 27012 52742
rect 27036 52740 27092 52742
rect 27116 52740 27172 52742
rect 27196 52740 27252 52742
rect 26956 51706 27012 51708
rect 27036 51706 27092 51708
rect 27116 51706 27172 51708
rect 27196 51706 27252 51708
rect 26956 51654 27002 51706
rect 27002 51654 27012 51706
rect 27036 51654 27066 51706
rect 27066 51654 27078 51706
rect 27078 51654 27092 51706
rect 27116 51654 27130 51706
rect 27130 51654 27142 51706
rect 27142 51654 27172 51706
rect 27196 51654 27206 51706
rect 27206 51654 27252 51706
rect 26956 51652 27012 51654
rect 27036 51652 27092 51654
rect 27116 51652 27172 51654
rect 27196 51652 27252 51654
rect 26956 50618 27012 50620
rect 27036 50618 27092 50620
rect 27116 50618 27172 50620
rect 27196 50618 27252 50620
rect 26956 50566 27002 50618
rect 27002 50566 27012 50618
rect 27036 50566 27066 50618
rect 27066 50566 27078 50618
rect 27078 50566 27092 50618
rect 27116 50566 27130 50618
rect 27130 50566 27142 50618
rect 27142 50566 27172 50618
rect 27196 50566 27206 50618
rect 27206 50566 27252 50618
rect 26956 50564 27012 50566
rect 27036 50564 27092 50566
rect 27116 50564 27172 50566
rect 27196 50564 27252 50566
rect 26956 49530 27012 49532
rect 27036 49530 27092 49532
rect 27116 49530 27172 49532
rect 27196 49530 27252 49532
rect 26956 49478 27002 49530
rect 27002 49478 27012 49530
rect 27036 49478 27066 49530
rect 27066 49478 27078 49530
rect 27078 49478 27092 49530
rect 27116 49478 27130 49530
rect 27130 49478 27142 49530
rect 27142 49478 27172 49530
rect 27196 49478 27206 49530
rect 27206 49478 27252 49530
rect 26956 49476 27012 49478
rect 27036 49476 27092 49478
rect 27116 49476 27172 49478
rect 27196 49476 27252 49478
rect 26956 48442 27012 48444
rect 27036 48442 27092 48444
rect 27116 48442 27172 48444
rect 27196 48442 27252 48444
rect 26956 48390 27002 48442
rect 27002 48390 27012 48442
rect 27036 48390 27066 48442
rect 27066 48390 27078 48442
rect 27078 48390 27092 48442
rect 27116 48390 27130 48442
rect 27130 48390 27142 48442
rect 27142 48390 27172 48442
rect 27196 48390 27206 48442
rect 27206 48390 27252 48442
rect 26956 48388 27012 48390
rect 27036 48388 27092 48390
rect 27116 48388 27172 48390
rect 27196 48388 27252 48390
rect 26956 47354 27012 47356
rect 27036 47354 27092 47356
rect 27116 47354 27172 47356
rect 27196 47354 27252 47356
rect 26956 47302 27002 47354
rect 27002 47302 27012 47354
rect 27036 47302 27066 47354
rect 27066 47302 27078 47354
rect 27078 47302 27092 47354
rect 27116 47302 27130 47354
rect 27130 47302 27142 47354
rect 27142 47302 27172 47354
rect 27196 47302 27206 47354
rect 27206 47302 27252 47354
rect 26956 47300 27012 47302
rect 27036 47300 27092 47302
rect 27116 47300 27172 47302
rect 27196 47300 27252 47302
rect 26956 46266 27012 46268
rect 27036 46266 27092 46268
rect 27116 46266 27172 46268
rect 27196 46266 27252 46268
rect 26956 46214 27002 46266
rect 27002 46214 27012 46266
rect 27036 46214 27066 46266
rect 27066 46214 27078 46266
rect 27078 46214 27092 46266
rect 27116 46214 27130 46266
rect 27130 46214 27142 46266
rect 27142 46214 27172 46266
rect 27196 46214 27206 46266
rect 27206 46214 27252 46266
rect 26956 46212 27012 46214
rect 27036 46212 27092 46214
rect 27116 46212 27172 46214
rect 27196 46212 27252 46214
rect 26956 45178 27012 45180
rect 27036 45178 27092 45180
rect 27116 45178 27172 45180
rect 27196 45178 27252 45180
rect 26956 45126 27002 45178
rect 27002 45126 27012 45178
rect 27036 45126 27066 45178
rect 27066 45126 27078 45178
rect 27078 45126 27092 45178
rect 27116 45126 27130 45178
rect 27130 45126 27142 45178
rect 27142 45126 27172 45178
rect 27196 45126 27206 45178
rect 27206 45126 27252 45178
rect 26956 45124 27012 45126
rect 27036 45124 27092 45126
rect 27116 45124 27172 45126
rect 27196 45124 27252 45126
rect 26956 44090 27012 44092
rect 27036 44090 27092 44092
rect 27116 44090 27172 44092
rect 27196 44090 27252 44092
rect 26956 44038 27002 44090
rect 27002 44038 27012 44090
rect 27036 44038 27066 44090
rect 27066 44038 27078 44090
rect 27078 44038 27092 44090
rect 27116 44038 27130 44090
rect 27130 44038 27142 44090
rect 27142 44038 27172 44090
rect 27196 44038 27206 44090
rect 27206 44038 27252 44090
rect 26956 44036 27012 44038
rect 27036 44036 27092 44038
rect 27116 44036 27172 44038
rect 27196 44036 27252 44038
rect 26956 43002 27012 43004
rect 27036 43002 27092 43004
rect 27116 43002 27172 43004
rect 27196 43002 27252 43004
rect 26956 42950 27002 43002
rect 27002 42950 27012 43002
rect 27036 42950 27066 43002
rect 27066 42950 27078 43002
rect 27078 42950 27092 43002
rect 27116 42950 27130 43002
rect 27130 42950 27142 43002
rect 27142 42950 27172 43002
rect 27196 42950 27206 43002
rect 27206 42950 27252 43002
rect 26956 42948 27012 42950
rect 27036 42948 27092 42950
rect 27116 42948 27172 42950
rect 27196 42948 27252 42950
rect 26956 41914 27012 41916
rect 27036 41914 27092 41916
rect 27116 41914 27172 41916
rect 27196 41914 27252 41916
rect 26956 41862 27002 41914
rect 27002 41862 27012 41914
rect 27036 41862 27066 41914
rect 27066 41862 27078 41914
rect 27078 41862 27092 41914
rect 27116 41862 27130 41914
rect 27130 41862 27142 41914
rect 27142 41862 27172 41914
rect 27196 41862 27206 41914
rect 27206 41862 27252 41914
rect 26956 41860 27012 41862
rect 27036 41860 27092 41862
rect 27116 41860 27172 41862
rect 27196 41860 27252 41862
rect 26956 40826 27012 40828
rect 27036 40826 27092 40828
rect 27116 40826 27172 40828
rect 27196 40826 27252 40828
rect 26956 40774 27002 40826
rect 27002 40774 27012 40826
rect 27036 40774 27066 40826
rect 27066 40774 27078 40826
rect 27078 40774 27092 40826
rect 27116 40774 27130 40826
rect 27130 40774 27142 40826
rect 27142 40774 27172 40826
rect 27196 40774 27206 40826
rect 27206 40774 27252 40826
rect 26956 40772 27012 40774
rect 27036 40772 27092 40774
rect 27116 40772 27172 40774
rect 27196 40772 27252 40774
rect 26956 39738 27012 39740
rect 27036 39738 27092 39740
rect 27116 39738 27172 39740
rect 27196 39738 27252 39740
rect 26956 39686 27002 39738
rect 27002 39686 27012 39738
rect 27036 39686 27066 39738
rect 27066 39686 27078 39738
rect 27078 39686 27092 39738
rect 27116 39686 27130 39738
rect 27130 39686 27142 39738
rect 27142 39686 27172 39738
rect 27196 39686 27206 39738
rect 27206 39686 27252 39738
rect 26956 39684 27012 39686
rect 27036 39684 27092 39686
rect 27116 39684 27172 39686
rect 27196 39684 27252 39686
rect 26956 38650 27012 38652
rect 27036 38650 27092 38652
rect 27116 38650 27172 38652
rect 27196 38650 27252 38652
rect 26956 38598 27002 38650
rect 27002 38598 27012 38650
rect 27036 38598 27066 38650
rect 27066 38598 27078 38650
rect 27078 38598 27092 38650
rect 27116 38598 27130 38650
rect 27130 38598 27142 38650
rect 27142 38598 27172 38650
rect 27196 38598 27206 38650
rect 27206 38598 27252 38650
rect 26956 38596 27012 38598
rect 27036 38596 27092 38598
rect 27116 38596 27172 38598
rect 27196 38596 27252 38598
rect 27616 59866 27672 59868
rect 27696 59866 27752 59868
rect 27776 59866 27832 59868
rect 27856 59866 27912 59868
rect 27616 59814 27662 59866
rect 27662 59814 27672 59866
rect 27696 59814 27726 59866
rect 27726 59814 27738 59866
rect 27738 59814 27752 59866
rect 27776 59814 27790 59866
rect 27790 59814 27802 59866
rect 27802 59814 27832 59866
rect 27856 59814 27866 59866
rect 27866 59814 27912 59866
rect 27616 59812 27672 59814
rect 27696 59812 27752 59814
rect 27776 59812 27832 59814
rect 27856 59812 27912 59814
rect 27616 58778 27672 58780
rect 27696 58778 27752 58780
rect 27776 58778 27832 58780
rect 27856 58778 27912 58780
rect 27616 58726 27662 58778
rect 27662 58726 27672 58778
rect 27696 58726 27726 58778
rect 27726 58726 27738 58778
rect 27738 58726 27752 58778
rect 27776 58726 27790 58778
rect 27790 58726 27802 58778
rect 27802 58726 27832 58778
rect 27856 58726 27866 58778
rect 27866 58726 27912 58778
rect 27616 58724 27672 58726
rect 27696 58724 27752 58726
rect 27776 58724 27832 58726
rect 27856 58724 27912 58726
rect 26956 37562 27012 37564
rect 27036 37562 27092 37564
rect 27116 37562 27172 37564
rect 27196 37562 27252 37564
rect 26956 37510 27002 37562
rect 27002 37510 27012 37562
rect 27036 37510 27066 37562
rect 27066 37510 27078 37562
rect 27078 37510 27092 37562
rect 27116 37510 27130 37562
rect 27130 37510 27142 37562
rect 27142 37510 27172 37562
rect 27196 37510 27206 37562
rect 27206 37510 27252 37562
rect 26956 37508 27012 37510
rect 27036 37508 27092 37510
rect 27116 37508 27172 37510
rect 27196 37508 27252 37510
rect 26956 36474 27012 36476
rect 27036 36474 27092 36476
rect 27116 36474 27172 36476
rect 27196 36474 27252 36476
rect 26956 36422 27002 36474
rect 27002 36422 27012 36474
rect 27036 36422 27066 36474
rect 27066 36422 27078 36474
rect 27078 36422 27092 36474
rect 27116 36422 27130 36474
rect 27130 36422 27142 36474
rect 27142 36422 27172 36474
rect 27196 36422 27206 36474
rect 27206 36422 27252 36474
rect 26956 36420 27012 36422
rect 27036 36420 27092 36422
rect 27116 36420 27172 36422
rect 27196 36420 27252 36422
rect 26956 35386 27012 35388
rect 27036 35386 27092 35388
rect 27116 35386 27172 35388
rect 27196 35386 27252 35388
rect 26956 35334 27002 35386
rect 27002 35334 27012 35386
rect 27036 35334 27066 35386
rect 27066 35334 27078 35386
rect 27078 35334 27092 35386
rect 27116 35334 27130 35386
rect 27130 35334 27142 35386
rect 27142 35334 27172 35386
rect 27196 35334 27206 35386
rect 27206 35334 27252 35386
rect 26956 35332 27012 35334
rect 27036 35332 27092 35334
rect 27116 35332 27172 35334
rect 27196 35332 27252 35334
rect 26956 34298 27012 34300
rect 27036 34298 27092 34300
rect 27116 34298 27172 34300
rect 27196 34298 27252 34300
rect 26956 34246 27002 34298
rect 27002 34246 27012 34298
rect 27036 34246 27066 34298
rect 27066 34246 27078 34298
rect 27078 34246 27092 34298
rect 27116 34246 27130 34298
rect 27130 34246 27142 34298
rect 27142 34246 27172 34298
rect 27196 34246 27206 34298
rect 27206 34246 27252 34298
rect 26956 34244 27012 34246
rect 27036 34244 27092 34246
rect 27116 34244 27172 34246
rect 27196 34244 27252 34246
rect 26956 33210 27012 33212
rect 27036 33210 27092 33212
rect 27116 33210 27172 33212
rect 27196 33210 27252 33212
rect 26956 33158 27002 33210
rect 27002 33158 27012 33210
rect 27036 33158 27066 33210
rect 27066 33158 27078 33210
rect 27078 33158 27092 33210
rect 27116 33158 27130 33210
rect 27130 33158 27142 33210
rect 27142 33158 27172 33210
rect 27196 33158 27206 33210
rect 27206 33158 27252 33210
rect 26956 33156 27012 33158
rect 27036 33156 27092 33158
rect 27116 33156 27172 33158
rect 27196 33156 27252 33158
rect 26956 32122 27012 32124
rect 27036 32122 27092 32124
rect 27116 32122 27172 32124
rect 27196 32122 27252 32124
rect 26956 32070 27002 32122
rect 27002 32070 27012 32122
rect 27036 32070 27066 32122
rect 27066 32070 27078 32122
rect 27078 32070 27092 32122
rect 27116 32070 27130 32122
rect 27130 32070 27142 32122
rect 27142 32070 27172 32122
rect 27196 32070 27206 32122
rect 27206 32070 27252 32122
rect 26956 32068 27012 32070
rect 27036 32068 27092 32070
rect 27116 32068 27172 32070
rect 27196 32068 27252 32070
rect 26956 31034 27012 31036
rect 27036 31034 27092 31036
rect 27116 31034 27172 31036
rect 27196 31034 27252 31036
rect 26956 30982 27002 31034
rect 27002 30982 27012 31034
rect 27036 30982 27066 31034
rect 27066 30982 27078 31034
rect 27078 30982 27092 31034
rect 27116 30982 27130 31034
rect 27130 30982 27142 31034
rect 27142 30982 27172 31034
rect 27196 30982 27206 31034
rect 27206 30982 27252 31034
rect 26956 30980 27012 30982
rect 27036 30980 27092 30982
rect 27116 30980 27172 30982
rect 27196 30980 27252 30982
rect 26956 29946 27012 29948
rect 27036 29946 27092 29948
rect 27116 29946 27172 29948
rect 27196 29946 27252 29948
rect 26956 29894 27002 29946
rect 27002 29894 27012 29946
rect 27036 29894 27066 29946
rect 27066 29894 27078 29946
rect 27078 29894 27092 29946
rect 27116 29894 27130 29946
rect 27130 29894 27142 29946
rect 27142 29894 27172 29946
rect 27196 29894 27206 29946
rect 27206 29894 27252 29946
rect 26956 29892 27012 29894
rect 27036 29892 27092 29894
rect 27116 29892 27172 29894
rect 27196 29892 27252 29894
rect 26956 28858 27012 28860
rect 27036 28858 27092 28860
rect 27116 28858 27172 28860
rect 27196 28858 27252 28860
rect 26956 28806 27002 28858
rect 27002 28806 27012 28858
rect 27036 28806 27066 28858
rect 27066 28806 27078 28858
rect 27078 28806 27092 28858
rect 27116 28806 27130 28858
rect 27130 28806 27142 28858
rect 27142 28806 27172 28858
rect 27196 28806 27206 28858
rect 27206 28806 27252 28858
rect 26956 28804 27012 28806
rect 27036 28804 27092 28806
rect 27116 28804 27172 28806
rect 27196 28804 27252 28806
rect 26956 27770 27012 27772
rect 27036 27770 27092 27772
rect 27116 27770 27172 27772
rect 27196 27770 27252 27772
rect 26956 27718 27002 27770
rect 27002 27718 27012 27770
rect 27036 27718 27066 27770
rect 27066 27718 27078 27770
rect 27078 27718 27092 27770
rect 27116 27718 27130 27770
rect 27130 27718 27142 27770
rect 27142 27718 27172 27770
rect 27196 27718 27206 27770
rect 27206 27718 27252 27770
rect 26956 27716 27012 27718
rect 27036 27716 27092 27718
rect 27116 27716 27172 27718
rect 27196 27716 27252 27718
rect 26956 26682 27012 26684
rect 27036 26682 27092 26684
rect 27116 26682 27172 26684
rect 27196 26682 27252 26684
rect 26956 26630 27002 26682
rect 27002 26630 27012 26682
rect 27036 26630 27066 26682
rect 27066 26630 27078 26682
rect 27078 26630 27092 26682
rect 27116 26630 27130 26682
rect 27130 26630 27142 26682
rect 27142 26630 27172 26682
rect 27196 26630 27206 26682
rect 27206 26630 27252 26682
rect 26956 26628 27012 26630
rect 27036 26628 27092 26630
rect 27116 26628 27172 26630
rect 27196 26628 27252 26630
rect 26956 25594 27012 25596
rect 27036 25594 27092 25596
rect 27116 25594 27172 25596
rect 27196 25594 27252 25596
rect 26956 25542 27002 25594
rect 27002 25542 27012 25594
rect 27036 25542 27066 25594
rect 27066 25542 27078 25594
rect 27078 25542 27092 25594
rect 27116 25542 27130 25594
rect 27130 25542 27142 25594
rect 27142 25542 27172 25594
rect 27196 25542 27206 25594
rect 27206 25542 27252 25594
rect 26956 25540 27012 25542
rect 27036 25540 27092 25542
rect 27116 25540 27172 25542
rect 27196 25540 27252 25542
rect 27616 57690 27672 57692
rect 27696 57690 27752 57692
rect 27776 57690 27832 57692
rect 27856 57690 27912 57692
rect 27616 57638 27662 57690
rect 27662 57638 27672 57690
rect 27696 57638 27726 57690
rect 27726 57638 27738 57690
rect 27738 57638 27752 57690
rect 27776 57638 27790 57690
rect 27790 57638 27802 57690
rect 27802 57638 27832 57690
rect 27856 57638 27866 57690
rect 27866 57638 27912 57690
rect 27616 57636 27672 57638
rect 27696 57636 27752 57638
rect 27776 57636 27832 57638
rect 27856 57636 27912 57638
rect 27616 56602 27672 56604
rect 27696 56602 27752 56604
rect 27776 56602 27832 56604
rect 27856 56602 27912 56604
rect 27616 56550 27662 56602
rect 27662 56550 27672 56602
rect 27696 56550 27726 56602
rect 27726 56550 27738 56602
rect 27738 56550 27752 56602
rect 27776 56550 27790 56602
rect 27790 56550 27802 56602
rect 27802 56550 27832 56602
rect 27856 56550 27866 56602
rect 27866 56550 27912 56602
rect 27616 56548 27672 56550
rect 27696 56548 27752 56550
rect 27776 56548 27832 56550
rect 27856 56548 27912 56550
rect 27616 55514 27672 55516
rect 27696 55514 27752 55516
rect 27776 55514 27832 55516
rect 27856 55514 27912 55516
rect 27616 55462 27662 55514
rect 27662 55462 27672 55514
rect 27696 55462 27726 55514
rect 27726 55462 27738 55514
rect 27738 55462 27752 55514
rect 27776 55462 27790 55514
rect 27790 55462 27802 55514
rect 27802 55462 27832 55514
rect 27856 55462 27866 55514
rect 27866 55462 27912 55514
rect 27616 55460 27672 55462
rect 27696 55460 27752 55462
rect 27776 55460 27832 55462
rect 27856 55460 27912 55462
rect 27616 54426 27672 54428
rect 27696 54426 27752 54428
rect 27776 54426 27832 54428
rect 27856 54426 27912 54428
rect 27616 54374 27662 54426
rect 27662 54374 27672 54426
rect 27696 54374 27726 54426
rect 27726 54374 27738 54426
rect 27738 54374 27752 54426
rect 27776 54374 27790 54426
rect 27790 54374 27802 54426
rect 27802 54374 27832 54426
rect 27856 54374 27866 54426
rect 27866 54374 27912 54426
rect 27616 54372 27672 54374
rect 27696 54372 27752 54374
rect 27776 54372 27832 54374
rect 27856 54372 27912 54374
rect 27616 53338 27672 53340
rect 27696 53338 27752 53340
rect 27776 53338 27832 53340
rect 27856 53338 27912 53340
rect 27616 53286 27662 53338
rect 27662 53286 27672 53338
rect 27696 53286 27726 53338
rect 27726 53286 27738 53338
rect 27738 53286 27752 53338
rect 27776 53286 27790 53338
rect 27790 53286 27802 53338
rect 27802 53286 27832 53338
rect 27856 53286 27866 53338
rect 27866 53286 27912 53338
rect 27616 53284 27672 53286
rect 27696 53284 27752 53286
rect 27776 53284 27832 53286
rect 27856 53284 27912 53286
rect 27616 52250 27672 52252
rect 27696 52250 27752 52252
rect 27776 52250 27832 52252
rect 27856 52250 27912 52252
rect 27616 52198 27662 52250
rect 27662 52198 27672 52250
rect 27696 52198 27726 52250
rect 27726 52198 27738 52250
rect 27738 52198 27752 52250
rect 27776 52198 27790 52250
rect 27790 52198 27802 52250
rect 27802 52198 27832 52250
rect 27856 52198 27866 52250
rect 27866 52198 27912 52250
rect 27616 52196 27672 52198
rect 27696 52196 27752 52198
rect 27776 52196 27832 52198
rect 27856 52196 27912 52198
rect 27616 51162 27672 51164
rect 27696 51162 27752 51164
rect 27776 51162 27832 51164
rect 27856 51162 27912 51164
rect 27616 51110 27662 51162
rect 27662 51110 27672 51162
rect 27696 51110 27726 51162
rect 27726 51110 27738 51162
rect 27738 51110 27752 51162
rect 27776 51110 27790 51162
rect 27790 51110 27802 51162
rect 27802 51110 27832 51162
rect 27856 51110 27866 51162
rect 27866 51110 27912 51162
rect 27616 51108 27672 51110
rect 27696 51108 27752 51110
rect 27776 51108 27832 51110
rect 27856 51108 27912 51110
rect 27616 50074 27672 50076
rect 27696 50074 27752 50076
rect 27776 50074 27832 50076
rect 27856 50074 27912 50076
rect 27616 50022 27662 50074
rect 27662 50022 27672 50074
rect 27696 50022 27726 50074
rect 27726 50022 27738 50074
rect 27738 50022 27752 50074
rect 27776 50022 27790 50074
rect 27790 50022 27802 50074
rect 27802 50022 27832 50074
rect 27856 50022 27866 50074
rect 27866 50022 27912 50074
rect 27616 50020 27672 50022
rect 27696 50020 27752 50022
rect 27776 50020 27832 50022
rect 27856 50020 27912 50022
rect 27616 48986 27672 48988
rect 27696 48986 27752 48988
rect 27776 48986 27832 48988
rect 27856 48986 27912 48988
rect 27616 48934 27662 48986
rect 27662 48934 27672 48986
rect 27696 48934 27726 48986
rect 27726 48934 27738 48986
rect 27738 48934 27752 48986
rect 27776 48934 27790 48986
rect 27790 48934 27802 48986
rect 27802 48934 27832 48986
rect 27856 48934 27866 48986
rect 27866 48934 27912 48986
rect 27616 48932 27672 48934
rect 27696 48932 27752 48934
rect 27776 48932 27832 48934
rect 27856 48932 27912 48934
rect 27616 47898 27672 47900
rect 27696 47898 27752 47900
rect 27776 47898 27832 47900
rect 27856 47898 27912 47900
rect 27616 47846 27662 47898
rect 27662 47846 27672 47898
rect 27696 47846 27726 47898
rect 27726 47846 27738 47898
rect 27738 47846 27752 47898
rect 27776 47846 27790 47898
rect 27790 47846 27802 47898
rect 27802 47846 27832 47898
rect 27856 47846 27866 47898
rect 27866 47846 27912 47898
rect 27616 47844 27672 47846
rect 27696 47844 27752 47846
rect 27776 47844 27832 47846
rect 27856 47844 27912 47846
rect 27616 46810 27672 46812
rect 27696 46810 27752 46812
rect 27776 46810 27832 46812
rect 27856 46810 27912 46812
rect 27616 46758 27662 46810
rect 27662 46758 27672 46810
rect 27696 46758 27726 46810
rect 27726 46758 27738 46810
rect 27738 46758 27752 46810
rect 27776 46758 27790 46810
rect 27790 46758 27802 46810
rect 27802 46758 27832 46810
rect 27856 46758 27866 46810
rect 27866 46758 27912 46810
rect 27616 46756 27672 46758
rect 27696 46756 27752 46758
rect 27776 46756 27832 46758
rect 27856 46756 27912 46758
rect 27616 45722 27672 45724
rect 27696 45722 27752 45724
rect 27776 45722 27832 45724
rect 27856 45722 27912 45724
rect 27616 45670 27662 45722
rect 27662 45670 27672 45722
rect 27696 45670 27726 45722
rect 27726 45670 27738 45722
rect 27738 45670 27752 45722
rect 27776 45670 27790 45722
rect 27790 45670 27802 45722
rect 27802 45670 27832 45722
rect 27856 45670 27866 45722
rect 27866 45670 27912 45722
rect 27616 45668 27672 45670
rect 27696 45668 27752 45670
rect 27776 45668 27832 45670
rect 27856 45668 27912 45670
rect 27616 44634 27672 44636
rect 27696 44634 27752 44636
rect 27776 44634 27832 44636
rect 27856 44634 27912 44636
rect 27616 44582 27662 44634
rect 27662 44582 27672 44634
rect 27696 44582 27726 44634
rect 27726 44582 27738 44634
rect 27738 44582 27752 44634
rect 27776 44582 27790 44634
rect 27790 44582 27802 44634
rect 27802 44582 27832 44634
rect 27856 44582 27866 44634
rect 27866 44582 27912 44634
rect 27616 44580 27672 44582
rect 27696 44580 27752 44582
rect 27776 44580 27832 44582
rect 27856 44580 27912 44582
rect 27616 43546 27672 43548
rect 27696 43546 27752 43548
rect 27776 43546 27832 43548
rect 27856 43546 27912 43548
rect 27616 43494 27662 43546
rect 27662 43494 27672 43546
rect 27696 43494 27726 43546
rect 27726 43494 27738 43546
rect 27738 43494 27752 43546
rect 27776 43494 27790 43546
rect 27790 43494 27802 43546
rect 27802 43494 27832 43546
rect 27856 43494 27866 43546
rect 27866 43494 27912 43546
rect 27616 43492 27672 43494
rect 27696 43492 27752 43494
rect 27776 43492 27832 43494
rect 27856 43492 27912 43494
rect 27616 42458 27672 42460
rect 27696 42458 27752 42460
rect 27776 42458 27832 42460
rect 27856 42458 27912 42460
rect 27616 42406 27662 42458
rect 27662 42406 27672 42458
rect 27696 42406 27726 42458
rect 27726 42406 27738 42458
rect 27738 42406 27752 42458
rect 27776 42406 27790 42458
rect 27790 42406 27802 42458
rect 27802 42406 27832 42458
rect 27856 42406 27866 42458
rect 27866 42406 27912 42458
rect 27616 42404 27672 42406
rect 27696 42404 27752 42406
rect 27776 42404 27832 42406
rect 27856 42404 27912 42406
rect 27616 41370 27672 41372
rect 27696 41370 27752 41372
rect 27776 41370 27832 41372
rect 27856 41370 27912 41372
rect 27616 41318 27662 41370
rect 27662 41318 27672 41370
rect 27696 41318 27726 41370
rect 27726 41318 27738 41370
rect 27738 41318 27752 41370
rect 27776 41318 27790 41370
rect 27790 41318 27802 41370
rect 27802 41318 27832 41370
rect 27856 41318 27866 41370
rect 27866 41318 27912 41370
rect 27616 41316 27672 41318
rect 27696 41316 27752 41318
rect 27776 41316 27832 41318
rect 27856 41316 27912 41318
rect 27616 40282 27672 40284
rect 27696 40282 27752 40284
rect 27776 40282 27832 40284
rect 27856 40282 27912 40284
rect 27616 40230 27662 40282
rect 27662 40230 27672 40282
rect 27696 40230 27726 40282
rect 27726 40230 27738 40282
rect 27738 40230 27752 40282
rect 27776 40230 27790 40282
rect 27790 40230 27802 40282
rect 27802 40230 27832 40282
rect 27856 40230 27866 40282
rect 27866 40230 27912 40282
rect 27616 40228 27672 40230
rect 27696 40228 27752 40230
rect 27776 40228 27832 40230
rect 27856 40228 27912 40230
rect 27616 39194 27672 39196
rect 27696 39194 27752 39196
rect 27776 39194 27832 39196
rect 27856 39194 27912 39196
rect 27616 39142 27662 39194
rect 27662 39142 27672 39194
rect 27696 39142 27726 39194
rect 27726 39142 27738 39194
rect 27738 39142 27752 39194
rect 27776 39142 27790 39194
rect 27790 39142 27802 39194
rect 27802 39142 27832 39194
rect 27856 39142 27866 39194
rect 27866 39142 27912 39194
rect 27616 39140 27672 39142
rect 27696 39140 27752 39142
rect 27776 39140 27832 39142
rect 27856 39140 27912 39142
rect 27616 38106 27672 38108
rect 27696 38106 27752 38108
rect 27776 38106 27832 38108
rect 27856 38106 27912 38108
rect 27616 38054 27662 38106
rect 27662 38054 27672 38106
rect 27696 38054 27726 38106
rect 27726 38054 27738 38106
rect 27738 38054 27752 38106
rect 27776 38054 27790 38106
rect 27790 38054 27802 38106
rect 27802 38054 27832 38106
rect 27856 38054 27866 38106
rect 27866 38054 27912 38106
rect 27616 38052 27672 38054
rect 27696 38052 27752 38054
rect 27776 38052 27832 38054
rect 27856 38052 27912 38054
rect 27616 37018 27672 37020
rect 27696 37018 27752 37020
rect 27776 37018 27832 37020
rect 27856 37018 27912 37020
rect 27616 36966 27662 37018
rect 27662 36966 27672 37018
rect 27696 36966 27726 37018
rect 27726 36966 27738 37018
rect 27738 36966 27752 37018
rect 27776 36966 27790 37018
rect 27790 36966 27802 37018
rect 27802 36966 27832 37018
rect 27856 36966 27866 37018
rect 27866 36966 27912 37018
rect 27616 36964 27672 36966
rect 27696 36964 27752 36966
rect 27776 36964 27832 36966
rect 27856 36964 27912 36966
rect 27616 35930 27672 35932
rect 27696 35930 27752 35932
rect 27776 35930 27832 35932
rect 27856 35930 27912 35932
rect 27616 35878 27662 35930
rect 27662 35878 27672 35930
rect 27696 35878 27726 35930
rect 27726 35878 27738 35930
rect 27738 35878 27752 35930
rect 27776 35878 27790 35930
rect 27790 35878 27802 35930
rect 27802 35878 27832 35930
rect 27856 35878 27866 35930
rect 27866 35878 27912 35930
rect 27616 35876 27672 35878
rect 27696 35876 27752 35878
rect 27776 35876 27832 35878
rect 27856 35876 27912 35878
rect 27616 34842 27672 34844
rect 27696 34842 27752 34844
rect 27776 34842 27832 34844
rect 27856 34842 27912 34844
rect 27616 34790 27662 34842
rect 27662 34790 27672 34842
rect 27696 34790 27726 34842
rect 27726 34790 27738 34842
rect 27738 34790 27752 34842
rect 27776 34790 27790 34842
rect 27790 34790 27802 34842
rect 27802 34790 27832 34842
rect 27856 34790 27866 34842
rect 27866 34790 27912 34842
rect 27616 34788 27672 34790
rect 27696 34788 27752 34790
rect 27776 34788 27832 34790
rect 27856 34788 27912 34790
rect 27616 33754 27672 33756
rect 27696 33754 27752 33756
rect 27776 33754 27832 33756
rect 27856 33754 27912 33756
rect 27616 33702 27662 33754
rect 27662 33702 27672 33754
rect 27696 33702 27726 33754
rect 27726 33702 27738 33754
rect 27738 33702 27752 33754
rect 27776 33702 27790 33754
rect 27790 33702 27802 33754
rect 27802 33702 27832 33754
rect 27856 33702 27866 33754
rect 27866 33702 27912 33754
rect 27616 33700 27672 33702
rect 27696 33700 27752 33702
rect 27776 33700 27832 33702
rect 27856 33700 27912 33702
rect 27616 32666 27672 32668
rect 27696 32666 27752 32668
rect 27776 32666 27832 32668
rect 27856 32666 27912 32668
rect 27616 32614 27662 32666
rect 27662 32614 27672 32666
rect 27696 32614 27726 32666
rect 27726 32614 27738 32666
rect 27738 32614 27752 32666
rect 27776 32614 27790 32666
rect 27790 32614 27802 32666
rect 27802 32614 27832 32666
rect 27856 32614 27866 32666
rect 27866 32614 27912 32666
rect 27616 32612 27672 32614
rect 27696 32612 27752 32614
rect 27776 32612 27832 32614
rect 27856 32612 27912 32614
rect 27616 31578 27672 31580
rect 27696 31578 27752 31580
rect 27776 31578 27832 31580
rect 27856 31578 27912 31580
rect 27616 31526 27662 31578
rect 27662 31526 27672 31578
rect 27696 31526 27726 31578
rect 27726 31526 27738 31578
rect 27738 31526 27752 31578
rect 27776 31526 27790 31578
rect 27790 31526 27802 31578
rect 27802 31526 27832 31578
rect 27856 31526 27866 31578
rect 27866 31526 27912 31578
rect 27616 31524 27672 31526
rect 27696 31524 27752 31526
rect 27776 31524 27832 31526
rect 27856 31524 27912 31526
rect 27616 30490 27672 30492
rect 27696 30490 27752 30492
rect 27776 30490 27832 30492
rect 27856 30490 27912 30492
rect 27616 30438 27662 30490
rect 27662 30438 27672 30490
rect 27696 30438 27726 30490
rect 27726 30438 27738 30490
rect 27738 30438 27752 30490
rect 27776 30438 27790 30490
rect 27790 30438 27802 30490
rect 27802 30438 27832 30490
rect 27856 30438 27866 30490
rect 27866 30438 27912 30490
rect 27616 30436 27672 30438
rect 27696 30436 27752 30438
rect 27776 30436 27832 30438
rect 27856 30436 27912 30438
rect 27616 29402 27672 29404
rect 27696 29402 27752 29404
rect 27776 29402 27832 29404
rect 27856 29402 27912 29404
rect 27616 29350 27662 29402
rect 27662 29350 27672 29402
rect 27696 29350 27726 29402
rect 27726 29350 27738 29402
rect 27738 29350 27752 29402
rect 27776 29350 27790 29402
rect 27790 29350 27802 29402
rect 27802 29350 27832 29402
rect 27856 29350 27866 29402
rect 27866 29350 27912 29402
rect 27616 29348 27672 29350
rect 27696 29348 27752 29350
rect 27776 29348 27832 29350
rect 27856 29348 27912 29350
rect 27616 28314 27672 28316
rect 27696 28314 27752 28316
rect 27776 28314 27832 28316
rect 27856 28314 27912 28316
rect 27616 28262 27662 28314
rect 27662 28262 27672 28314
rect 27696 28262 27726 28314
rect 27726 28262 27738 28314
rect 27738 28262 27752 28314
rect 27776 28262 27790 28314
rect 27790 28262 27802 28314
rect 27802 28262 27832 28314
rect 27856 28262 27866 28314
rect 27866 28262 27912 28314
rect 27616 28260 27672 28262
rect 27696 28260 27752 28262
rect 27776 28260 27832 28262
rect 27856 28260 27912 28262
rect 27616 27226 27672 27228
rect 27696 27226 27752 27228
rect 27776 27226 27832 27228
rect 27856 27226 27912 27228
rect 27616 27174 27662 27226
rect 27662 27174 27672 27226
rect 27696 27174 27726 27226
rect 27726 27174 27738 27226
rect 27738 27174 27752 27226
rect 27776 27174 27790 27226
rect 27790 27174 27802 27226
rect 27802 27174 27832 27226
rect 27856 27174 27866 27226
rect 27866 27174 27912 27226
rect 27616 27172 27672 27174
rect 27696 27172 27752 27174
rect 27776 27172 27832 27174
rect 27856 27172 27912 27174
rect 27616 26138 27672 26140
rect 27696 26138 27752 26140
rect 27776 26138 27832 26140
rect 27856 26138 27912 26140
rect 27616 26086 27662 26138
rect 27662 26086 27672 26138
rect 27696 26086 27726 26138
rect 27726 26086 27738 26138
rect 27738 26086 27752 26138
rect 27776 26086 27790 26138
rect 27790 26086 27802 26138
rect 27802 26086 27832 26138
rect 27856 26086 27866 26138
rect 27866 26086 27912 26138
rect 27616 26084 27672 26086
rect 27696 26084 27752 26086
rect 27776 26084 27832 26086
rect 27856 26084 27912 26086
rect 27616 25050 27672 25052
rect 27696 25050 27752 25052
rect 27776 25050 27832 25052
rect 27856 25050 27912 25052
rect 27616 24998 27662 25050
rect 27662 24998 27672 25050
rect 27696 24998 27726 25050
rect 27726 24998 27738 25050
rect 27738 24998 27752 25050
rect 27776 24998 27790 25050
rect 27790 24998 27802 25050
rect 27802 24998 27832 25050
rect 27856 24998 27866 25050
rect 27866 24998 27912 25050
rect 27616 24996 27672 24998
rect 27696 24996 27752 24998
rect 27776 24996 27832 24998
rect 27856 24996 27912 24998
rect 26956 24506 27012 24508
rect 27036 24506 27092 24508
rect 27116 24506 27172 24508
rect 27196 24506 27252 24508
rect 26956 24454 27002 24506
rect 27002 24454 27012 24506
rect 27036 24454 27066 24506
rect 27066 24454 27078 24506
rect 27078 24454 27092 24506
rect 27116 24454 27130 24506
rect 27130 24454 27142 24506
rect 27142 24454 27172 24506
rect 27196 24454 27206 24506
rect 27206 24454 27252 24506
rect 26956 24452 27012 24454
rect 27036 24452 27092 24454
rect 27116 24452 27172 24454
rect 27196 24452 27252 24454
rect 26956 23418 27012 23420
rect 27036 23418 27092 23420
rect 27116 23418 27172 23420
rect 27196 23418 27252 23420
rect 26956 23366 27002 23418
rect 27002 23366 27012 23418
rect 27036 23366 27066 23418
rect 27066 23366 27078 23418
rect 27078 23366 27092 23418
rect 27116 23366 27130 23418
rect 27130 23366 27142 23418
rect 27142 23366 27172 23418
rect 27196 23366 27206 23418
rect 27206 23366 27252 23418
rect 26956 23364 27012 23366
rect 27036 23364 27092 23366
rect 27116 23364 27172 23366
rect 27196 23364 27252 23366
rect 26956 22330 27012 22332
rect 27036 22330 27092 22332
rect 27116 22330 27172 22332
rect 27196 22330 27252 22332
rect 26956 22278 27002 22330
rect 27002 22278 27012 22330
rect 27036 22278 27066 22330
rect 27066 22278 27078 22330
rect 27078 22278 27092 22330
rect 27116 22278 27130 22330
rect 27130 22278 27142 22330
rect 27142 22278 27172 22330
rect 27196 22278 27206 22330
rect 27206 22278 27252 22330
rect 26956 22276 27012 22278
rect 27036 22276 27092 22278
rect 27116 22276 27172 22278
rect 27196 22276 27252 22278
rect 26956 21242 27012 21244
rect 27036 21242 27092 21244
rect 27116 21242 27172 21244
rect 27196 21242 27252 21244
rect 26956 21190 27002 21242
rect 27002 21190 27012 21242
rect 27036 21190 27066 21242
rect 27066 21190 27078 21242
rect 27078 21190 27092 21242
rect 27116 21190 27130 21242
rect 27130 21190 27142 21242
rect 27142 21190 27172 21242
rect 27196 21190 27206 21242
rect 27206 21190 27252 21242
rect 26956 21188 27012 21190
rect 27036 21188 27092 21190
rect 27116 21188 27172 21190
rect 27196 21188 27252 21190
rect 27616 23962 27672 23964
rect 27696 23962 27752 23964
rect 27776 23962 27832 23964
rect 27856 23962 27912 23964
rect 27616 23910 27662 23962
rect 27662 23910 27672 23962
rect 27696 23910 27726 23962
rect 27726 23910 27738 23962
rect 27738 23910 27752 23962
rect 27776 23910 27790 23962
rect 27790 23910 27802 23962
rect 27802 23910 27832 23962
rect 27856 23910 27866 23962
rect 27866 23910 27912 23962
rect 27616 23908 27672 23910
rect 27696 23908 27752 23910
rect 27776 23908 27832 23910
rect 27856 23908 27912 23910
rect 27616 22874 27672 22876
rect 27696 22874 27752 22876
rect 27776 22874 27832 22876
rect 27856 22874 27912 22876
rect 27616 22822 27662 22874
rect 27662 22822 27672 22874
rect 27696 22822 27726 22874
rect 27726 22822 27738 22874
rect 27738 22822 27752 22874
rect 27776 22822 27790 22874
rect 27790 22822 27802 22874
rect 27802 22822 27832 22874
rect 27856 22822 27866 22874
rect 27866 22822 27912 22874
rect 27616 22820 27672 22822
rect 27696 22820 27752 22822
rect 27776 22820 27832 22822
rect 27856 22820 27912 22822
rect 27616 21786 27672 21788
rect 27696 21786 27752 21788
rect 27776 21786 27832 21788
rect 27856 21786 27912 21788
rect 27616 21734 27662 21786
rect 27662 21734 27672 21786
rect 27696 21734 27726 21786
rect 27726 21734 27738 21786
rect 27738 21734 27752 21786
rect 27776 21734 27790 21786
rect 27790 21734 27802 21786
rect 27802 21734 27832 21786
rect 27856 21734 27866 21786
rect 27866 21734 27912 21786
rect 27616 21732 27672 21734
rect 27696 21732 27752 21734
rect 27776 21732 27832 21734
rect 27856 21732 27912 21734
rect 27616 20698 27672 20700
rect 27696 20698 27752 20700
rect 27776 20698 27832 20700
rect 27856 20698 27912 20700
rect 27616 20646 27662 20698
rect 27662 20646 27672 20698
rect 27696 20646 27726 20698
rect 27726 20646 27738 20698
rect 27738 20646 27752 20698
rect 27776 20646 27790 20698
rect 27790 20646 27802 20698
rect 27802 20646 27832 20698
rect 27856 20646 27866 20698
rect 27866 20646 27912 20698
rect 27616 20644 27672 20646
rect 27696 20644 27752 20646
rect 27776 20644 27832 20646
rect 27856 20644 27912 20646
rect 26956 20154 27012 20156
rect 27036 20154 27092 20156
rect 27116 20154 27172 20156
rect 27196 20154 27252 20156
rect 26956 20102 27002 20154
rect 27002 20102 27012 20154
rect 27036 20102 27066 20154
rect 27066 20102 27078 20154
rect 27078 20102 27092 20154
rect 27116 20102 27130 20154
rect 27130 20102 27142 20154
rect 27142 20102 27172 20154
rect 27196 20102 27206 20154
rect 27206 20102 27252 20154
rect 26956 20100 27012 20102
rect 27036 20100 27092 20102
rect 27116 20100 27172 20102
rect 27196 20100 27252 20102
rect 26956 19066 27012 19068
rect 27036 19066 27092 19068
rect 27116 19066 27172 19068
rect 27196 19066 27252 19068
rect 26956 19014 27002 19066
rect 27002 19014 27012 19066
rect 27036 19014 27066 19066
rect 27066 19014 27078 19066
rect 27078 19014 27092 19066
rect 27116 19014 27130 19066
rect 27130 19014 27142 19066
rect 27142 19014 27172 19066
rect 27196 19014 27206 19066
rect 27206 19014 27252 19066
rect 26956 19012 27012 19014
rect 27036 19012 27092 19014
rect 27116 19012 27172 19014
rect 27196 19012 27252 19014
rect 26956 17978 27012 17980
rect 27036 17978 27092 17980
rect 27116 17978 27172 17980
rect 27196 17978 27252 17980
rect 26956 17926 27002 17978
rect 27002 17926 27012 17978
rect 27036 17926 27066 17978
rect 27066 17926 27078 17978
rect 27078 17926 27092 17978
rect 27116 17926 27130 17978
rect 27130 17926 27142 17978
rect 27142 17926 27172 17978
rect 27196 17926 27206 17978
rect 27206 17926 27252 17978
rect 26956 17924 27012 17926
rect 27036 17924 27092 17926
rect 27116 17924 27172 17926
rect 27196 17924 27252 17926
rect 26956 16890 27012 16892
rect 27036 16890 27092 16892
rect 27116 16890 27172 16892
rect 27196 16890 27252 16892
rect 26956 16838 27002 16890
rect 27002 16838 27012 16890
rect 27036 16838 27066 16890
rect 27066 16838 27078 16890
rect 27078 16838 27092 16890
rect 27116 16838 27130 16890
rect 27130 16838 27142 16890
rect 27142 16838 27172 16890
rect 27196 16838 27206 16890
rect 27206 16838 27252 16890
rect 26956 16836 27012 16838
rect 27036 16836 27092 16838
rect 27116 16836 27172 16838
rect 27196 16836 27252 16838
rect 26956 15802 27012 15804
rect 27036 15802 27092 15804
rect 27116 15802 27172 15804
rect 27196 15802 27252 15804
rect 26956 15750 27002 15802
rect 27002 15750 27012 15802
rect 27036 15750 27066 15802
rect 27066 15750 27078 15802
rect 27078 15750 27092 15802
rect 27116 15750 27130 15802
rect 27130 15750 27142 15802
rect 27142 15750 27172 15802
rect 27196 15750 27206 15802
rect 27206 15750 27252 15802
rect 26956 15748 27012 15750
rect 27036 15748 27092 15750
rect 27116 15748 27172 15750
rect 27196 15748 27252 15750
rect 26956 14714 27012 14716
rect 27036 14714 27092 14716
rect 27116 14714 27172 14716
rect 27196 14714 27252 14716
rect 26956 14662 27002 14714
rect 27002 14662 27012 14714
rect 27036 14662 27066 14714
rect 27066 14662 27078 14714
rect 27078 14662 27092 14714
rect 27116 14662 27130 14714
rect 27130 14662 27142 14714
rect 27142 14662 27172 14714
rect 27196 14662 27206 14714
rect 27206 14662 27252 14714
rect 26956 14660 27012 14662
rect 27036 14660 27092 14662
rect 27116 14660 27172 14662
rect 27196 14660 27252 14662
rect 26956 13626 27012 13628
rect 27036 13626 27092 13628
rect 27116 13626 27172 13628
rect 27196 13626 27252 13628
rect 26956 13574 27002 13626
rect 27002 13574 27012 13626
rect 27036 13574 27066 13626
rect 27066 13574 27078 13626
rect 27078 13574 27092 13626
rect 27116 13574 27130 13626
rect 27130 13574 27142 13626
rect 27142 13574 27172 13626
rect 27196 13574 27206 13626
rect 27206 13574 27252 13626
rect 26956 13572 27012 13574
rect 27036 13572 27092 13574
rect 27116 13572 27172 13574
rect 27196 13572 27252 13574
rect 26956 12538 27012 12540
rect 27036 12538 27092 12540
rect 27116 12538 27172 12540
rect 27196 12538 27252 12540
rect 26956 12486 27002 12538
rect 27002 12486 27012 12538
rect 27036 12486 27066 12538
rect 27066 12486 27078 12538
rect 27078 12486 27092 12538
rect 27116 12486 27130 12538
rect 27130 12486 27142 12538
rect 27142 12486 27172 12538
rect 27196 12486 27206 12538
rect 27206 12486 27252 12538
rect 26956 12484 27012 12486
rect 27036 12484 27092 12486
rect 27116 12484 27172 12486
rect 27196 12484 27252 12486
rect 26956 11450 27012 11452
rect 27036 11450 27092 11452
rect 27116 11450 27172 11452
rect 27196 11450 27252 11452
rect 26956 11398 27002 11450
rect 27002 11398 27012 11450
rect 27036 11398 27066 11450
rect 27066 11398 27078 11450
rect 27078 11398 27092 11450
rect 27116 11398 27130 11450
rect 27130 11398 27142 11450
rect 27142 11398 27172 11450
rect 27196 11398 27206 11450
rect 27206 11398 27252 11450
rect 26956 11396 27012 11398
rect 27036 11396 27092 11398
rect 27116 11396 27172 11398
rect 27196 11396 27252 11398
rect 26956 10362 27012 10364
rect 27036 10362 27092 10364
rect 27116 10362 27172 10364
rect 27196 10362 27252 10364
rect 26956 10310 27002 10362
rect 27002 10310 27012 10362
rect 27036 10310 27066 10362
rect 27066 10310 27078 10362
rect 27078 10310 27092 10362
rect 27116 10310 27130 10362
rect 27130 10310 27142 10362
rect 27142 10310 27172 10362
rect 27196 10310 27206 10362
rect 27206 10310 27252 10362
rect 26956 10308 27012 10310
rect 27036 10308 27092 10310
rect 27116 10308 27172 10310
rect 27196 10308 27252 10310
rect 26956 9274 27012 9276
rect 27036 9274 27092 9276
rect 27116 9274 27172 9276
rect 27196 9274 27252 9276
rect 26956 9222 27002 9274
rect 27002 9222 27012 9274
rect 27036 9222 27066 9274
rect 27066 9222 27078 9274
rect 27078 9222 27092 9274
rect 27116 9222 27130 9274
rect 27130 9222 27142 9274
rect 27142 9222 27172 9274
rect 27196 9222 27206 9274
rect 27206 9222 27252 9274
rect 26956 9220 27012 9222
rect 27036 9220 27092 9222
rect 27116 9220 27172 9222
rect 27196 9220 27252 9222
rect 27616 19610 27672 19612
rect 27696 19610 27752 19612
rect 27776 19610 27832 19612
rect 27856 19610 27912 19612
rect 27616 19558 27662 19610
rect 27662 19558 27672 19610
rect 27696 19558 27726 19610
rect 27726 19558 27738 19610
rect 27738 19558 27752 19610
rect 27776 19558 27790 19610
rect 27790 19558 27802 19610
rect 27802 19558 27832 19610
rect 27856 19558 27866 19610
rect 27866 19558 27912 19610
rect 27616 19556 27672 19558
rect 27696 19556 27752 19558
rect 27776 19556 27832 19558
rect 27856 19556 27912 19558
rect 27616 18522 27672 18524
rect 27696 18522 27752 18524
rect 27776 18522 27832 18524
rect 27856 18522 27912 18524
rect 27616 18470 27662 18522
rect 27662 18470 27672 18522
rect 27696 18470 27726 18522
rect 27726 18470 27738 18522
rect 27738 18470 27752 18522
rect 27776 18470 27790 18522
rect 27790 18470 27802 18522
rect 27802 18470 27832 18522
rect 27856 18470 27866 18522
rect 27866 18470 27912 18522
rect 27616 18468 27672 18470
rect 27696 18468 27752 18470
rect 27776 18468 27832 18470
rect 27856 18468 27912 18470
rect 27616 17434 27672 17436
rect 27696 17434 27752 17436
rect 27776 17434 27832 17436
rect 27856 17434 27912 17436
rect 27616 17382 27662 17434
rect 27662 17382 27672 17434
rect 27696 17382 27726 17434
rect 27726 17382 27738 17434
rect 27738 17382 27752 17434
rect 27776 17382 27790 17434
rect 27790 17382 27802 17434
rect 27802 17382 27832 17434
rect 27856 17382 27866 17434
rect 27866 17382 27912 17434
rect 27616 17380 27672 17382
rect 27696 17380 27752 17382
rect 27776 17380 27832 17382
rect 27856 17380 27912 17382
rect 29090 38956 29146 38992
rect 29090 38936 29092 38956
rect 29092 38936 29144 38956
rect 29144 38936 29146 38956
rect 28998 38664 29054 38720
rect 29366 38936 29422 38992
rect 29550 38664 29606 38720
rect 27616 16346 27672 16348
rect 27696 16346 27752 16348
rect 27776 16346 27832 16348
rect 27856 16346 27912 16348
rect 27616 16294 27662 16346
rect 27662 16294 27672 16346
rect 27696 16294 27726 16346
rect 27726 16294 27738 16346
rect 27738 16294 27752 16346
rect 27776 16294 27790 16346
rect 27790 16294 27802 16346
rect 27802 16294 27832 16346
rect 27856 16294 27866 16346
rect 27866 16294 27912 16346
rect 27616 16292 27672 16294
rect 27696 16292 27752 16294
rect 27776 16292 27832 16294
rect 27856 16292 27912 16294
rect 27616 15258 27672 15260
rect 27696 15258 27752 15260
rect 27776 15258 27832 15260
rect 27856 15258 27912 15260
rect 27616 15206 27662 15258
rect 27662 15206 27672 15258
rect 27696 15206 27726 15258
rect 27726 15206 27738 15258
rect 27738 15206 27752 15258
rect 27776 15206 27790 15258
rect 27790 15206 27802 15258
rect 27802 15206 27832 15258
rect 27856 15206 27866 15258
rect 27866 15206 27912 15258
rect 27616 15204 27672 15206
rect 27696 15204 27752 15206
rect 27776 15204 27832 15206
rect 27856 15204 27912 15206
rect 27616 14170 27672 14172
rect 27696 14170 27752 14172
rect 27776 14170 27832 14172
rect 27856 14170 27912 14172
rect 27616 14118 27662 14170
rect 27662 14118 27672 14170
rect 27696 14118 27726 14170
rect 27726 14118 27738 14170
rect 27738 14118 27752 14170
rect 27776 14118 27790 14170
rect 27790 14118 27802 14170
rect 27802 14118 27832 14170
rect 27856 14118 27866 14170
rect 27866 14118 27912 14170
rect 27616 14116 27672 14118
rect 27696 14116 27752 14118
rect 27776 14116 27832 14118
rect 27856 14116 27912 14118
rect 27616 13082 27672 13084
rect 27696 13082 27752 13084
rect 27776 13082 27832 13084
rect 27856 13082 27912 13084
rect 27616 13030 27662 13082
rect 27662 13030 27672 13082
rect 27696 13030 27726 13082
rect 27726 13030 27738 13082
rect 27738 13030 27752 13082
rect 27776 13030 27790 13082
rect 27790 13030 27802 13082
rect 27802 13030 27832 13082
rect 27856 13030 27866 13082
rect 27866 13030 27912 13082
rect 27616 13028 27672 13030
rect 27696 13028 27752 13030
rect 27776 13028 27832 13030
rect 27856 13028 27912 13030
rect 27616 11994 27672 11996
rect 27696 11994 27752 11996
rect 27776 11994 27832 11996
rect 27856 11994 27912 11996
rect 27616 11942 27662 11994
rect 27662 11942 27672 11994
rect 27696 11942 27726 11994
rect 27726 11942 27738 11994
rect 27738 11942 27752 11994
rect 27776 11942 27790 11994
rect 27790 11942 27802 11994
rect 27802 11942 27832 11994
rect 27856 11942 27866 11994
rect 27866 11942 27912 11994
rect 27616 11940 27672 11942
rect 27696 11940 27752 11942
rect 27776 11940 27832 11942
rect 27856 11940 27912 11942
rect 27616 10906 27672 10908
rect 27696 10906 27752 10908
rect 27776 10906 27832 10908
rect 27856 10906 27912 10908
rect 27616 10854 27662 10906
rect 27662 10854 27672 10906
rect 27696 10854 27726 10906
rect 27726 10854 27738 10906
rect 27738 10854 27752 10906
rect 27776 10854 27790 10906
rect 27790 10854 27802 10906
rect 27802 10854 27832 10906
rect 27856 10854 27866 10906
rect 27866 10854 27912 10906
rect 27616 10852 27672 10854
rect 27696 10852 27752 10854
rect 27776 10852 27832 10854
rect 27856 10852 27912 10854
rect 27616 9818 27672 9820
rect 27696 9818 27752 9820
rect 27776 9818 27832 9820
rect 27856 9818 27912 9820
rect 27616 9766 27662 9818
rect 27662 9766 27672 9818
rect 27696 9766 27726 9818
rect 27726 9766 27738 9818
rect 27738 9766 27752 9818
rect 27776 9766 27790 9818
rect 27790 9766 27802 9818
rect 27802 9766 27832 9818
rect 27856 9766 27866 9818
rect 27866 9766 27912 9818
rect 27616 9764 27672 9766
rect 27696 9764 27752 9766
rect 27776 9764 27832 9766
rect 27856 9764 27912 9766
rect 26956 8186 27012 8188
rect 27036 8186 27092 8188
rect 27116 8186 27172 8188
rect 27196 8186 27252 8188
rect 26956 8134 27002 8186
rect 27002 8134 27012 8186
rect 27036 8134 27066 8186
rect 27066 8134 27078 8186
rect 27078 8134 27092 8186
rect 27116 8134 27130 8186
rect 27130 8134 27142 8186
rect 27142 8134 27172 8186
rect 27196 8134 27206 8186
rect 27206 8134 27252 8186
rect 26956 8132 27012 8134
rect 27036 8132 27092 8134
rect 27116 8132 27172 8134
rect 27196 8132 27252 8134
rect 26956 7098 27012 7100
rect 27036 7098 27092 7100
rect 27116 7098 27172 7100
rect 27196 7098 27252 7100
rect 26956 7046 27002 7098
rect 27002 7046 27012 7098
rect 27036 7046 27066 7098
rect 27066 7046 27078 7098
rect 27078 7046 27092 7098
rect 27116 7046 27130 7098
rect 27130 7046 27142 7098
rect 27142 7046 27172 7098
rect 27196 7046 27206 7098
rect 27206 7046 27252 7098
rect 26956 7044 27012 7046
rect 27036 7044 27092 7046
rect 27116 7044 27172 7046
rect 27196 7044 27252 7046
rect 26956 6010 27012 6012
rect 27036 6010 27092 6012
rect 27116 6010 27172 6012
rect 27196 6010 27252 6012
rect 26956 5958 27002 6010
rect 27002 5958 27012 6010
rect 27036 5958 27066 6010
rect 27066 5958 27078 6010
rect 27078 5958 27092 6010
rect 27116 5958 27130 6010
rect 27130 5958 27142 6010
rect 27142 5958 27172 6010
rect 27196 5958 27206 6010
rect 27206 5958 27252 6010
rect 26956 5956 27012 5958
rect 27036 5956 27092 5958
rect 27116 5956 27172 5958
rect 27196 5956 27252 5958
rect 26956 4922 27012 4924
rect 27036 4922 27092 4924
rect 27116 4922 27172 4924
rect 27196 4922 27252 4924
rect 26956 4870 27002 4922
rect 27002 4870 27012 4922
rect 27036 4870 27066 4922
rect 27066 4870 27078 4922
rect 27078 4870 27092 4922
rect 27116 4870 27130 4922
rect 27130 4870 27142 4922
rect 27142 4870 27172 4922
rect 27196 4870 27206 4922
rect 27206 4870 27252 4922
rect 26956 4868 27012 4870
rect 27036 4868 27092 4870
rect 27116 4868 27172 4870
rect 27196 4868 27252 4870
rect 26956 3834 27012 3836
rect 27036 3834 27092 3836
rect 27116 3834 27172 3836
rect 27196 3834 27252 3836
rect 26956 3782 27002 3834
rect 27002 3782 27012 3834
rect 27036 3782 27066 3834
rect 27066 3782 27078 3834
rect 27078 3782 27092 3834
rect 27116 3782 27130 3834
rect 27130 3782 27142 3834
rect 27142 3782 27172 3834
rect 27196 3782 27206 3834
rect 27206 3782 27252 3834
rect 26956 3780 27012 3782
rect 27036 3780 27092 3782
rect 27116 3780 27172 3782
rect 27196 3780 27252 3782
rect 27616 8730 27672 8732
rect 27696 8730 27752 8732
rect 27776 8730 27832 8732
rect 27856 8730 27912 8732
rect 27616 8678 27662 8730
rect 27662 8678 27672 8730
rect 27696 8678 27726 8730
rect 27726 8678 27738 8730
rect 27738 8678 27752 8730
rect 27776 8678 27790 8730
rect 27790 8678 27802 8730
rect 27802 8678 27832 8730
rect 27856 8678 27866 8730
rect 27866 8678 27912 8730
rect 27616 8676 27672 8678
rect 27696 8676 27752 8678
rect 27776 8676 27832 8678
rect 27856 8676 27912 8678
rect 27616 7642 27672 7644
rect 27696 7642 27752 7644
rect 27776 7642 27832 7644
rect 27856 7642 27912 7644
rect 27616 7590 27662 7642
rect 27662 7590 27672 7642
rect 27696 7590 27726 7642
rect 27726 7590 27738 7642
rect 27738 7590 27752 7642
rect 27776 7590 27790 7642
rect 27790 7590 27802 7642
rect 27802 7590 27832 7642
rect 27856 7590 27866 7642
rect 27866 7590 27912 7642
rect 27616 7588 27672 7590
rect 27696 7588 27752 7590
rect 27776 7588 27832 7590
rect 27856 7588 27912 7590
rect 27616 6554 27672 6556
rect 27696 6554 27752 6556
rect 27776 6554 27832 6556
rect 27856 6554 27912 6556
rect 27616 6502 27662 6554
rect 27662 6502 27672 6554
rect 27696 6502 27726 6554
rect 27726 6502 27738 6554
rect 27738 6502 27752 6554
rect 27776 6502 27790 6554
rect 27790 6502 27802 6554
rect 27802 6502 27832 6554
rect 27856 6502 27866 6554
rect 27866 6502 27912 6554
rect 27616 6500 27672 6502
rect 27696 6500 27752 6502
rect 27776 6500 27832 6502
rect 27856 6500 27912 6502
rect 27616 5466 27672 5468
rect 27696 5466 27752 5468
rect 27776 5466 27832 5468
rect 27856 5466 27912 5468
rect 27616 5414 27662 5466
rect 27662 5414 27672 5466
rect 27696 5414 27726 5466
rect 27726 5414 27738 5466
rect 27738 5414 27752 5466
rect 27776 5414 27790 5466
rect 27790 5414 27802 5466
rect 27802 5414 27832 5466
rect 27856 5414 27866 5466
rect 27866 5414 27912 5466
rect 27616 5412 27672 5414
rect 27696 5412 27752 5414
rect 27776 5412 27832 5414
rect 27856 5412 27912 5414
rect 27616 4378 27672 4380
rect 27696 4378 27752 4380
rect 27776 4378 27832 4380
rect 27856 4378 27912 4380
rect 27616 4326 27662 4378
rect 27662 4326 27672 4378
rect 27696 4326 27726 4378
rect 27726 4326 27738 4378
rect 27738 4326 27752 4378
rect 27776 4326 27790 4378
rect 27790 4326 27802 4378
rect 27802 4326 27832 4378
rect 27856 4326 27866 4378
rect 27866 4326 27912 4378
rect 27616 4324 27672 4326
rect 27696 4324 27752 4326
rect 27776 4324 27832 4326
rect 27856 4324 27912 4326
rect 27616 3290 27672 3292
rect 27696 3290 27752 3292
rect 27776 3290 27832 3292
rect 27856 3290 27912 3292
rect 27616 3238 27662 3290
rect 27662 3238 27672 3290
rect 27696 3238 27726 3290
rect 27726 3238 27738 3290
rect 27738 3238 27752 3290
rect 27776 3238 27790 3290
rect 27790 3238 27802 3290
rect 27802 3238 27832 3290
rect 27856 3238 27866 3290
rect 27866 3238 27912 3290
rect 27616 3236 27672 3238
rect 27696 3236 27752 3238
rect 27776 3236 27832 3238
rect 27856 3236 27912 3238
rect 30562 40024 30618 40080
rect 32616 68570 32672 68572
rect 32696 68570 32752 68572
rect 32776 68570 32832 68572
rect 32856 68570 32912 68572
rect 32616 68518 32662 68570
rect 32662 68518 32672 68570
rect 32696 68518 32726 68570
rect 32726 68518 32738 68570
rect 32738 68518 32752 68570
rect 32776 68518 32790 68570
rect 32790 68518 32802 68570
rect 32802 68518 32832 68570
rect 32856 68518 32866 68570
rect 32866 68518 32912 68570
rect 32616 68516 32672 68518
rect 32696 68516 32752 68518
rect 32776 68516 32832 68518
rect 32856 68516 32912 68518
rect 31956 68026 32012 68028
rect 32036 68026 32092 68028
rect 32116 68026 32172 68028
rect 32196 68026 32252 68028
rect 31956 67974 32002 68026
rect 32002 67974 32012 68026
rect 32036 67974 32066 68026
rect 32066 67974 32078 68026
rect 32078 67974 32092 68026
rect 32116 67974 32130 68026
rect 32130 67974 32142 68026
rect 32142 67974 32172 68026
rect 32196 67974 32206 68026
rect 32206 67974 32252 68026
rect 31956 67972 32012 67974
rect 32036 67972 32092 67974
rect 32116 67972 32172 67974
rect 32196 67972 32252 67974
rect 32616 67482 32672 67484
rect 32696 67482 32752 67484
rect 32776 67482 32832 67484
rect 32856 67482 32912 67484
rect 32616 67430 32662 67482
rect 32662 67430 32672 67482
rect 32696 67430 32726 67482
rect 32726 67430 32738 67482
rect 32738 67430 32752 67482
rect 32776 67430 32790 67482
rect 32790 67430 32802 67482
rect 32802 67430 32832 67482
rect 32856 67430 32866 67482
rect 32866 67430 32912 67482
rect 32616 67428 32672 67430
rect 32696 67428 32752 67430
rect 32776 67428 32832 67430
rect 32856 67428 32912 67430
rect 31956 66938 32012 66940
rect 32036 66938 32092 66940
rect 32116 66938 32172 66940
rect 32196 66938 32252 66940
rect 31956 66886 32002 66938
rect 32002 66886 32012 66938
rect 32036 66886 32066 66938
rect 32066 66886 32078 66938
rect 32078 66886 32092 66938
rect 32116 66886 32130 66938
rect 32130 66886 32142 66938
rect 32142 66886 32172 66938
rect 32196 66886 32206 66938
rect 32206 66886 32252 66938
rect 31956 66884 32012 66886
rect 32036 66884 32092 66886
rect 32116 66884 32172 66886
rect 32196 66884 32252 66886
rect 32616 66394 32672 66396
rect 32696 66394 32752 66396
rect 32776 66394 32832 66396
rect 32856 66394 32912 66396
rect 32616 66342 32662 66394
rect 32662 66342 32672 66394
rect 32696 66342 32726 66394
rect 32726 66342 32738 66394
rect 32738 66342 32752 66394
rect 32776 66342 32790 66394
rect 32790 66342 32802 66394
rect 32802 66342 32832 66394
rect 32856 66342 32866 66394
rect 32866 66342 32912 66394
rect 32616 66340 32672 66342
rect 32696 66340 32752 66342
rect 32776 66340 32832 66342
rect 32856 66340 32912 66342
rect 31956 65850 32012 65852
rect 32036 65850 32092 65852
rect 32116 65850 32172 65852
rect 32196 65850 32252 65852
rect 31956 65798 32002 65850
rect 32002 65798 32012 65850
rect 32036 65798 32066 65850
rect 32066 65798 32078 65850
rect 32078 65798 32092 65850
rect 32116 65798 32130 65850
rect 32130 65798 32142 65850
rect 32142 65798 32172 65850
rect 32196 65798 32206 65850
rect 32206 65798 32252 65850
rect 31956 65796 32012 65798
rect 32036 65796 32092 65798
rect 32116 65796 32172 65798
rect 32196 65796 32252 65798
rect 32616 65306 32672 65308
rect 32696 65306 32752 65308
rect 32776 65306 32832 65308
rect 32856 65306 32912 65308
rect 32616 65254 32662 65306
rect 32662 65254 32672 65306
rect 32696 65254 32726 65306
rect 32726 65254 32738 65306
rect 32738 65254 32752 65306
rect 32776 65254 32790 65306
rect 32790 65254 32802 65306
rect 32802 65254 32832 65306
rect 32856 65254 32866 65306
rect 32866 65254 32912 65306
rect 32616 65252 32672 65254
rect 32696 65252 32752 65254
rect 32776 65252 32832 65254
rect 32856 65252 32912 65254
rect 31956 64762 32012 64764
rect 32036 64762 32092 64764
rect 32116 64762 32172 64764
rect 32196 64762 32252 64764
rect 31956 64710 32002 64762
rect 32002 64710 32012 64762
rect 32036 64710 32066 64762
rect 32066 64710 32078 64762
rect 32078 64710 32092 64762
rect 32116 64710 32130 64762
rect 32130 64710 32142 64762
rect 32142 64710 32172 64762
rect 32196 64710 32206 64762
rect 32206 64710 32252 64762
rect 31956 64708 32012 64710
rect 32036 64708 32092 64710
rect 32116 64708 32172 64710
rect 32196 64708 32252 64710
rect 31956 63674 32012 63676
rect 32036 63674 32092 63676
rect 32116 63674 32172 63676
rect 32196 63674 32252 63676
rect 31956 63622 32002 63674
rect 32002 63622 32012 63674
rect 32036 63622 32066 63674
rect 32066 63622 32078 63674
rect 32078 63622 32092 63674
rect 32116 63622 32130 63674
rect 32130 63622 32142 63674
rect 32142 63622 32172 63674
rect 32196 63622 32206 63674
rect 32206 63622 32252 63674
rect 31956 63620 32012 63622
rect 32036 63620 32092 63622
rect 32116 63620 32172 63622
rect 32196 63620 32252 63622
rect 31956 62586 32012 62588
rect 32036 62586 32092 62588
rect 32116 62586 32172 62588
rect 32196 62586 32252 62588
rect 31956 62534 32002 62586
rect 32002 62534 32012 62586
rect 32036 62534 32066 62586
rect 32066 62534 32078 62586
rect 32078 62534 32092 62586
rect 32116 62534 32130 62586
rect 32130 62534 32142 62586
rect 32142 62534 32172 62586
rect 32196 62534 32206 62586
rect 32206 62534 32252 62586
rect 31956 62532 32012 62534
rect 32036 62532 32092 62534
rect 32116 62532 32172 62534
rect 32196 62532 32252 62534
rect 31956 61498 32012 61500
rect 32036 61498 32092 61500
rect 32116 61498 32172 61500
rect 32196 61498 32252 61500
rect 31956 61446 32002 61498
rect 32002 61446 32012 61498
rect 32036 61446 32066 61498
rect 32066 61446 32078 61498
rect 32078 61446 32092 61498
rect 32116 61446 32130 61498
rect 32130 61446 32142 61498
rect 32142 61446 32172 61498
rect 32196 61446 32206 61498
rect 32206 61446 32252 61498
rect 31956 61444 32012 61446
rect 32036 61444 32092 61446
rect 32116 61444 32172 61446
rect 32196 61444 32252 61446
rect 31956 60410 32012 60412
rect 32036 60410 32092 60412
rect 32116 60410 32172 60412
rect 32196 60410 32252 60412
rect 31956 60358 32002 60410
rect 32002 60358 32012 60410
rect 32036 60358 32066 60410
rect 32066 60358 32078 60410
rect 32078 60358 32092 60410
rect 32116 60358 32130 60410
rect 32130 60358 32142 60410
rect 32142 60358 32172 60410
rect 32196 60358 32206 60410
rect 32206 60358 32252 60410
rect 31956 60356 32012 60358
rect 32036 60356 32092 60358
rect 32116 60356 32172 60358
rect 32196 60356 32252 60358
rect 31956 59322 32012 59324
rect 32036 59322 32092 59324
rect 32116 59322 32172 59324
rect 32196 59322 32252 59324
rect 31956 59270 32002 59322
rect 32002 59270 32012 59322
rect 32036 59270 32066 59322
rect 32066 59270 32078 59322
rect 32078 59270 32092 59322
rect 32116 59270 32130 59322
rect 32130 59270 32142 59322
rect 32142 59270 32172 59322
rect 32196 59270 32206 59322
rect 32206 59270 32252 59322
rect 31956 59268 32012 59270
rect 32036 59268 32092 59270
rect 32116 59268 32172 59270
rect 32196 59268 32252 59270
rect 31956 58234 32012 58236
rect 32036 58234 32092 58236
rect 32116 58234 32172 58236
rect 32196 58234 32252 58236
rect 31956 58182 32002 58234
rect 32002 58182 32012 58234
rect 32036 58182 32066 58234
rect 32066 58182 32078 58234
rect 32078 58182 32092 58234
rect 32116 58182 32130 58234
rect 32130 58182 32142 58234
rect 32142 58182 32172 58234
rect 32196 58182 32206 58234
rect 32206 58182 32252 58234
rect 31956 58180 32012 58182
rect 32036 58180 32092 58182
rect 32116 58180 32172 58182
rect 32196 58180 32252 58182
rect 31956 57146 32012 57148
rect 32036 57146 32092 57148
rect 32116 57146 32172 57148
rect 32196 57146 32252 57148
rect 31956 57094 32002 57146
rect 32002 57094 32012 57146
rect 32036 57094 32066 57146
rect 32066 57094 32078 57146
rect 32078 57094 32092 57146
rect 32116 57094 32130 57146
rect 32130 57094 32142 57146
rect 32142 57094 32172 57146
rect 32196 57094 32206 57146
rect 32206 57094 32252 57146
rect 31956 57092 32012 57094
rect 32036 57092 32092 57094
rect 32116 57092 32172 57094
rect 32196 57092 32252 57094
rect 31956 56058 32012 56060
rect 32036 56058 32092 56060
rect 32116 56058 32172 56060
rect 32196 56058 32252 56060
rect 31956 56006 32002 56058
rect 32002 56006 32012 56058
rect 32036 56006 32066 56058
rect 32066 56006 32078 56058
rect 32078 56006 32092 56058
rect 32116 56006 32130 56058
rect 32130 56006 32142 56058
rect 32142 56006 32172 56058
rect 32196 56006 32206 56058
rect 32206 56006 32252 56058
rect 31956 56004 32012 56006
rect 32036 56004 32092 56006
rect 32116 56004 32172 56006
rect 32196 56004 32252 56006
rect 31956 54970 32012 54972
rect 32036 54970 32092 54972
rect 32116 54970 32172 54972
rect 32196 54970 32252 54972
rect 31956 54918 32002 54970
rect 32002 54918 32012 54970
rect 32036 54918 32066 54970
rect 32066 54918 32078 54970
rect 32078 54918 32092 54970
rect 32116 54918 32130 54970
rect 32130 54918 32142 54970
rect 32142 54918 32172 54970
rect 32196 54918 32206 54970
rect 32206 54918 32252 54970
rect 31956 54916 32012 54918
rect 32036 54916 32092 54918
rect 32116 54916 32172 54918
rect 32196 54916 32252 54918
rect 31956 53882 32012 53884
rect 32036 53882 32092 53884
rect 32116 53882 32172 53884
rect 32196 53882 32252 53884
rect 31956 53830 32002 53882
rect 32002 53830 32012 53882
rect 32036 53830 32066 53882
rect 32066 53830 32078 53882
rect 32078 53830 32092 53882
rect 32116 53830 32130 53882
rect 32130 53830 32142 53882
rect 32142 53830 32172 53882
rect 32196 53830 32206 53882
rect 32206 53830 32252 53882
rect 31956 53828 32012 53830
rect 32036 53828 32092 53830
rect 32116 53828 32172 53830
rect 32196 53828 32252 53830
rect 31956 52794 32012 52796
rect 32036 52794 32092 52796
rect 32116 52794 32172 52796
rect 32196 52794 32252 52796
rect 31956 52742 32002 52794
rect 32002 52742 32012 52794
rect 32036 52742 32066 52794
rect 32066 52742 32078 52794
rect 32078 52742 32092 52794
rect 32116 52742 32130 52794
rect 32130 52742 32142 52794
rect 32142 52742 32172 52794
rect 32196 52742 32206 52794
rect 32206 52742 32252 52794
rect 31956 52740 32012 52742
rect 32036 52740 32092 52742
rect 32116 52740 32172 52742
rect 32196 52740 32252 52742
rect 31956 51706 32012 51708
rect 32036 51706 32092 51708
rect 32116 51706 32172 51708
rect 32196 51706 32252 51708
rect 31956 51654 32002 51706
rect 32002 51654 32012 51706
rect 32036 51654 32066 51706
rect 32066 51654 32078 51706
rect 32078 51654 32092 51706
rect 32116 51654 32130 51706
rect 32130 51654 32142 51706
rect 32142 51654 32172 51706
rect 32196 51654 32206 51706
rect 32206 51654 32252 51706
rect 31956 51652 32012 51654
rect 32036 51652 32092 51654
rect 32116 51652 32172 51654
rect 32196 51652 32252 51654
rect 32616 64218 32672 64220
rect 32696 64218 32752 64220
rect 32776 64218 32832 64220
rect 32856 64218 32912 64220
rect 32616 64166 32662 64218
rect 32662 64166 32672 64218
rect 32696 64166 32726 64218
rect 32726 64166 32738 64218
rect 32738 64166 32752 64218
rect 32776 64166 32790 64218
rect 32790 64166 32802 64218
rect 32802 64166 32832 64218
rect 32856 64166 32866 64218
rect 32866 64166 32912 64218
rect 32616 64164 32672 64166
rect 32696 64164 32752 64166
rect 32776 64164 32832 64166
rect 32856 64164 32912 64166
rect 32616 63130 32672 63132
rect 32696 63130 32752 63132
rect 32776 63130 32832 63132
rect 32856 63130 32912 63132
rect 32616 63078 32662 63130
rect 32662 63078 32672 63130
rect 32696 63078 32726 63130
rect 32726 63078 32738 63130
rect 32738 63078 32752 63130
rect 32776 63078 32790 63130
rect 32790 63078 32802 63130
rect 32802 63078 32832 63130
rect 32856 63078 32866 63130
rect 32866 63078 32912 63130
rect 32616 63076 32672 63078
rect 32696 63076 32752 63078
rect 32776 63076 32832 63078
rect 32856 63076 32912 63078
rect 33598 62736 33654 62792
rect 32616 62042 32672 62044
rect 32696 62042 32752 62044
rect 32776 62042 32832 62044
rect 32856 62042 32912 62044
rect 32616 61990 32662 62042
rect 32662 61990 32672 62042
rect 32696 61990 32726 62042
rect 32726 61990 32738 62042
rect 32738 61990 32752 62042
rect 32776 61990 32790 62042
rect 32790 61990 32802 62042
rect 32802 61990 32832 62042
rect 32856 61990 32866 62042
rect 32866 61990 32912 62042
rect 32616 61988 32672 61990
rect 32696 61988 32752 61990
rect 32776 61988 32832 61990
rect 32856 61988 32912 61990
rect 32616 60954 32672 60956
rect 32696 60954 32752 60956
rect 32776 60954 32832 60956
rect 32856 60954 32912 60956
rect 32616 60902 32662 60954
rect 32662 60902 32672 60954
rect 32696 60902 32726 60954
rect 32726 60902 32738 60954
rect 32738 60902 32752 60954
rect 32776 60902 32790 60954
rect 32790 60902 32802 60954
rect 32802 60902 32832 60954
rect 32856 60902 32866 60954
rect 32866 60902 32912 60954
rect 32616 60900 32672 60902
rect 32696 60900 32752 60902
rect 32776 60900 32832 60902
rect 32856 60900 32912 60902
rect 32616 59866 32672 59868
rect 32696 59866 32752 59868
rect 32776 59866 32832 59868
rect 32856 59866 32912 59868
rect 32616 59814 32662 59866
rect 32662 59814 32672 59866
rect 32696 59814 32726 59866
rect 32726 59814 32738 59866
rect 32738 59814 32752 59866
rect 32776 59814 32790 59866
rect 32790 59814 32802 59866
rect 32802 59814 32832 59866
rect 32856 59814 32866 59866
rect 32866 59814 32912 59866
rect 32616 59812 32672 59814
rect 32696 59812 32752 59814
rect 32776 59812 32832 59814
rect 32856 59812 32912 59814
rect 32616 58778 32672 58780
rect 32696 58778 32752 58780
rect 32776 58778 32832 58780
rect 32856 58778 32912 58780
rect 32616 58726 32662 58778
rect 32662 58726 32672 58778
rect 32696 58726 32726 58778
rect 32726 58726 32738 58778
rect 32738 58726 32752 58778
rect 32776 58726 32790 58778
rect 32790 58726 32802 58778
rect 32802 58726 32832 58778
rect 32856 58726 32866 58778
rect 32866 58726 32912 58778
rect 32616 58724 32672 58726
rect 32696 58724 32752 58726
rect 32776 58724 32832 58726
rect 32856 58724 32912 58726
rect 32616 57690 32672 57692
rect 32696 57690 32752 57692
rect 32776 57690 32832 57692
rect 32856 57690 32912 57692
rect 32616 57638 32662 57690
rect 32662 57638 32672 57690
rect 32696 57638 32726 57690
rect 32726 57638 32738 57690
rect 32738 57638 32752 57690
rect 32776 57638 32790 57690
rect 32790 57638 32802 57690
rect 32802 57638 32832 57690
rect 32856 57638 32866 57690
rect 32866 57638 32912 57690
rect 32616 57636 32672 57638
rect 32696 57636 32752 57638
rect 32776 57636 32832 57638
rect 32856 57636 32912 57638
rect 32616 56602 32672 56604
rect 32696 56602 32752 56604
rect 32776 56602 32832 56604
rect 32856 56602 32912 56604
rect 32616 56550 32662 56602
rect 32662 56550 32672 56602
rect 32696 56550 32726 56602
rect 32726 56550 32738 56602
rect 32738 56550 32752 56602
rect 32776 56550 32790 56602
rect 32790 56550 32802 56602
rect 32802 56550 32832 56602
rect 32856 56550 32866 56602
rect 32866 56550 32912 56602
rect 32616 56548 32672 56550
rect 32696 56548 32752 56550
rect 32776 56548 32832 56550
rect 32856 56548 32912 56550
rect 32616 55514 32672 55516
rect 32696 55514 32752 55516
rect 32776 55514 32832 55516
rect 32856 55514 32912 55516
rect 32616 55462 32662 55514
rect 32662 55462 32672 55514
rect 32696 55462 32726 55514
rect 32726 55462 32738 55514
rect 32738 55462 32752 55514
rect 32776 55462 32790 55514
rect 32790 55462 32802 55514
rect 32802 55462 32832 55514
rect 32856 55462 32866 55514
rect 32866 55462 32912 55514
rect 32616 55460 32672 55462
rect 32696 55460 32752 55462
rect 32776 55460 32832 55462
rect 32856 55460 32912 55462
rect 32616 54426 32672 54428
rect 32696 54426 32752 54428
rect 32776 54426 32832 54428
rect 32856 54426 32912 54428
rect 32616 54374 32662 54426
rect 32662 54374 32672 54426
rect 32696 54374 32726 54426
rect 32726 54374 32738 54426
rect 32738 54374 32752 54426
rect 32776 54374 32790 54426
rect 32790 54374 32802 54426
rect 32802 54374 32832 54426
rect 32856 54374 32866 54426
rect 32866 54374 32912 54426
rect 32616 54372 32672 54374
rect 32696 54372 32752 54374
rect 32776 54372 32832 54374
rect 32856 54372 32912 54374
rect 32616 53338 32672 53340
rect 32696 53338 32752 53340
rect 32776 53338 32832 53340
rect 32856 53338 32912 53340
rect 32616 53286 32662 53338
rect 32662 53286 32672 53338
rect 32696 53286 32726 53338
rect 32726 53286 32738 53338
rect 32738 53286 32752 53338
rect 32776 53286 32790 53338
rect 32790 53286 32802 53338
rect 32802 53286 32832 53338
rect 32856 53286 32866 53338
rect 32866 53286 32912 53338
rect 32616 53284 32672 53286
rect 32696 53284 32752 53286
rect 32776 53284 32832 53286
rect 32856 53284 32912 53286
rect 32616 52250 32672 52252
rect 32696 52250 32752 52252
rect 32776 52250 32832 52252
rect 32856 52250 32912 52252
rect 32616 52198 32662 52250
rect 32662 52198 32672 52250
rect 32696 52198 32726 52250
rect 32726 52198 32738 52250
rect 32738 52198 32752 52250
rect 32776 52198 32790 52250
rect 32790 52198 32802 52250
rect 32802 52198 32832 52250
rect 32856 52198 32866 52250
rect 32866 52198 32912 52250
rect 32616 52196 32672 52198
rect 32696 52196 32752 52198
rect 32776 52196 32832 52198
rect 32856 52196 32912 52198
rect 32616 51162 32672 51164
rect 32696 51162 32752 51164
rect 32776 51162 32832 51164
rect 32856 51162 32912 51164
rect 32616 51110 32662 51162
rect 32662 51110 32672 51162
rect 32696 51110 32726 51162
rect 32726 51110 32738 51162
rect 32738 51110 32752 51162
rect 32776 51110 32790 51162
rect 32790 51110 32802 51162
rect 32802 51110 32832 51162
rect 32856 51110 32866 51162
rect 32866 51110 32912 51162
rect 32616 51108 32672 51110
rect 32696 51108 32752 51110
rect 32776 51108 32832 51110
rect 32856 51108 32912 51110
rect 31956 50618 32012 50620
rect 32036 50618 32092 50620
rect 32116 50618 32172 50620
rect 32196 50618 32252 50620
rect 31956 50566 32002 50618
rect 32002 50566 32012 50618
rect 32036 50566 32066 50618
rect 32066 50566 32078 50618
rect 32078 50566 32092 50618
rect 32116 50566 32130 50618
rect 32130 50566 32142 50618
rect 32142 50566 32172 50618
rect 32196 50566 32206 50618
rect 32206 50566 32252 50618
rect 31956 50564 32012 50566
rect 32036 50564 32092 50566
rect 32116 50564 32172 50566
rect 32196 50564 32252 50566
rect 32616 50074 32672 50076
rect 32696 50074 32752 50076
rect 32776 50074 32832 50076
rect 32856 50074 32912 50076
rect 32616 50022 32662 50074
rect 32662 50022 32672 50074
rect 32696 50022 32726 50074
rect 32726 50022 32738 50074
rect 32738 50022 32752 50074
rect 32776 50022 32790 50074
rect 32790 50022 32802 50074
rect 32802 50022 32832 50074
rect 32856 50022 32866 50074
rect 32866 50022 32912 50074
rect 32616 50020 32672 50022
rect 32696 50020 32752 50022
rect 32776 50020 32832 50022
rect 32856 50020 32912 50022
rect 31956 49530 32012 49532
rect 32036 49530 32092 49532
rect 32116 49530 32172 49532
rect 32196 49530 32252 49532
rect 31956 49478 32002 49530
rect 32002 49478 32012 49530
rect 32036 49478 32066 49530
rect 32066 49478 32078 49530
rect 32078 49478 32092 49530
rect 32116 49478 32130 49530
rect 32130 49478 32142 49530
rect 32142 49478 32172 49530
rect 32196 49478 32206 49530
rect 32206 49478 32252 49530
rect 31956 49476 32012 49478
rect 32036 49476 32092 49478
rect 32116 49476 32172 49478
rect 32196 49476 32252 49478
rect 32616 48986 32672 48988
rect 32696 48986 32752 48988
rect 32776 48986 32832 48988
rect 32856 48986 32912 48988
rect 32616 48934 32662 48986
rect 32662 48934 32672 48986
rect 32696 48934 32726 48986
rect 32726 48934 32738 48986
rect 32738 48934 32752 48986
rect 32776 48934 32790 48986
rect 32790 48934 32802 48986
rect 32802 48934 32832 48986
rect 32856 48934 32866 48986
rect 32866 48934 32912 48986
rect 32616 48932 32672 48934
rect 32696 48932 32752 48934
rect 32776 48932 32832 48934
rect 32856 48932 32912 48934
rect 31956 48442 32012 48444
rect 32036 48442 32092 48444
rect 32116 48442 32172 48444
rect 32196 48442 32252 48444
rect 31956 48390 32002 48442
rect 32002 48390 32012 48442
rect 32036 48390 32066 48442
rect 32066 48390 32078 48442
rect 32078 48390 32092 48442
rect 32116 48390 32130 48442
rect 32130 48390 32142 48442
rect 32142 48390 32172 48442
rect 32196 48390 32206 48442
rect 32206 48390 32252 48442
rect 31956 48388 32012 48390
rect 32036 48388 32092 48390
rect 32116 48388 32172 48390
rect 32196 48388 32252 48390
rect 32616 47898 32672 47900
rect 32696 47898 32752 47900
rect 32776 47898 32832 47900
rect 32856 47898 32912 47900
rect 32616 47846 32662 47898
rect 32662 47846 32672 47898
rect 32696 47846 32726 47898
rect 32726 47846 32738 47898
rect 32738 47846 32752 47898
rect 32776 47846 32790 47898
rect 32790 47846 32802 47898
rect 32802 47846 32832 47898
rect 32856 47846 32866 47898
rect 32866 47846 32912 47898
rect 32616 47844 32672 47846
rect 32696 47844 32752 47846
rect 32776 47844 32832 47846
rect 32856 47844 32912 47846
rect 31956 47354 32012 47356
rect 32036 47354 32092 47356
rect 32116 47354 32172 47356
rect 32196 47354 32252 47356
rect 31956 47302 32002 47354
rect 32002 47302 32012 47354
rect 32036 47302 32066 47354
rect 32066 47302 32078 47354
rect 32078 47302 32092 47354
rect 32116 47302 32130 47354
rect 32130 47302 32142 47354
rect 32142 47302 32172 47354
rect 32196 47302 32206 47354
rect 32206 47302 32252 47354
rect 31956 47300 32012 47302
rect 32036 47300 32092 47302
rect 32116 47300 32172 47302
rect 32196 47300 32252 47302
rect 32616 46810 32672 46812
rect 32696 46810 32752 46812
rect 32776 46810 32832 46812
rect 32856 46810 32912 46812
rect 32616 46758 32662 46810
rect 32662 46758 32672 46810
rect 32696 46758 32726 46810
rect 32726 46758 32738 46810
rect 32738 46758 32752 46810
rect 32776 46758 32790 46810
rect 32790 46758 32802 46810
rect 32802 46758 32832 46810
rect 32856 46758 32866 46810
rect 32866 46758 32912 46810
rect 32616 46756 32672 46758
rect 32696 46756 32752 46758
rect 32776 46756 32832 46758
rect 32856 46756 32912 46758
rect 31956 46266 32012 46268
rect 32036 46266 32092 46268
rect 32116 46266 32172 46268
rect 32196 46266 32252 46268
rect 31956 46214 32002 46266
rect 32002 46214 32012 46266
rect 32036 46214 32066 46266
rect 32066 46214 32078 46266
rect 32078 46214 32092 46266
rect 32116 46214 32130 46266
rect 32130 46214 32142 46266
rect 32142 46214 32172 46266
rect 32196 46214 32206 46266
rect 32206 46214 32252 46266
rect 31956 46212 32012 46214
rect 32036 46212 32092 46214
rect 32116 46212 32172 46214
rect 32196 46212 32252 46214
rect 32616 45722 32672 45724
rect 32696 45722 32752 45724
rect 32776 45722 32832 45724
rect 32856 45722 32912 45724
rect 32616 45670 32662 45722
rect 32662 45670 32672 45722
rect 32696 45670 32726 45722
rect 32726 45670 32738 45722
rect 32738 45670 32752 45722
rect 32776 45670 32790 45722
rect 32790 45670 32802 45722
rect 32802 45670 32832 45722
rect 32856 45670 32866 45722
rect 32866 45670 32912 45722
rect 32616 45668 32672 45670
rect 32696 45668 32752 45670
rect 32776 45668 32832 45670
rect 32856 45668 32912 45670
rect 31956 45178 32012 45180
rect 32036 45178 32092 45180
rect 32116 45178 32172 45180
rect 32196 45178 32252 45180
rect 31956 45126 32002 45178
rect 32002 45126 32012 45178
rect 32036 45126 32066 45178
rect 32066 45126 32078 45178
rect 32078 45126 32092 45178
rect 32116 45126 32130 45178
rect 32130 45126 32142 45178
rect 32142 45126 32172 45178
rect 32196 45126 32206 45178
rect 32206 45126 32252 45178
rect 31956 45124 32012 45126
rect 32036 45124 32092 45126
rect 32116 45124 32172 45126
rect 32196 45124 32252 45126
rect 31956 44090 32012 44092
rect 32036 44090 32092 44092
rect 32116 44090 32172 44092
rect 32196 44090 32252 44092
rect 31956 44038 32002 44090
rect 32002 44038 32012 44090
rect 32036 44038 32066 44090
rect 32066 44038 32078 44090
rect 32078 44038 32092 44090
rect 32116 44038 32130 44090
rect 32130 44038 32142 44090
rect 32142 44038 32172 44090
rect 32196 44038 32206 44090
rect 32206 44038 32252 44090
rect 31956 44036 32012 44038
rect 32036 44036 32092 44038
rect 32116 44036 32172 44038
rect 32196 44036 32252 44038
rect 31956 43002 32012 43004
rect 32036 43002 32092 43004
rect 32116 43002 32172 43004
rect 32196 43002 32252 43004
rect 31956 42950 32002 43002
rect 32002 42950 32012 43002
rect 32036 42950 32066 43002
rect 32066 42950 32078 43002
rect 32078 42950 32092 43002
rect 32116 42950 32130 43002
rect 32130 42950 32142 43002
rect 32142 42950 32172 43002
rect 32196 42950 32206 43002
rect 32206 42950 32252 43002
rect 31956 42948 32012 42950
rect 32036 42948 32092 42950
rect 32116 42948 32172 42950
rect 32196 42948 32252 42950
rect 31956 41914 32012 41916
rect 32036 41914 32092 41916
rect 32116 41914 32172 41916
rect 32196 41914 32252 41916
rect 31956 41862 32002 41914
rect 32002 41862 32012 41914
rect 32036 41862 32066 41914
rect 32066 41862 32078 41914
rect 32078 41862 32092 41914
rect 32116 41862 32130 41914
rect 32130 41862 32142 41914
rect 32142 41862 32172 41914
rect 32196 41862 32206 41914
rect 32206 41862 32252 41914
rect 31956 41860 32012 41862
rect 32036 41860 32092 41862
rect 32116 41860 32172 41862
rect 32196 41860 32252 41862
rect 31956 40826 32012 40828
rect 32036 40826 32092 40828
rect 32116 40826 32172 40828
rect 32196 40826 32252 40828
rect 31956 40774 32002 40826
rect 32002 40774 32012 40826
rect 32036 40774 32066 40826
rect 32066 40774 32078 40826
rect 32078 40774 32092 40826
rect 32116 40774 32130 40826
rect 32130 40774 32142 40826
rect 32142 40774 32172 40826
rect 32196 40774 32206 40826
rect 32206 40774 32252 40826
rect 31956 40772 32012 40774
rect 32036 40772 32092 40774
rect 32116 40772 32172 40774
rect 32196 40772 32252 40774
rect 32616 44634 32672 44636
rect 32696 44634 32752 44636
rect 32776 44634 32832 44636
rect 32856 44634 32912 44636
rect 32616 44582 32662 44634
rect 32662 44582 32672 44634
rect 32696 44582 32726 44634
rect 32726 44582 32738 44634
rect 32738 44582 32752 44634
rect 32776 44582 32790 44634
rect 32790 44582 32802 44634
rect 32802 44582 32832 44634
rect 32856 44582 32866 44634
rect 32866 44582 32912 44634
rect 32616 44580 32672 44582
rect 32696 44580 32752 44582
rect 32776 44580 32832 44582
rect 32856 44580 32912 44582
rect 31956 39738 32012 39740
rect 32036 39738 32092 39740
rect 32116 39738 32172 39740
rect 32196 39738 32252 39740
rect 31956 39686 32002 39738
rect 32002 39686 32012 39738
rect 32036 39686 32066 39738
rect 32066 39686 32078 39738
rect 32078 39686 32092 39738
rect 32116 39686 32130 39738
rect 32130 39686 32142 39738
rect 32142 39686 32172 39738
rect 32196 39686 32206 39738
rect 32206 39686 32252 39738
rect 31956 39684 32012 39686
rect 32036 39684 32092 39686
rect 32116 39684 32172 39686
rect 32196 39684 32252 39686
rect 31956 38650 32012 38652
rect 32036 38650 32092 38652
rect 32116 38650 32172 38652
rect 32196 38650 32252 38652
rect 31956 38598 32002 38650
rect 32002 38598 32012 38650
rect 32036 38598 32066 38650
rect 32066 38598 32078 38650
rect 32078 38598 32092 38650
rect 32116 38598 32130 38650
rect 32130 38598 32142 38650
rect 32142 38598 32172 38650
rect 32196 38598 32206 38650
rect 32206 38598 32252 38650
rect 31956 38596 32012 38598
rect 32036 38596 32092 38598
rect 32116 38596 32172 38598
rect 32196 38596 32252 38598
rect 31956 37562 32012 37564
rect 32036 37562 32092 37564
rect 32116 37562 32172 37564
rect 32196 37562 32252 37564
rect 31956 37510 32002 37562
rect 32002 37510 32012 37562
rect 32036 37510 32066 37562
rect 32066 37510 32078 37562
rect 32078 37510 32092 37562
rect 32116 37510 32130 37562
rect 32130 37510 32142 37562
rect 32142 37510 32172 37562
rect 32196 37510 32206 37562
rect 32206 37510 32252 37562
rect 31956 37508 32012 37510
rect 32036 37508 32092 37510
rect 32116 37508 32172 37510
rect 32196 37508 32252 37510
rect 31956 36474 32012 36476
rect 32036 36474 32092 36476
rect 32116 36474 32172 36476
rect 32196 36474 32252 36476
rect 31956 36422 32002 36474
rect 32002 36422 32012 36474
rect 32036 36422 32066 36474
rect 32066 36422 32078 36474
rect 32078 36422 32092 36474
rect 32116 36422 32130 36474
rect 32130 36422 32142 36474
rect 32142 36422 32172 36474
rect 32196 36422 32206 36474
rect 32206 36422 32252 36474
rect 31956 36420 32012 36422
rect 32036 36420 32092 36422
rect 32116 36420 32172 36422
rect 32196 36420 32252 36422
rect 31956 35386 32012 35388
rect 32036 35386 32092 35388
rect 32116 35386 32172 35388
rect 32196 35386 32252 35388
rect 31956 35334 32002 35386
rect 32002 35334 32012 35386
rect 32036 35334 32066 35386
rect 32066 35334 32078 35386
rect 32078 35334 32092 35386
rect 32116 35334 32130 35386
rect 32130 35334 32142 35386
rect 32142 35334 32172 35386
rect 32196 35334 32206 35386
rect 32206 35334 32252 35386
rect 31956 35332 32012 35334
rect 32036 35332 32092 35334
rect 32116 35332 32172 35334
rect 32196 35332 32252 35334
rect 31956 34298 32012 34300
rect 32036 34298 32092 34300
rect 32116 34298 32172 34300
rect 32196 34298 32252 34300
rect 31956 34246 32002 34298
rect 32002 34246 32012 34298
rect 32036 34246 32066 34298
rect 32066 34246 32078 34298
rect 32078 34246 32092 34298
rect 32116 34246 32130 34298
rect 32130 34246 32142 34298
rect 32142 34246 32172 34298
rect 32196 34246 32206 34298
rect 32206 34246 32252 34298
rect 31956 34244 32012 34246
rect 32036 34244 32092 34246
rect 32116 34244 32172 34246
rect 32196 34244 32252 34246
rect 31956 33210 32012 33212
rect 32036 33210 32092 33212
rect 32116 33210 32172 33212
rect 32196 33210 32252 33212
rect 31956 33158 32002 33210
rect 32002 33158 32012 33210
rect 32036 33158 32066 33210
rect 32066 33158 32078 33210
rect 32078 33158 32092 33210
rect 32116 33158 32130 33210
rect 32130 33158 32142 33210
rect 32142 33158 32172 33210
rect 32196 33158 32206 33210
rect 32206 33158 32252 33210
rect 31956 33156 32012 33158
rect 32036 33156 32092 33158
rect 32116 33156 32172 33158
rect 32196 33156 32252 33158
rect 31956 32122 32012 32124
rect 32036 32122 32092 32124
rect 32116 32122 32172 32124
rect 32196 32122 32252 32124
rect 31956 32070 32002 32122
rect 32002 32070 32012 32122
rect 32036 32070 32066 32122
rect 32066 32070 32078 32122
rect 32078 32070 32092 32122
rect 32116 32070 32130 32122
rect 32130 32070 32142 32122
rect 32142 32070 32172 32122
rect 32196 32070 32206 32122
rect 32206 32070 32252 32122
rect 31956 32068 32012 32070
rect 32036 32068 32092 32070
rect 32116 32068 32172 32070
rect 32196 32068 32252 32070
rect 31956 31034 32012 31036
rect 32036 31034 32092 31036
rect 32116 31034 32172 31036
rect 32196 31034 32252 31036
rect 31956 30982 32002 31034
rect 32002 30982 32012 31034
rect 32036 30982 32066 31034
rect 32066 30982 32078 31034
rect 32078 30982 32092 31034
rect 32116 30982 32130 31034
rect 32130 30982 32142 31034
rect 32142 30982 32172 31034
rect 32196 30982 32206 31034
rect 32206 30982 32252 31034
rect 31956 30980 32012 30982
rect 32036 30980 32092 30982
rect 32116 30980 32172 30982
rect 32196 30980 32252 30982
rect 31956 29946 32012 29948
rect 32036 29946 32092 29948
rect 32116 29946 32172 29948
rect 32196 29946 32252 29948
rect 31956 29894 32002 29946
rect 32002 29894 32012 29946
rect 32036 29894 32066 29946
rect 32066 29894 32078 29946
rect 32078 29894 32092 29946
rect 32116 29894 32130 29946
rect 32130 29894 32142 29946
rect 32142 29894 32172 29946
rect 32196 29894 32206 29946
rect 32206 29894 32252 29946
rect 31956 29892 32012 29894
rect 32036 29892 32092 29894
rect 32116 29892 32172 29894
rect 32196 29892 32252 29894
rect 31956 28858 32012 28860
rect 32036 28858 32092 28860
rect 32116 28858 32172 28860
rect 32196 28858 32252 28860
rect 31956 28806 32002 28858
rect 32002 28806 32012 28858
rect 32036 28806 32066 28858
rect 32066 28806 32078 28858
rect 32078 28806 32092 28858
rect 32116 28806 32130 28858
rect 32130 28806 32142 28858
rect 32142 28806 32172 28858
rect 32196 28806 32206 28858
rect 32206 28806 32252 28858
rect 31956 28804 32012 28806
rect 32036 28804 32092 28806
rect 32116 28804 32172 28806
rect 32196 28804 32252 28806
rect 31956 27770 32012 27772
rect 32036 27770 32092 27772
rect 32116 27770 32172 27772
rect 32196 27770 32252 27772
rect 31956 27718 32002 27770
rect 32002 27718 32012 27770
rect 32036 27718 32066 27770
rect 32066 27718 32078 27770
rect 32078 27718 32092 27770
rect 32116 27718 32130 27770
rect 32130 27718 32142 27770
rect 32142 27718 32172 27770
rect 32196 27718 32206 27770
rect 32206 27718 32252 27770
rect 31956 27716 32012 27718
rect 32036 27716 32092 27718
rect 32116 27716 32172 27718
rect 32196 27716 32252 27718
rect 31956 26682 32012 26684
rect 32036 26682 32092 26684
rect 32116 26682 32172 26684
rect 32196 26682 32252 26684
rect 31956 26630 32002 26682
rect 32002 26630 32012 26682
rect 32036 26630 32066 26682
rect 32066 26630 32078 26682
rect 32078 26630 32092 26682
rect 32116 26630 32130 26682
rect 32130 26630 32142 26682
rect 32142 26630 32172 26682
rect 32196 26630 32206 26682
rect 32206 26630 32252 26682
rect 31956 26628 32012 26630
rect 32036 26628 32092 26630
rect 32116 26628 32172 26630
rect 32196 26628 32252 26630
rect 31956 25594 32012 25596
rect 32036 25594 32092 25596
rect 32116 25594 32172 25596
rect 32196 25594 32252 25596
rect 31956 25542 32002 25594
rect 32002 25542 32012 25594
rect 32036 25542 32066 25594
rect 32066 25542 32078 25594
rect 32078 25542 32092 25594
rect 32116 25542 32130 25594
rect 32130 25542 32142 25594
rect 32142 25542 32172 25594
rect 32196 25542 32206 25594
rect 32206 25542 32252 25594
rect 31956 25540 32012 25542
rect 32036 25540 32092 25542
rect 32116 25540 32172 25542
rect 32196 25540 32252 25542
rect 31956 24506 32012 24508
rect 32036 24506 32092 24508
rect 32116 24506 32172 24508
rect 32196 24506 32252 24508
rect 31956 24454 32002 24506
rect 32002 24454 32012 24506
rect 32036 24454 32066 24506
rect 32066 24454 32078 24506
rect 32078 24454 32092 24506
rect 32116 24454 32130 24506
rect 32130 24454 32142 24506
rect 32142 24454 32172 24506
rect 32196 24454 32206 24506
rect 32206 24454 32252 24506
rect 31956 24452 32012 24454
rect 32036 24452 32092 24454
rect 32116 24452 32172 24454
rect 32196 24452 32252 24454
rect 31956 23418 32012 23420
rect 32036 23418 32092 23420
rect 32116 23418 32172 23420
rect 32196 23418 32252 23420
rect 31956 23366 32002 23418
rect 32002 23366 32012 23418
rect 32036 23366 32066 23418
rect 32066 23366 32078 23418
rect 32078 23366 32092 23418
rect 32116 23366 32130 23418
rect 32130 23366 32142 23418
rect 32142 23366 32172 23418
rect 32196 23366 32206 23418
rect 32206 23366 32252 23418
rect 31956 23364 32012 23366
rect 32036 23364 32092 23366
rect 32116 23364 32172 23366
rect 32196 23364 32252 23366
rect 31956 22330 32012 22332
rect 32036 22330 32092 22332
rect 32116 22330 32172 22332
rect 32196 22330 32252 22332
rect 31956 22278 32002 22330
rect 32002 22278 32012 22330
rect 32036 22278 32066 22330
rect 32066 22278 32078 22330
rect 32078 22278 32092 22330
rect 32116 22278 32130 22330
rect 32130 22278 32142 22330
rect 32142 22278 32172 22330
rect 32196 22278 32206 22330
rect 32206 22278 32252 22330
rect 31956 22276 32012 22278
rect 32036 22276 32092 22278
rect 32116 22276 32172 22278
rect 32196 22276 32252 22278
rect 31956 21242 32012 21244
rect 32036 21242 32092 21244
rect 32116 21242 32172 21244
rect 32196 21242 32252 21244
rect 31956 21190 32002 21242
rect 32002 21190 32012 21242
rect 32036 21190 32066 21242
rect 32066 21190 32078 21242
rect 32078 21190 32092 21242
rect 32116 21190 32130 21242
rect 32130 21190 32142 21242
rect 32142 21190 32172 21242
rect 32196 21190 32206 21242
rect 32206 21190 32252 21242
rect 31956 21188 32012 21190
rect 32036 21188 32092 21190
rect 32116 21188 32172 21190
rect 32196 21188 32252 21190
rect 31956 20154 32012 20156
rect 32036 20154 32092 20156
rect 32116 20154 32172 20156
rect 32196 20154 32252 20156
rect 31956 20102 32002 20154
rect 32002 20102 32012 20154
rect 32036 20102 32066 20154
rect 32066 20102 32078 20154
rect 32078 20102 32092 20154
rect 32116 20102 32130 20154
rect 32130 20102 32142 20154
rect 32142 20102 32172 20154
rect 32196 20102 32206 20154
rect 32206 20102 32252 20154
rect 31956 20100 32012 20102
rect 32036 20100 32092 20102
rect 32116 20100 32172 20102
rect 32196 20100 32252 20102
rect 31956 19066 32012 19068
rect 32036 19066 32092 19068
rect 32116 19066 32172 19068
rect 32196 19066 32252 19068
rect 31956 19014 32002 19066
rect 32002 19014 32012 19066
rect 32036 19014 32066 19066
rect 32066 19014 32078 19066
rect 32078 19014 32092 19066
rect 32116 19014 32130 19066
rect 32130 19014 32142 19066
rect 32142 19014 32172 19066
rect 32196 19014 32206 19066
rect 32206 19014 32252 19066
rect 31956 19012 32012 19014
rect 32036 19012 32092 19014
rect 32116 19012 32172 19014
rect 32196 19012 32252 19014
rect 31956 17978 32012 17980
rect 32036 17978 32092 17980
rect 32116 17978 32172 17980
rect 32196 17978 32252 17980
rect 31956 17926 32002 17978
rect 32002 17926 32012 17978
rect 32036 17926 32066 17978
rect 32066 17926 32078 17978
rect 32078 17926 32092 17978
rect 32116 17926 32130 17978
rect 32130 17926 32142 17978
rect 32142 17926 32172 17978
rect 32196 17926 32206 17978
rect 32206 17926 32252 17978
rect 31956 17924 32012 17926
rect 32036 17924 32092 17926
rect 32116 17924 32172 17926
rect 32196 17924 32252 17926
rect 31956 16890 32012 16892
rect 32036 16890 32092 16892
rect 32116 16890 32172 16892
rect 32196 16890 32252 16892
rect 31956 16838 32002 16890
rect 32002 16838 32012 16890
rect 32036 16838 32066 16890
rect 32066 16838 32078 16890
rect 32078 16838 32092 16890
rect 32116 16838 32130 16890
rect 32130 16838 32142 16890
rect 32142 16838 32172 16890
rect 32196 16838 32206 16890
rect 32206 16838 32252 16890
rect 31956 16836 32012 16838
rect 32036 16836 32092 16838
rect 32116 16836 32172 16838
rect 32196 16836 32252 16838
rect 31956 15802 32012 15804
rect 32036 15802 32092 15804
rect 32116 15802 32172 15804
rect 32196 15802 32252 15804
rect 31956 15750 32002 15802
rect 32002 15750 32012 15802
rect 32036 15750 32066 15802
rect 32066 15750 32078 15802
rect 32078 15750 32092 15802
rect 32116 15750 32130 15802
rect 32130 15750 32142 15802
rect 32142 15750 32172 15802
rect 32196 15750 32206 15802
rect 32206 15750 32252 15802
rect 31956 15748 32012 15750
rect 32036 15748 32092 15750
rect 32116 15748 32172 15750
rect 32196 15748 32252 15750
rect 31956 14714 32012 14716
rect 32036 14714 32092 14716
rect 32116 14714 32172 14716
rect 32196 14714 32252 14716
rect 31956 14662 32002 14714
rect 32002 14662 32012 14714
rect 32036 14662 32066 14714
rect 32066 14662 32078 14714
rect 32078 14662 32092 14714
rect 32116 14662 32130 14714
rect 32130 14662 32142 14714
rect 32142 14662 32172 14714
rect 32196 14662 32206 14714
rect 32206 14662 32252 14714
rect 31956 14660 32012 14662
rect 32036 14660 32092 14662
rect 32116 14660 32172 14662
rect 32196 14660 32252 14662
rect 32616 43546 32672 43548
rect 32696 43546 32752 43548
rect 32776 43546 32832 43548
rect 32856 43546 32912 43548
rect 32616 43494 32662 43546
rect 32662 43494 32672 43546
rect 32696 43494 32726 43546
rect 32726 43494 32738 43546
rect 32738 43494 32752 43546
rect 32776 43494 32790 43546
rect 32790 43494 32802 43546
rect 32802 43494 32832 43546
rect 32856 43494 32866 43546
rect 32866 43494 32912 43546
rect 32616 43492 32672 43494
rect 32696 43492 32752 43494
rect 32776 43492 32832 43494
rect 32856 43492 32912 43494
rect 32616 42458 32672 42460
rect 32696 42458 32752 42460
rect 32776 42458 32832 42460
rect 32856 42458 32912 42460
rect 32616 42406 32662 42458
rect 32662 42406 32672 42458
rect 32696 42406 32726 42458
rect 32726 42406 32738 42458
rect 32738 42406 32752 42458
rect 32776 42406 32790 42458
rect 32790 42406 32802 42458
rect 32802 42406 32832 42458
rect 32856 42406 32866 42458
rect 32866 42406 32912 42458
rect 32616 42404 32672 42406
rect 32696 42404 32752 42406
rect 32776 42404 32832 42406
rect 32856 42404 32912 42406
rect 32616 41370 32672 41372
rect 32696 41370 32752 41372
rect 32776 41370 32832 41372
rect 32856 41370 32912 41372
rect 32616 41318 32662 41370
rect 32662 41318 32672 41370
rect 32696 41318 32726 41370
rect 32726 41318 32738 41370
rect 32738 41318 32752 41370
rect 32776 41318 32790 41370
rect 32790 41318 32802 41370
rect 32802 41318 32832 41370
rect 32856 41318 32866 41370
rect 32866 41318 32912 41370
rect 32616 41316 32672 41318
rect 32696 41316 32752 41318
rect 32776 41316 32832 41318
rect 32856 41316 32912 41318
rect 32616 40282 32672 40284
rect 32696 40282 32752 40284
rect 32776 40282 32832 40284
rect 32856 40282 32912 40284
rect 32616 40230 32662 40282
rect 32662 40230 32672 40282
rect 32696 40230 32726 40282
rect 32726 40230 32738 40282
rect 32738 40230 32752 40282
rect 32776 40230 32790 40282
rect 32790 40230 32802 40282
rect 32802 40230 32832 40282
rect 32856 40230 32866 40282
rect 32866 40230 32912 40282
rect 32616 40228 32672 40230
rect 32696 40228 32752 40230
rect 32776 40228 32832 40230
rect 32856 40228 32912 40230
rect 32616 39194 32672 39196
rect 32696 39194 32752 39196
rect 32776 39194 32832 39196
rect 32856 39194 32912 39196
rect 32616 39142 32662 39194
rect 32662 39142 32672 39194
rect 32696 39142 32726 39194
rect 32726 39142 32738 39194
rect 32738 39142 32752 39194
rect 32776 39142 32790 39194
rect 32790 39142 32802 39194
rect 32802 39142 32832 39194
rect 32856 39142 32866 39194
rect 32866 39142 32912 39194
rect 32616 39140 32672 39142
rect 32696 39140 32752 39142
rect 32776 39140 32832 39142
rect 32856 39140 32912 39142
rect 32616 38106 32672 38108
rect 32696 38106 32752 38108
rect 32776 38106 32832 38108
rect 32856 38106 32912 38108
rect 32616 38054 32662 38106
rect 32662 38054 32672 38106
rect 32696 38054 32726 38106
rect 32726 38054 32738 38106
rect 32738 38054 32752 38106
rect 32776 38054 32790 38106
rect 32790 38054 32802 38106
rect 32802 38054 32832 38106
rect 32856 38054 32866 38106
rect 32866 38054 32912 38106
rect 32616 38052 32672 38054
rect 32696 38052 32752 38054
rect 32776 38052 32832 38054
rect 32856 38052 32912 38054
rect 32616 37018 32672 37020
rect 32696 37018 32752 37020
rect 32776 37018 32832 37020
rect 32856 37018 32912 37020
rect 32616 36966 32662 37018
rect 32662 36966 32672 37018
rect 32696 36966 32726 37018
rect 32726 36966 32738 37018
rect 32738 36966 32752 37018
rect 32776 36966 32790 37018
rect 32790 36966 32802 37018
rect 32802 36966 32832 37018
rect 32856 36966 32866 37018
rect 32866 36966 32912 37018
rect 32616 36964 32672 36966
rect 32696 36964 32752 36966
rect 32776 36964 32832 36966
rect 32856 36964 32912 36966
rect 32616 35930 32672 35932
rect 32696 35930 32752 35932
rect 32776 35930 32832 35932
rect 32856 35930 32912 35932
rect 32616 35878 32662 35930
rect 32662 35878 32672 35930
rect 32696 35878 32726 35930
rect 32726 35878 32738 35930
rect 32738 35878 32752 35930
rect 32776 35878 32790 35930
rect 32790 35878 32802 35930
rect 32802 35878 32832 35930
rect 32856 35878 32866 35930
rect 32866 35878 32912 35930
rect 32616 35876 32672 35878
rect 32696 35876 32752 35878
rect 32776 35876 32832 35878
rect 32856 35876 32912 35878
rect 32616 34842 32672 34844
rect 32696 34842 32752 34844
rect 32776 34842 32832 34844
rect 32856 34842 32912 34844
rect 32616 34790 32662 34842
rect 32662 34790 32672 34842
rect 32696 34790 32726 34842
rect 32726 34790 32738 34842
rect 32738 34790 32752 34842
rect 32776 34790 32790 34842
rect 32790 34790 32802 34842
rect 32802 34790 32832 34842
rect 32856 34790 32866 34842
rect 32866 34790 32912 34842
rect 32616 34788 32672 34790
rect 32696 34788 32752 34790
rect 32776 34788 32832 34790
rect 32856 34788 32912 34790
rect 32616 33754 32672 33756
rect 32696 33754 32752 33756
rect 32776 33754 32832 33756
rect 32856 33754 32912 33756
rect 32616 33702 32662 33754
rect 32662 33702 32672 33754
rect 32696 33702 32726 33754
rect 32726 33702 32738 33754
rect 32738 33702 32752 33754
rect 32776 33702 32790 33754
rect 32790 33702 32802 33754
rect 32802 33702 32832 33754
rect 32856 33702 32866 33754
rect 32866 33702 32912 33754
rect 32616 33700 32672 33702
rect 32696 33700 32752 33702
rect 32776 33700 32832 33702
rect 32856 33700 32912 33702
rect 32616 32666 32672 32668
rect 32696 32666 32752 32668
rect 32776 32666 32832 32668
rect 32856 32666 32912 32668
rect 32616 32614 32662 32666
rect 32662 32614 32672 32666
rect 32696 32614 32726 32666
rect 32726 32614 32738 32666
rect 32738 32614 32752 32666
rect 32776 32614 32790 32666
rect 32790 32614 32802 32666
rect 32802 32614 32832 32666
rect 32856 32614 32866 32666
rect 32866 32614 32912 32666
rect 32616 32612 32672 32614
rect 32696 32612 32752 32614
rect 32776 32612 32832 32614
rect 32856 32612 32912 32614
rect 32616 31578 32672 31580
rect 32696 31578 32752 31580
rect 32776 31578 32832 31580
rect 32856 31578 32912 31580
rect 32616 31526 32662 31578
rect 32662 31526 32672 31578
rect 32696 31526 32726 31578
rect 32726 31526 32738 31578
rect 32738 31526 32752 31578
rect 32776 31526 32790 31578
rect 32790 31526 32802 31578
rect 32802 31526 32832 31578
rect 32856 31526 32866 31578
rect 32866 31526 32912 31578
rect 32616 31524 32672 31526
rect 32696 31524 32752 31526
rect 32776 31524 32832 31526
rect 32856 31524 32912 31526
rect 32616 30490 32672 30492
rect 32696 30490 32752 30492
rect 32776 30490 32832 30492
rect 32856 30490 32912 30492
rect 32616 30438 32662 30490
rect 32662 30438 32672 30490
rect 32696 30438 32726 30490
rect 32726 30438 32738 30490
rect 32738 30438 32752 30490
rect 32776 30438 32790 30490
rect 32790 30438 32802 30490
rect 32802 30438 32832 30490
rect 32856 30438 32866 30490
rect 32866 30438 32912 30490
rect 32616 30436 32672 30438
rect 32696 30436 32752 30438
rect 32776 30436 32832 30438
rect 32856 30436 32912 30438
rect 32616 29402 32672 29404
rect 32696 29402 32752 29404
rect 32776 29402 32832 29404
rect 32856 29402 32912 29404
rect 32616 29350 32662 29402
rect 32662 29350 32672 29402
rect 32696 29350 32726 29402
rect 32726 29350 32738 29402
rect 32738 29350 32752 29402
rect 32776 29350 32790 29402
rect 32790 29350 32802 29402
rect 32802 29350 32832 29402
rect 32856 29350 32866 29402
rect 32866 29350 32912 29402
rect 32616 29348 32672 29350
rect 32696 29348 32752 29350
rect 32776 29348 32832 29350
rect 32856 29348 32912 29350
rect 32616 28314 32672 28316
rect 32696 28314 32752 28316
rect 32776 28314 32832 28316
rect 32856 28314 32912 28316
rect 32616 28262 32662 28314
rect 32662 28262 32672 28314
rect 32696 28262 32726 28314
rect 32726 28262 32738 28314
rect 32738 28262 32752 28314
rect 32776 28262 32790 28314
rect 32790 28262 32802 28314
rect 32802 28262 32832 28314
rect 32856 28262 32866 28314
rect 32866 28262 32912 28314
rect 32616 28260 32672 28262
rect 32696 28260 32752 28262
rect 32776 28260 32832 28262
rect 32856 28260 32912 28262
rect 32616 27226 32672 27228
rect 32696 27226 32752 27228
rect 32776 27226 32832 27228
rect 32856 27226 32912 27228
rect 32616 27174 32662 27226
rect 32662 27174 32672 27226
rect 32696 27174 32726 27226
rect 32726 27174 32738 27226
rect 32738 27174 32752 27226
rect 32776 27174 32790 27226
rect 32790 27174 32802 27226
rect 32802 27174 32832 27226
rect 32856 27174 32866 27226
rect 32866 27174 32912 27226
rect 32616 27172 32672 27174
rect 32696 27172 32752 27174
rect 32776 27172 32832 27174
rect 32856 27172 32912 27174
rect 32616 26138 32672 26140
rect 32696 26138 32752 26140
rect 32776 26138 32832 26140
rect 32856 26138 32912 26140
rect 32616 26086 32662 26138
rect 32662 26086 32672 26138
rect 32696 26086 32726 26138
rect 32726 26086 32738 26138
rect 32738 26086 32752 26138
rect 32776 26086 32790 26138
rect 32790 26086 32802 26138
rect 32802 26086 32832 26138
rect 32856 26086 32866 26138
rect 32866 26086 32912 26138
rect 32616 26084 32672 26086
rect 32696 26084 32752 26086
rect 32776 26084 32832 26086
rect 32856 26084 32912 26086
rect 32616 25050 32672 25052
rect 32696 25050 32752 25052
rect 32776 25050 32832 25052
rect 32856 25050 32912 25052
rect 32616 24998 32662 25050
rect 32662 24998 32672 25050
rect 32696 24998 32726 25050
rect 32726 24998 32738 25050
rect 32738 24998 32752 25050
rect 32776 24998 32790 25050
rect 32790 24998 32802 25050
rect 32802 24998 32832 25050
rect 32856 24998 32866 25050
rect 32866 24998 32912 25050
rect 32616 24996 32672 24998
rect 32696 24996 32752 24998
rect 32776 24996 32832 24998
rect 32856 24996 32912 24998
rect 32616 23962 32672 23964
rect 32696 23962 32752 23964
rect 32776 23962 32832 23964
rect 32856 23962 32912 23964
rect 32616 23910 32662 23962
rect 32662 23910 32672 23962
rect 32696 23910 32726 23962
rect 32726 23910 32738 23962
rect 32738 23910 32752 23962
rect 32776 23910 32790 23962
rect 32790 23910 32802 23962
rect 32802 23910 32832 23962
rect 32856 23910 32866 23962
rect 32866 23910 32912 23962
rect 32616 23908 32672 23910
rect 32696 23908 32752 23910
rect 32776 23908 32832 23910
rect 32856 23908 32912 23910
rect 32616 22874 32672 22876
rect 32696 22874 32752 22876
rect 32776 22874 32832 22876
rect 32856 22874 32912 22876
rect 32616 22822 32662 22874
rect 32662 22822 32672 22874
rect 32696 22822 32726 22874
rect 32726 22822 32738 22874
rect 32738 22822 32752 22874
rect 32776 22822 32790 22874
rect 32790 22822 32802 22874
rect 32802 22822 32832 22874
rect 32856 22822 32866 22874
rect 32866 22822 32912 22874
rect 32616 22820 32672 22822
rect 32696 22820 32752 22822
rect 32776 22820 32832 22822
rect 32856 22820 32912 22822
rect 32616 21786 32672 21788
rect 32696 21786 32752 21788
rect 32776 21786 32832 21788
rect 32856 21786 32912 21788
rect 32616 21734 32662 21786
rect 32662 21734 32672 21786
rect 32696 21734 32726 21786
rect 32726 21734 32738 21786
rect 32738 21734 32752 21786
rect 32776 21734 32790 21786
rect 32790 21734 32802 21786
rect 32802 21734 32832 21786
rect 32856 21734 32866 21786
rect 32866 21734 32912 21786
rect 32616 21732 32672 21734
rect 32696 21732 32752 21734
rect 32776 21732 32832 21734
rect 32856 21732 32912 21734
rect 32616 20698 32672 20700
rect 32696 20698 32752 20700
rect 32776 20698 32832 20700
rect 32856 20698 32912 20700
rect 32616 20646 32662 20698
rect 32662 20646 32672 20698
rect 32696 20646 32726 20698
rect 32726 20646 32738 20698
rect 32738 20646 32752 20698
rect 32776 20646 32790 20698
rect 32790 20646 32802 20698
rect 32802 20646 32832 20698
rect 32856 20646 32866 20698
rect 32866 20646 32912 20698
rect 32616 20644 32672 20646
rect 32696 20644 32752 20646
rect 32776 20644 32832 20646
rect 32856 20644 32912 20646
rect 32616 19610 32672 19612
rect 32696 19610 32752 19612
rect 32776 19610 32832 19612
rect 32856 19610 32912 19612
rect 32616 19558 32662 19610
rect 32662 19558 32672 19610
rect 32696 19558 32726 19610
rect 32726 19558 32738 19610
rect 32738 19558 32752 19610
rect 32776 19558 32790 19610
rect 32790 19558 32802 19610
rect 32802 19558 32832 19610
rect 32856 19558 32866 19610
rect 32866 19558 32912 19610
rect 32616 19556 32672 19558
rect 32696 19556 32752 19558
rect 32776 19556 32832 19558
rect 32856 19556 32912 19558
rect 32616 18522 32672 18524
rect 32696 18522 32752 18524
rect 32776 18522 32832 18524
rect 32856 18522 32912 18524
rect 32616 18470 32662 18522
rect 32662 18470 32672 18522
rect 32696 18470 32726 18522
rect 32726 18470 32738 18522
rect 32738 18470 32752 18522
rect 32776 18470 32790 18522
rect 32790 18470 32802 18522
rect 32802 18470 32832 18522
rect 32856 18470 32866 18522
rect 32866 18470 32912 18522
rect 32616 18468 32672 18470
rect 32696 18468 32752 18470
rect 32776 18468 32832 18470
rect 32856 18468 32912 18470
rect 32616 17434 32672 17436
rect 32696 17434 32752 17436
rect 32776 17434 32832 17436
rect 32856 17434 32912 17436
rect 32616 17382 32662 17434
rect 32662 17382 32672 17434
rect 32696 17382 32726 17434
rect 32726 17382 32738 17434
rect 32738 17382 32752 17434
rect 32776 17382 32790 17434
rect 32790 17382 32802 17434
rect 32802 17382 32832 17434
rect 32856 17382 32866 17434
rect 32866 17382 32912 17434
rect 32616 17380 32672 17382
rect 32696 17380 32752 17382
rect 32776 17380 32832 17382
rect 32856 17380 32912 17382
rect 32616 16346 32672 16348
rect 32696 16346 32752 16348
rect 32776 16346 32832 16348
rect 32856 16346 32912 16348
rect 32616 16294 32662 16346
rect 32662 16294 32672 16346
rect 32696 16294 32726 16346
rect 32726 16294 32738 16346
rect 32738 16294 32752 16346
rect 32776 16294 32790 16346
rect 32790 16294 32802 16346
rect 32802 16294 32832 16346
rect 32856 16294 32866 16346
rect 32866 16294 32912 16346
rect 32616 16292 32672 16294
rect 32696 16292 32752 16294
rect 32776 16292 32832 16294
rect 32856 16292 32912 16294
rect 32616 15258 32672 15260
rect 32696 15258 32752 15260
rect 32776 15258 32832 15260
rect 32856 15258 32912 15260
rect 32616 15206 32662 15258
rect 32662 15206 32672 15258
rect 32696 15206 32726 15258
rect 32726 15206 32738 15258
rect 32738 15206 32752 15258
rect 32776 15206 32790 15258
rect 32790 15206 32802 15258
rect 32802 15206 32832 15258
rect 32856 15206 32866 15258
rect 32866 15206 32912 15258
rect 32616 15204 32672 15206
rect 32696 15204 32752 15206
rect 32776 15204 32832 15206
rect 32856 15204 32912 15206
rect 31956 13626 32012 13628
rect 32036 13626 32092 13628
rect 32116 13626 32172 13628
rect 32196 13626 32252 13628
rect 31956 13574 32002 13626
rect 32002 13574 32012 13626
rect 32036 13574 32066 13626
rect 32066 13574 32078 13626
rect 32078 13574 32092 13626
rect 32116 13574 32130 13626
rect 32130 13574 32142 13626
rect 32142 13574 32172 13626
rect 32196 13574 32206 13626
rect 32206 13574 32252 13626
rect 31956 13572 32012 13574
rect 32036 13572 32092 13574
rect 32116 13572 32172 13574
rect 32196 13572 32252 13574
rect 31956 12538 32012 12540
rect 32036 12538 32092 12540
rect 32116 12538 32172 12540
rect 32196 12538 32252 12540
rect 31956 12486 32002 12538
rect 32002 12486 32012 12538
rect 32036 12486 32066 12538
rect 32066 12486 32078 12538
rect 32078 12486 32092 12538
rect 32116 12486 32130 12538
rect 32130 12486 32142 12538
rect 32142 12486 32172 12538
rect 32196 12486 32206 12538
rect 32206 12486 32252 12538
rect 31956 12484 32012 12486
rect 32036 12484 32092 12486
rect 32116 12484 32172 12486
rect 32196 12484 32252 12486
rect 31956 11450 32012 11452
rect 32036 11450 32092 11452
rect 32116 11450 32172 11452
rect 32196 11450 32252 11452
rect 31956 11398 32002 11450
rect 32002 11398 32012 11450
rect 32036 11398 32066 11450
rect 32066 11398 32078 11450
rect 32078 11398 32092 11450
rect 32116 11398 32130 11450
rect 32130 11398 32142 11450
rect 32142 11398 32172 11450
rect 32196 11398 32206 11450
rect 32206 11398 32252 11450
rect 31956 11396 32012 11398
rect 32036 11396 32092 11398
rect 32116 11396 32172 11398
rect 32196 11396 32252 11398
rect 32616 14170 32672 14172
rect 32696 14170 32752 14172
rect 32776 14170 32832 14172
rect 32856 14170 32912 14172
rect 32616 14118 32662 14170
rect 32662 14118 32672 14170
rect 32696 14118 32726 14170
rect 32726 14118 32738 14170
rect 32738 14118 32752 14170
rect 32776 14118 32790 14170
rect 32790 14118 32802 14170
rect 32802 14118 32832 14170
rect 32856 14118 32866 14170
rect 32866 14118 32912 14170
rect 32616 14116 32672 14118
rect 32696 14116 32752 14118
rect 32776 14116 32832 14118
rect 32856 14116 32912 14118
rect 32616 13082 32672 13084
rect 32696 13082 32752 13084
rect 32776 13082 32832 13084
rect 32856 13082 32912 13084
rect 32616 13030 32662 13082
rect 32662 13030 32672 13082
rect 32696 13030 32726 13082
rect 32726 13030 32738 13082
rect 32738 13030 32752 13082
rect 32776 13030 32790 13082
rect 32790 13030 32802 13082
rect 32802 13030 32832 13082
rect 32856 13030 32866 13082
rect 32866 13030 32912 13082
rect 32616 13028 32672 13030
rect 32696 13028 32752 13030
rect 32776 13028 32832 13030
rect 32856 13028 32912 13030
rect 32616 11994 32672 11996
rect 32696 11994 32752 11996
rect 32776 11994 32832 11996
rect 32856 11994 32912 11996
rect 32616 11942 32662 11994
rect 32662 11942 32672 11994
rect 32696 11942 32726 11994
rect 32726 11942 32738 11994
rect 32738 11942 32752 11994
rect 32776 11942 32790 11994
rect 32790 11942 32802 11994
rect 32802 11942 32832 11994
rect 32856 11942 32866 11994
rect 32866 11942 32912 11994
rect 32616 11940 32672 11942
rect 32696 11940 32752 11942
rect 32776 11940 32832 11942
rect 32856 11940 32912 11942
rect 31956 10362 32012 10364
rect 32036 10362 32092 10364
rect 32116 10362 32172 10364
rect 32196 10362 32252 10364
rect 31956 10310 32002 10362
rect 32002 10310 32012 10362
rect 32036 10310 32066 10362
rect 32066 10310 32078 10362
rect 32078 10310 32092 10362
rect 32116 10310 32130 10362
rect 32130 10310 32142 10362
rect 32142 10310 32172 10362
rect 32196 10310 32206 10362
rect 32206 10310 32252 10362
rect 31956 10308 32012 10310
rect 32036 10308 32092 10310
rect 32116 10308 32172 10310
rect 32196 10308 32252 10310
rect 32616 10906 32672 10908
rect 32696 10906 32752 10908
rect 32776 10906 32832 10908
rect 32856 10906 32912 10908
rect 32616 10854 32662 10906
rect 32662 10854 32672 10906
rect 32696 10854 32726 10906
rect 32726 10854 32738 10906
rect 32738 10854 32752 10906
rect 32776 10854 32790 10906
rect 32790 10854 32802 10906
rect 32802 10854 32832 10906
rect 32856 10854 32866 10906
rect 32866 10854 32912 10906
rect 32616 10852 32672 10854
rect 32696 10852 32752 10854
rect 32776 10852 32832 10854
rect 32856 10852 32912 10854
rect 32616 9818 32672 9820
rect 32696 9818 32752 9820
rect 32776 9818 32832 9820
rect 32856 9818 32912 9820
rect 32616 9766 32662 9818
rect 32662 9766 32672 9818
rect 32696 9766 32726 9818
rect 32726 9766 32738 9818
rect 32738 9766 32752 9818
rect 32776 9766 32790 9818
rect 32790 9766 32802 9818
rect 32802 9766 32832 9818
rect 32856 9766 32866 9818
rect 32866 9766 32912 9818
rect 32616 9764 32672 9766
rect 32696 9764 32752 9766
rect 32776 9764 32832 9766
rect 32856 9764 32912 9766
rect 31956 9274 32012 9276
rect 32036 9274 32092 9276
rect 32116 9274 32172 9276
rect 32196 9274 32252 9276
rect 31956 9222 32002 9274
rect 32002 9222 32012 9274
rect 32036 9222 32066 9274
rect 32066 9222 32078 9274
rect 32078 9222 32092 9274
rect 32116 9222 32130 9274
rect 32130 9222 32142 9274
rect 32142 9222 32172 9274
rect 32196 9222 32206 9274
rect 32206 9222 32252 9274
rect 31956 9220 32012 9222
rect 32036 9220 32092 9222
rect 32116 9220 32172 9222
rect 32196 9220 32252 9222
rect 32616 8730 32672 8732
rect 32696 8730 32752 8732
rect 32776 8730 32832 8732
rect 32856 8730 32912 8732
rect 32616 8678 32662 8730
rect 32662 8678 32672 8730
rect 32696 8678 32726 8730
rect 32726 8678 32738 8730
rect 32738 8678 32752 8730
rect 32776 8678 32790 8730
rect 32790 8678 32802 8730
rect 32802 8678 32832 8730
rect 32856 8678 32866 8730
rect 32866 8678 32912 8730
rect 32616 8676 32672 8678
rect 32696 8676 32752 8678
rect 32776 8676 32832 8678
rect 32856 8676 32912 8678
rect 31956 8186 32012 8188
rect 32036 8186 32092 8188
rect 32116 8186 32172 8188
rect 32196 8186 32252 8188
rect 31956 8134 32002 8186
rect 32002 8134 32012 8186
rect 32036 8134 32066 8186
rect 32066 8134 32078 8186
rect 32078 8134 32092 8186
rect 32116 8134 32130 8186
rect 32130 8134 32142 8186
rect 32142 8134 32172 8186
rect 32196 8134 32206 8186
rect 32206 8134 32252 8186
rect 31956 8132 32012 8134
rect 32036 8132 32092 8134
rect 32116 8132 32172 8134
rect 32196 8132 32252 8134
rect 32616 7642 32672 7644
rect 32696 7642 32752 7644
rect 32776 7642 32832 7644
rect 32856 7642 32912 7644
rect 32616 7590 32662 7642
rect 32662 7590 32672 7642
rect 32696 7590 32726 7642
rect 32726 7590 32738 7642
rect 32738 7590 32752 7642
rect 32776 7590 32790 7642
rect 32790 7590 32802 7642
rect 32802 7590 32832 7642
rect 32856 7590 32866 7642
rect 32866 7590 32912 7642
rect 32616 7588 32672 7590
rect 32696 7588 32752 7590
rect 32776 7588 32832 7590
rect 32856 7588 32912 7590
rect 31956 7098 32012 7100
rect 32036 7098 32092 7100
rect 32116 7098 32172 7100
rect 32196 7098 32252 7100
rect 31956 7046 32002 7098
rect 32002 7046 32012 7098
rect 32036 7046 32066 7098
rect 32066 7046 32078 7098
rect 32078 7046 32092 7098
rect 32116 7046 32130 7098
rect 32130 7046 32142 7098
rect 32142 7046 32172 7098
rect 32196 7046 32206 7098
rect 32206 7046 32252 7098
rect 31956 7044 32012 7046
rect 32036 7044 32092 7046
rect 32116 7044 32172 7046
rect 32196 7044 32252 7046
rect 32616 6554 32672 6556
rect 32696 6554 32752 6556
rect 32776 6554 32832 6556
rect 32856 6554 32912 6556
rect 32616 6502 32662 6554
rect 32662 6502 32672 6554
rect 32696 6502 32726 6554
rect 32726 6502 32738 6554
rect 32738 6502 32752 6554
rect 32776 6502 32790 6554
rect 32790 6502 32802 6554
rect 32802 6502 32832 6554
rect 32856 6502 32866 6554
rect 32866 6502 32912 6554
rect 32616 6500 32672 6502
rect 32696 6500 32752 6502
rect 32776 6500 32832 6502
rect 32856 6500 32912 6502
rect 31956 6010 32012 6012
rect 32036 6010 32092 6012
rect 32116 6010 32172 6012
rect 32196 6010 32252 6012
rect 31956 5958 32002 6010
rect 32002 5958 32012 6010
rect 32036 5958 32066 6010
rect 32066 5958 32078 6010
rect 32078 5958 32092 6010
rect 32116 5958 32130 6010
rect 32130 5958 32142 6010
rect 32142 5958 32172 6010
rect 32196 5958 32206 6010
rect 32206 5958 32252 6010
rect 31956 5956 32012 5958
rect 32036 5956 32092 5958
rect 32116 5956 32172 5958
rect 32196 5956 32252 5958
rect 32616 5466 32672 5468
rect 32696 5466 32752 5468
rect 32776 5466 32832 5468
rect 32856 5466 32912 5468
rect 32616 5414 32662 5466
rect 32662 5414 32672 5466
rect 32696 5414 32726 5466
rect 32726 5414 32738 5466
rect 32738 5414 32752 5466
rect 32776 5414 32790 5466
rect 32790 5414 32802 5466
rect 32802 5414 32832 5466
rect 32856 5414 32866 5466
rect 32866 5414 32912 5466
rect 32616 5412 32672 5414
rect 32696 5412 32752 5414
rect 32776 5412 32832 5414
rect 32856 5412 32912 5414
rect 31956 4922 32012 4924
rect 32036 4922 32092 4924
rect 32116 4922 32172 4924
rect 32196 4922 32252 4924
rect 31956 4870 32002 4922
rect 32002 4870 32012 4922
rect 32036 4870 32066 4922
rect 32066 4870 32078 4922
rect 32078 4870 32092 4922
rect 32116 4870 32130 4922
rect 32130 4870 32142 4922
rect 32142 4870 32172 4922
rect 32196 4870 32206 4922
rect 32206 4870 32252 4922
rect 31956 4868 32012 4870
rect 32036 4868 32092 4870
rect 32116 4868 32172 4870
rect 32196 4868 32252 4870
rect 32616 4378 32672 4380
rect 32696 4378 32752 4380
rect 32776 4378 32832 4380
rect 32856 4378 32912 4380
rect 32616 4326 32662 4378
rect 32662 4326 32672 4378
rect 32696 4326 32726 4378
rect 32726 4326 32738 4378
rect 32738 4326 32752 4378
rect 32776 4326 32790 4378
rect 32790 4326 32802 4378
rect 32802 4326 32832 4378
rect 32856 4326 32866 4378
rect 32866 4326 32912 4378
rect 32616 4324 32672 4326
rect 32696 4324 32752 4326
rect 32776 4324 32832 4326
rect 32856 4324 32912 4326
rect 31956 3834 32012 3836
rect 32036 3834 32092 3836
rect 32116 3834 32172 3836
rect 32196 3834 32252 3836
rect 31956 3782 32002 3834
rect 32002 3782 32012 3834
rect 32036 3782 32066 3834
rect 32066 3782 32078 3834
rect 32078 3782 32092 3834
rect 32116 3782 32130 3834
rect 32130 3782 32142 3834
rect 32142 3782 32172 3834
rect 32196 3782 32206 3834
rect 32206 3782 32252 3834
rect 31956 3780 32012 3782
rect 32036 3780 32092 3782
rect 32116 3780 32172 3782
rect 32196 3780 32252 3782
rect 32616 3290 32672 3292
rect 32696 3290 32752 3292
rect 32776 3290 32832 3292
rect 32856 3290 32912 3292
rect 32616 3238 32662 3290
rect 32662 3238 32672 3290
rect 32696 3238 32726 3290
rect 32726 3238 32738 3290
rect 32738 3238 32752 3290
rect 32776 3238 32790 3290
rect 32790 3238 32802 3290
rect 32802 3238 32832 3290
rect 32856 3238 32866 3290
rect 32866 3238 32912 3290
rect 32616 3236 32672 3238
rect 32696 3236 32752 3238
rect 32776 3236 32832 3238
rect 32856 3236 32912 3238
rect 34702 51040 34758 51096
rect 26956 2746 27012 2748
rect 27036 2746 27092 2748
rect 27116 2746 27172 2748
rect 27196 2746 27252 2748
rect 26956 2694 27002 2746
rect 27002 2694 27012 2746
rect 27036 2694 27066 2746
rect 27066 2694 27078 2746
rect 27078 2694 27092 2746
rect 27116 2694 27130 2746
rect 27130 2694 27142 2746
rect 27142 2694 27172 2746
rect 27196 2694 27206 2746
rect 27206 2694 27252 2746
rect 26956 2692 27012 2694
rect 27036 2692 27092 2694
rect 27116 2692 27172 2694
rect 27196 2692 27252 2694
rect 31956 2746 32012 2748
rect 32036 2746 32092 2748
rect 32116 2746 32172 2748
rect 32196 2746 32252 2748
rect 31956 2694 32002 2746
rect 32002 2694 32012 2746
rect 32036 2694 32066 2746
rect 32066 2694 32078 2746
rect 32078 2694 32092 2746
rect 32116 2694 32130 2746
rect 32130 2694 32142 2746
rect 32142 2694 32172 2746
rect 32196 2694 32206 2746
rect 32206 2694 32252 2746
rect 31956 2692 32012 2694
rect 32036 2692 32092 2694
rect 32116 2692 32172 2694
rect 32196 2692 32252 2694
rect 35254 61648 35310 61704
rect 36956 69114 37012 69116
rect 37036 69114 37092 69116
rect 37116 69114 37172 69116
rect 37196 69114 37252 69116
rect 36956 69062 37002 69114
rect 37002 69062 37012 69114
rect 37036 69062 37066 69114
rect 37066 69062 37078 69114
rect 37078 69062 37092 69114
rect 37116 69062 37130 69114
rect 37130 69062 37142 69114
rect 37142 69062 37172 69114
rect 37196 69062 37206 69114
rect 37206 69062 37252 69114
rect 36956 69060 37012 69062
rect 37036 69060 37092 69062
rect 37116 69060 37172 69062
rect 37196 69060 37252 69062
rect 37616 68570 37672 68572
rect 37696 68570 37752 68572
rect 37776 68570 37832 68572
rect 37856 68570 37912 68572
rect 37616 68518 37662 68570
rect 37662 68518 37672 68570
rect 37696 68518 37726 68570
rect 37726 68518 37738 68570
rect 37738 68518 37752 68570
rect 37776 68518 37790 68570
rect 37790 68518 37802 68570
rect 37802 68518 37832 68570
rect 37856 68518 37866 68570
rect 37866 68518 37912 68570
rect 37616 68516 37672 68518
rect 37696 68516 37752 68518
rect 37776 68516 37832 68518
rect 37856 68516 37912 68518
rect 36956 68026 37012 68028
rect 37036 68026 37092 68028
rect 37116 68026 37172 68028
rect 37196 68026 37252 68028
rect 36956 67974 37002 68026
rect 37002 67974 37012 68026
rect 37036 67974 37066 68026
rect 37066 67974 37078 68026
rect 37078 67974 37092 68026
rect 37116 67974 37130 68026
rect 37130 67974 37142 68026
rect 37142 67974 37172 68026
rect 37196 67974 37206 68026
rect 37206 67974 37252 68026
rect 36956 67972 37012 67974
rect 37036 67972 37092 67974
rect 37116 67972 37172 67974
rect 37196 67972 37252 67974
rect 38014 67804 38016 67824
rect 38016 67804 38068 67824
rect 38068 67804 38070 67824
rect 38014 67768 38070 67804
rect 37094 67668 37096 67688
rect 37096 67668 37148 67688
rect 37148 67668 37150 67688
rect 37094 67632 37150 67668
rect 35346 15020 35402 15056
rect 35346 15000 35348 15020
rect 35348 15000 35400 15020
rect 35400 15000 35402 15020
rect 37616 67482 37672 67484
rect 37696 67482 37752 67484
rect 37776 67482 37832 67484
rect 37856 67482 37912 67484
rect 37616 67430 37662 67482
rect 37662 67430 37672 67482
rect 37696 67430 37726 67482
rect 37726 67430 37738 67482
rect 37738 67430 37752 67482
rect 37776 67430 37790 67482
rect 37790 67430 37802 67482
rect 37802 67430 37832 67482
rect 37856 67430 37866 67482
rect 37866 67430 37912 67482
rect 37616 67428 37672 67430
rect 37696 67428 37752 67430
rect 37776 67428 37832 67430
rect 37856 67428 37912 67430
rect 36956 66938 37012 66940
rect 37036 66938 37092 66940
rect 37116 66938 37172 66940
rect 37196 66938 37252 66940
rect 36956 66886 37002 66938
rect 37002 66886 37012 66938
rect 37036 66886 37066 66938
rect 37066 66886 37078 66938
rect 37078 66886 37092 66938
rect 37116 66886 37130 66938
rect 37130 66886 37142 66938
rect 37142 66886 37172 66938
rect 37196 66886 37206 66938
rect 37206 66886 37252 66938
rect 36956 66884 37012 66886
rect 37036 66884 37092 66886
rect 37116 66884 37172 66886
rect 37196 66884 37252 66886
rect 36956 65850 37012 65852
rect 37036 65850 37092 65852
rect 37116 65850 37172 65852
rect 37196 65850 37252 65852
rect 36956 65798 37002 65850
rect 37002 65798 37012 65850
rect 37036 65798 37066 65850
rect 37066 65798 37078 65850
rect 37078 65798 37092 65850
rect 37116 65798 37130 65850
rect 37130 65798 37142 65850
rect 37142 65798 37172 65850
rect 37196 65798 37206 65850
rect 37206 65798 37252 65850
rect 36956 65796 37012 65798
rect 37036 65796 37092 65798
rect 37116 65796 37172 65798
rect 37196 65796 37252 65798
rect 37616 66394 37672 66396
rect 37696 66394 37752 66396
rect 37776 66394 37832 66396
rect 37856 66394 37912 66396
rect 37616 66342 37662 66394
rect 37662 66342 37672 66394
rect 37696 66342 37726 66394
rect 37726 66342 37738 66394
rect 37738 66342 37752 66394
rect 37776 66342 37790 66394
rect 37790 66342 37802 66394
rect 37802 66342 37832 66394
rect 37856 66342 37866 66394
rect 37866 66342 37912 66394
rect 37616 66340 37672 66342
rect 37696 66340 37752 66342
rect 37776 66340 37832 66342
rect 37856 66340 37912 66342
rect 37616 65306 37672 65308
rect 37696 65306 37752 65308
rect 37776 65306 37832 65308
rect 37856 65306 37912 65308
rect 37616 65254 37662 65306
rect 37662 65254 37672 65306
rect 37696 65254 37726 65306
rect 37726 65254 37738 65306
rect 37738 65254 37752 65306
rect 37776 65254 37790 65306
rect 37790 65254 37802 65306
rect 37802 65254 37832 65306
rect 37856 65254 37866 65306
rect 37866 65254 37912 65306
rect 37616 65252 37672 65254
rect 37696 65252 37752 65254
rect 37776 65252 37832 65254
rect 37856 65252 37912 65254
rect 36956 64762 37012 64764
rect 37036 64762 37092 64764
rect 37116 64762 37172 64764
rect 37196 64762 37252 64764
rect 36956 64710 37002 64762
rect 37002 64710 37012 64762
rect 37036 64710 37066 64762
rect 37066 64710 37078 64762
rect 37078 64710 37092 64762
rect 37116 64710 37130 64762
rect 37130 64710 37142 64762
rect 37142 64710 37172 64762
rect 37196 64710 37206 64762
rect 37206 64710 37252 64762
rect 36956 64708 37012 64710
rect 37036 64708 37092 64710
rect 37116 64708 37172 64710
rect 37196 64708 37252 64710
rect 37616 64218 37672 64220
rect 37696 64218 37752 64220
rect 37776 64218 37832 64220
rect 37856 64218 37912 64220
rect 37616 64166 37662 64218
rect 37662 64166 37672 64218
rect 37696 64166 37726 64218
rect 37726 64166 37738 64218
rect 37738 64166 37752 64218
rect 37776 64166 37790 64218
rect 37790 64166 37802 64218
rect 37802 64166 37832 64218
rect 37856 64166 37866 64218
rect 37866 64166 37912 64218
rect 37616 64164 37672 64166
rect 37696 64164 37752 64166
rect 37776 64164 37832 64166
rect 37856 64164 37912 64166
rect 36956 63674 37012 63676
rect 37036 63674 37092 63676
rect 37116 63674 37172 63676
rect 37196 63674 37252 63676
rect 36956 63622 37002 63674
rect 37002 63622 37012 63674
rect 37036 63622 37066 63674
rect 37066 63622 37078 63674
rect 37078 63622 37092 63674
rect 37116 63622 37130 63674
rect 37130 63622 37142 63674
rect 37142 63622 37172 63674
rect 37196 63622 37206 63674
rect 37206 63622 37252 63674
rect 36956 63620 37012 63622
rect 37036 63620 37092 63622
rect 37116 63620 37172 63622
rect 37196 63620 37252 63622
rect 36956 62586 37012 62588
rect 37036 62586 37092 62588
rect 37116 62586 37172 62588
rect 37196 62586 37252 62588
rect 36956 62534 37002 62586
rect 37002 62534 37012 62586
rect 37036 62534 37066 62586
rect 37066 62534 37078 62586
rect 37078 62534 37092 62586
rect 37116 62534 37130 62586
rect 37130 62534 37142 62586
rect 37142 62534 37172 62586
rect 37196 62534 37206 62586
rect 37206 62534 37252 62586
rect 36956 62532 37012 62534
rect 37036 62532 37092 62534
rect 37116 62532 37172 62534
rect 37196 62532 37252 62534
rect 36956 61498 37012 61500
rect 37036 61498 37092 61500
rect 37116 61498 37172 61500
rect 37196 61498 37252 61500
rect 36956 61446 37002 61498
rect 37002 61446 37012 61498
rect 37036 61446 37066 61498
rect 37066 61446 37078 61498
rect 37078 61446 37092 61498
rect 37116 61446 37130 61498
rect 37130 61446 37142 61498
rect 37142 61446 37172 61498
rect 37196 61446 37206 61498
rect 37206 61446 37252 61498
rect 36956 61444 37012 61446
rect 37036 61444 37092 61446
rect 37116 61444 37172 61446
rect 37196 61444 37252 61446
rect 36956 60410 37012 60412
rect 37036 60410 37092 60412
rect 37116 60410 37172 60412
rect 37196 60410 37252 60412
rect 36956 60358 37002 60410
rect 37002 60358 37012 60410
rect 37036 60358 37066 60410
rect 37066 60358 37078 60410
rect 37078 60358 37092 60410
rect 37116 60358 37130 60410
rect 37130 60358 37142 60410
rect 37142 60358 37172 60410
rect 37196 60358 37206 60410
rect 37206 60358 37252 60410
rect 36956 60356 37012 60358
rect 37036 60356 37092 60358
rect 37116 60356 37172 60358
rect 37196 60356 37252 60358
rect 36956 59322 37012 59324
rect 37036 59322 37092 59324
rect 37116 59322 37172 59324
rect 37196 59322 37252 59324
rect 36956 59270 37002 59322
rect 37002 59270 37012 59322
rect 37036 59270 37066 59322
rect 37066 59270 37078 59322
rect 37078 59270 37092 59322
rect 37116 59270 37130 59322
rect 37130 59270 37142 59322
rect 37142 59270 37172 59322
rect 37196 59270 37206 59322
rect 37206 59270 37252 59322
rect 36956 59268 37012 59270
rect 37036 59268 37092 59270
rect 37116 59268 37172 59270
rect 37196 59268 37252 59270
rect 36956 58234 37012 58236
rect 37036 58234 37092 58236
rect 37116 58234 37172 58236
rect 37196 58234 37252 58236
rect 36956 58182 37002 58234
rect 37002 58182 37012 58234
rect 37036 58182 37066 58234
rect 37066 58182 37078 58234
rect 37078 58182 37092 58234
rect 37116 58182 37130 58234
rect 37130 58182 37142 58234
rect 37142 58182 37172 58234
rect 37196 58182 37206 58234
rect 37206 58182 37252 58234
rect 36956 58180 37012 58182
rect 37036 58180 37092 58182
rect 37116 58180 37172 58182
rect 37196 58180 37252 58182
rect 36956 57146 37012 57148
rect 37036 57146 37092 57148
rect 37116 57146 37172 57148
rect 37196 57146 37252 57148
rect 36956 57094 37002 57146
rect 37002 57094 37012 57146
rect 37036 57094 37066 57146
rect 37066 57094 37078 57146
rect 37078 57094 37092 57146
rect 37116 57094 37130 57146
rect 37130 57094 37142 57146
rect 37142 57094 37172 57146
rect 37196 57094 37206 57146
rect 37206 57094 37252 57146
rect 36956 57092 37012 57094
rect 37036 57092 37092 57094
rect 37116 57092 37172 57094
rect 37196 57092 37252 57094
rect 36956 56058 37012 56060
rect 37036 56058 37092 56060
rect 37116 56058 37172 56060
rect 37196 56058 37252 56060
rect 36956 56006 37002 56058
rect 37002 56006 37012 56058
rect 37036 56006 37066 56058
rect 37066 56006 37078 56058
rect 37078 56006 37092 56058
rect 37116 56006 37130 56058
rect 37130 56006 37142 56058
rect 37142 56006 37172 56058
rect 37196 56006 37206 56058
rect 37206 56006 37252 56058
rect 36956 56004 37012 56006
rect 37036 56004 37092 56006
rect 37116 56004 37172 56006
rect 37196 56004 37252 56006
rect 37616 63130 37672 63132
rect 37696 63130 37752 63132
rect 37776 63130 37832 63132
rect 37856 63130 37912 63132
rect 37616 63078 37662 63130
rect 37662 63078 37672 63130
rect 37696 63078 37726 63130
rect 37726 63078 37738 63130
rect 37738 63078 37752 63130
rect 37776 63078 37790 63130
rect 37790 63078 37802 63130
rect 37802 63078 37832 63130
rect 37856 63078 37866 63130
rect 37866 63078 37912 63130
rect 37616 63076 37672 63078
rect 37696 63076 37752 63078
rect 37776 63076 37832 63078
rect 37856 63076 37912 63078
rect 37616 62042 37672 62044
rect 37696 62042 37752 62044
rect 37776 62042 37832 62044
rect 37856 62042 37912 62044
rect 37616 61990 37662 62042
rect 37662 61990 37672 62042
rect 37696 61990 37726 62042
rect 37726 61990 37738 62042
rect 37738 61990 37752 62042
rect 37776 61990 37790 62042
rect 37790 61990 37802 62042
rect 37802 61990 37832 62042
rect 37856 61990 37866 62042
rect 37866 61990 37912 62042
rect 37616 61988 37672 61990
rect 37696 61988 37752 61990
rect 37776 61988 37832 61990
rect 37856 61988 37912 61990
rect 37616 60954 37672 60956
rect 37696 60954 37752 60956
rect 37776 60954 37832 60956
rect 37856 60954 37912 60956
rect 37616 60902 37662 60954
rect 37662 60902 37672 60954
rect 37696 60902 37726 60954
rect 37726 60902 37738 60954
rect 37738 60902 37752 60954
rect 37776 60902 37790 60954
rect 37790 60902 37802 60954
rect 37802 60902 37832 60954
rect 37856 60902 37866 60954
rect 37866 60902 37912 60954
rect 37616 60900 37672 60902
rect 37696 60900 37752 60902
rect 37776 60900 37832 60902
rect 37856 60900 37912 60902
rect 37616 59866 37672 59868
rect 37696 59866 37752 59868
rect 37776 59866 37832 59868
rect 37856 59866 37912 59868
rect 37616 59814 37662 59866
rect 37662 59814 37672 59866
rect 37696 59814 37726 59866
rect 37726 59814 37738 59866
rect 37738 59814 37752 59866
rect 37776 59814 37790 59866
rect 37790 59814 37802 59866
rect 37802 59814 37832 59866
rect 37856 59814 37866 59866
rect 37866 59814 37912 59866
rect 37616 59812 37672 59814
rect 37696 59812 37752 59814
rect 37776 59812 37832 59814
rect 37856 59812 37912 59814
rect 37616 58778 37672 58780
rect 37696 58778 37752 58780
rect 37776 58778 37832 58780
rect 37856 58778 37912 58780
rect 37616 58726 37662 58778
rect 37662 58726 37672 58778
rect 37696 58726 37726 58778
rect 37726 58726 37738 58778
rect 37738 58726 37752 58778
rect 37776 58726 37790 58778
rect 37790 58726 37802 58778
rect 37802 58726 37832 58778
rect 37856 58726 37866 58778
rect 37866 58726 37912 58778
rect 37616 58724 37672 58726
rect 37696 58724 37752 58726
rect 37776 58724 37832 58726
rect 37856 58724 37912 58726
rect 37616 57690 37672 57692
rect 37696 57690 37752 57692
rect 37776 57690 37832 57692
rect 37856 57690 37912 57692
rect 37616 57638 37662 57690
rect 37662 57638 37672 57690
rect 37696 57638 37726 57690
rect 37726 57638 37738 57690
rect 37738 57638 37752 57690
rect 37776 57638 37790 57690
rect 37790 57638 37802 57690
rect 37802 57638 37832 57690
rect 37856 57638 37866 57690
rect 37866 57638 37912 57690
rect 37616 57636 37672 57638
rect 37696 57636 37752 57638
rect 37776 57636 37832 57638
rect 37856 57636 37912 57638
rect 37616 56602 37672 56604
rect 37696 56602 37752 56604
rect 37776 56602 37832 56604
rect 37856 56602 37912 56604
rect 37616 56550 37662 56602
rect 37662 56550 37672 56602
rect 37696 56550 37726 56602
rect 37726 56550 37738 56602
rect 37738 56550 37752 56602
rect 37776 56550 37790 56602
rect 37790 56550 37802 56602
rect 37802 56550 37832 56602
rect 37856 56550 37866 56602
rect 37866 56550 37912 56602
rect 37616 56548 37672 56550
rect 37696 56548 37752 56550
rect 37776 56548 37832 56550
rect 37856 56548 37912 56550
rect 37616 55514 37672 55516
rect 37696 55514 37752 55516
rect 37776 55514 37832 55516
rect 37856 55514 37912 55516
rect 37616 55462 37662 55514
rect 37662 55462 37672 55514
rect 37696 55462 37726 55514
rect 37726 55462 37738 55514
rect 37738 55462 37752 55514
rect 37776 55462 37790 55514
rect 37790 55462 37802 55514
rect 37802 55462 37832 55514
rect 37856 55462 37866 55514
rect 37866 55462 37912 55514
rect 37616 55460 37672 55462
rect 37696 55460 37752 55462
rect 37776 55460 37832 55462
rect 37856 55460 37912 55462
rect 36956 54970 37012 54972
rect 37036 54970 37092 54972
rect 37116 54970 37172 54972
rect 37196 54970 37252 54972
rect 36956 54918 37002 54970
rect 37002 54918 37012 54970
rect 37036 54918 37066 54970
rect 37066 54918 37078 54970
rect 37078 54918 37092 54970
rect 37116 54918 37130 54970
rect 37130 54918 37142 54970
rect 37142 54918 37172 54970
rect 37196 54918 37206 54970
rect 37206 54918 37252 54970
rect 36956 54916 37012 54918
rect 37036 54916 37092 54918
rect 37116 54916 37172 54918
rect 37196 54916 37252 54918
rect 36956 53882 37012 53884
rect 37036 53882 37092 53884
rect 37116 53882 37172 53884
rect 37196 53882 37252 53884
rect 36956 53830 37002 53882
rect 37002 53830 37012 53882
rect 37036 53830 37066 53882
rect 37066 53830 37078 53882
rect 37078 53830 37092 53882
rect 37116 53830 37130 53882
rect 37130 53830 37142 53882
rect 37142 53830 37172 53882
rect 37196 53830 37206 53882
rect 37206 53830 37252 53882
rect 36956 53828 37012 53830
rect 37036 53828 37092 53830
rect 37116 53828 37172 53830
rect 37196 53828 37252 53830
rect 36956 52794 37012 52796
rect 37036 52794 37092 52796
rect 37116 52794 37172 52796
rect 37196 52794 37252 52796
rect 36956 52742 37002 52794
rect 37002 52742 37012 52794
rect 37036 52742 37066 52794
rect 37066 52742 37078 52794
rect 37078 52742 37092 52794
rect 37116 52742 37130 52794
rect 37130 52742 37142 52794
rect 37142 52742 37172 52794
rect 37196 52742 37206 52794
rect 37206 52742 37252 52794
rect 36956 52740 37012 52742
rect 37036 52740 37092 52742
rect 37116 52740 37172 52742
rect 37196 52740 37252 52742
rect 36956 51706 37012 51708
rect 37036 51706 37092 51708
rect 37116 51706 37172 51708
rect 37196 51706 37252 51708
rect 36956 51654 37002 51706
rect 37002 51654 37012 51706
rect 37036 51654 37066 51706
rect 37066 51654 37078 51706
rect 37078 51654 37092 51706
rect 37116 51654 37130 51706
rect 37130 51654 37142 51706
rect 37142 51654 37172 51706
rect 37196 51654 37206 51706
rect 37206 51654 37252 51706
rect 36956 51652 37012 51654
rect 37036 51652 37092 51654
rect 37116 51652 37172 51654
rect 37196 51652 37252 51654
rect 36956 50618 37012 50620
rect 37036 50618 37092 50620
rect 37116 50618 37172 50620
rect 37196 50618 37252 50620
rect 36956 50566 37002 50618
rect 37002 50566 37012 50618
rect 37036 50566 37066 50618
rect 37066 50566 37078 50618
rect 37078 50566 37092 50618
rect 37116 50566 37130 50618
rect 37130 50566 37142 50618
rect 37142 50566 37172 50618
rect 37196 50566 37206 50618
rect 37206 50566 37252 50618
rect 36956 50564 37012 50566
rect 37036 50564 37092 50566
rect 37116 50564 37172 50566
rect 37196 50564 37252 50566
rect 36956 49530 37012 49532
rect 37036 49530 37092 49532
rect 37116 49530 37172 49532
rect 37196 49530 37252 49532
rect 36956 49478 37002 49530
rect 37002 49478 37012 49530
rect 37036 49478 37066 49530
rect 37066 49478 37078 49530
rect 37078 49478 37092 49530
rect 37116 49478 37130 49530
rect 37130 49478 37142 49530
rect 37142 49478 37172 49530
rect 37196 49478 37206 49530
rect 37206 49478 37252 49530
rect 36956 49476 37012 49478
rect 37036 49476 37092 49478
rect 37116 49476 37172 49478
rect 37196 49476 37252 49478
rect 36956 48442 37012 48444
rect 37036 48442 37092 48444
rect 37116 48442 37172 48444
rect 37196 48442 37252 48444
rect 36956 48390 37002 48442
rect 37002 48390 37012 48442
rect 37036 48390 37066 48442
rect 37066 48390 37078 48442
rect 37078 48390 37092 48442
rect 37116 48390 37130 48442
rect 37130 48390 37142 48442
rect 37142 48390 37172 48442
rect 37196 48390 37206 48442
rect 37206 48390 37252 48442
rect 36956 48388 37012 48390
rect 37036 48388 37092 48390
rect 37116 48388 37172 48390
rect 37196 48388 37252 48390
rect 36956 47354 37012 47356
rect 37036 47354 37092 47356
rect 37116 47354 37172 47356
rect 37196 47354 37252 47356
rect 36956 47302 37002 47354
rect 37002 47302 37012 47354
rect 37036 47302 37066 47354
rect 37066 47302 37078 47354
rect 37078 47302 37092 47354
rect 37116 47302 37130 47354
rect 37130 47302 37142 47354
rect 37142 47302 37172 47354
rect 37196 47302 37206 47354
rect 37206 47302 37252 47354
rect 36956 47300 37012 47302
rect 37036 47300 37092 47302
rect 37116 47300 37172 47302
rect 37196 47300 37252 47302
rect 36956 46266 37012 46268
rect 37036 46266 37092 46268
rect 37116 46266 37172 46268
rect 37196 46266 37252 46268
rect 36956 46214 37002 46266
rect 37002 46214 37012 46266
rect 37036 46214 37066 46266
rect 37066 46214 37078 46266
rect 37078 46214 37092 46266
rect 37116 46214 37130 46266
rect 37130 46214 37142 46266
rect 37142 46214 37172 46266
rect 37196 46214 37206 46266
rect 37206 46214 37252 46266
rect 36956 46212 37012 46214
rect 37036 46212 37092 46214
rect 37116 46212 37172 46214
rect 37196 46212 37252 46214
rect 36956 45178 37012 45180
rect 37036 45178 37092 45180
rect 37116 45178 37172 45180
rect 37196 45178 37252 45180
rect 36956 45126 37002 45178
rect 37002 45126 37012 45178
rect 37036 45126 37066 45178
rect 37066 45126 37078 45178
rect 37078 45126 37092 45178
rect 37116 45126 37130 45178
rect 37130 45126 37142 45178
rect 37142 45126 37172 45178
rect 37196 45126 37206 45178
rect 37206 45126 37252 45178
rect 36956 45124 37012 45126
rect 37036 45124 37092 45126
rect 37116 45124 37172 45126
rect 37196 45124 37252 45126
rect 36956 44090 37012 44092
rect 37036 44090 37092 44092
rect 37116 44090 37172 44092
rect 37196 44090 37252 44092
rect 36956 44038 37002 44090
rect 37002 44038 37012 44090
rect 37036 44038 37066 44090
rect 37066 44038 37078 44090
rect 37078 44038 37092 44090
rect 37116 44038 37130 44090
rect 37130 44038 37142 44090
rect 37142 44038 37172 44090
rect 37196 44038 37206 44090
rect 37206 44038 37252 44090
rect 36956 44036 37012 44038
rect 37036 44036 37092 44038
rect 37116 44036 37172 44038
rect 37196 44036 37252 44038
rect 36956 43002 37012 43004
rect 37036 43002 37092 43004
rect 37116 43002 37172 43004
rect 37196 43002 37252 43004
rect 36956 42950 37002 43002
rect 37002 42950 37012 43002
rect 37036 42950 37066 43002
rect 37066 42950 37078 43002
rect 37078 42950 37092 43002
rect 37116 42950 37130 43002
rect 37130 42950 37142 43002
rect 37142 42950 37172 43002
rect 37196 42950 37206 43002
rect 37206 42950 37252 43002
rect 36956 42948 37012 42950
rect 37036 42948 37092 42950
rect 37116 42948 37172 42950
rect 37196 42948 37252 42950
rect 36956 41914 37012 41916
rect 37036 41914 37092 41916
rect 37116 41914 37172 41916
rect 37196 41914 37252 41916
rect 36956 41862 37002 41914
rect 37002 41862 37012 41914
rect 37036 41862 37066 41914
rect 37066 41862 37078 41914
rect 37078 41862 37092 41914
rect 37116 41862 37130 41914
rect 37130 41862 37142 41914
rect 37142 41862 37172 41914
rect 37196 41862 37206 41914
rect 37206 41862 37252 41914
rect 36956 41860 37012 41862
rect 37036 41860 37092 41862
rect 37116 41860 37172 41862
rect 37196 41860 37252 41862
rect 36956 40826 37012 40828
rect 37036 40826 37092 40828
rect 37116 40826 37172 40828
rect 37196 40826 37252 40828
rect 36956 40774 37002 40826
rect 37002 40774 37012 40826
rect 37036 40774 37066 40826
rect 37066 40774 37078 40826
rect 37078 40774 37092 40826
rect 37116 40774 37130 40826
rect 37130 40774 37142 40826
rect 37142 40774 37172 40826
rect 37196 40774 37206 40826
rect 37206 40774 37252 40826
rect 36956 40772 37012 40774
rect 37036 40772 37092 40774
rect 37116 40772 37172 40774
rect 37196 40772 37252 40774
rect 36956 39738 37012 39740
rect 37036 39738 37092 39740
rect 37116 39738 37172 39740
rect 37196 39738 37252 39740
rect 36956 39686 37002 39738
rect 37002 39686 37012 39738
rect 37036 39686 37066 39738
rect 37066 39686 37078 39738
rect 37078 39686 37092 39738
rect 37116 39686 37130 39738
rect 37130 39686 37142 39738
rect 37142 39686 37172 39738
rect 37196 39686 37206 39738
rect 37206 39686 37252 39738
rect 36956 39684 37012 39686
rect 37036 39684 37092 39686
rect 37116 39684 37172 39686
rect 37196 39684 37252 39686
rect 36956 38650 37012 38652
rect 37036 38650 37092 38652
rect 37116 38650 37172 38652
rect 37196 38650 37252 38652
rect 36956 38598 37002 38650
rect 37002 38598 37012 38650
rect 37036 38598 37066 38650
rect 37066 38598 37078 38650
rect 37078 38598 37092 38650
rect 37116 38598 37130 38650
rect 37130 38598 37142 38650
rect 37142 38598 37172 38650
rect 37196 38598 37206 38650
rect 37206 38598 37252 38650
rect 36956 38596 37012 38598
rect 37036 38596 37092 38598
rect 37116 38596 37172 38598
rect 37196 38596 37252 38598
rect 36956 37562 37012 37564
rect 37036 37562 37092 37564
rect 37116 37562 37172 37564
rect 37196 37562 37252 37564
rect 36956 37510 37002 37562
rect 37002 37510 37012 37562
rect 37036 37510 37066 37562
rect 37066 37510 37078 37562
rect 37078 37510 37092 37562
rect 37116 37510 37130 37562
rect 37130 37510 37142 37562
rect 37142 37510 37172 37562
rect 37196 37510 37206 37562
rect 37206 37510 37252 37562
rect 36956 37508 37012 37510
rect 37036 37508 37092 37510
rect 37116 37508 37172 37510
rect 37196 37508 37252 37510
rect 36956 36474 37012 36476
rect 37036 36474 37092 36476
rect 37116 36474 37172 36476
rect 37196 36474 37252 36476
rect 36956 36422 37002 36474
rect 37002 36422 37012 36474
rect 37036 36422 37066 36474
rect 37066 36422 37078 36474
rect 37078 36422 37092 36474
rect 37116 36422 37130 36474
rect 37130 36422 37142 36474
rect 37142 36422 37172 36474
rect 37196 36422 37206 36474
rect 37206 36422 37252 36474
rect 36956 36420 37012 36422
rect 37036 36420 37092 36422
rect 37116 36420 37172 36422
rect 37196 36420 37252 36422
rect 36956 35386 37012 35388
rect 37036 35386 37092 35388
rect 37116 35386 37172 35388
rect 37196 35386 37252 35388
rect 36956 35334 37002 35386
rect 37002 35334 37012 35386
rect 37036 35334 37066 35386
rect 37066 35334 37078 35386
rect 37078 35334 37092 35386
rect 37116 35334 37130 35386
rect 37130 35334 37142 35386
rect 37142 35334 37172 35386
rect 37196 35334 37206 35386
rect 37206 35334 37252 35386
rect 36956 35332 37012 35334
rect 37036 35332 37092 35334
rect 37116 35332 37172 35334
rect 37196 35332 37252 35334
rect 36956 34298 37012 34300
rect 37036 34298 37092 34300
rect 37116 34298 37172 34300
rect 37196 34298 37252 34300
rect 36956 34246 37002 34298
rect 37002 34246 37012 34298
rect 37036 34246 37066 34298
rect 37066 34246 37078 34298
rect 37078 34246 37092 34298
rect 37116 34246 37130 34298
rect 37130 34246 37142 34298
rect 37142 34246 37172 34298
rect 37196 34246 37206 34298
rect 37206 34246 37252 34298
rect 36956 34244 37012 34246
rect 37036 34244 37092 34246
rect 37116 34244 37172 34246
rect 37196 34244 37252 34246
rect 36956 33210 37012 33212
rect 37036 33210 37092 33212
rect 37116 33210 37172 33212
rect 37196 33210 37252 33212
rect 36956 33158 37002 33210
rect 37002 33158 37012 33210
rect 37036 33158 37066 33210
rect 37066 33158 37078 33210
rect 37078 33158 37092 33210
rect 37116 33158 37130 33210
rect 37130 33158 37142 33210
rect 37142 33158 37172 33210
rect 37196 33158 37206 33210
rect 37206 33158 37252 33210
rect 36956 33156 37012 33158
rect 37036 33156 37092 33158
rect 37116 33156 37172 33158
rect 37196 33156 37252 33158
rect 36956 32122 37012 32124
rect 37036 32122 37092 32124
rect 37116 32122 37172 32124
rect 37196 32122 37252 32124
rect 36956 32070 37002 32122
rect 37002 32070 37012 32122
rect 37036 32070 37066 32122
rect 37066 32070 37078 32122
rect 37078 32070 37092 32122
rect 37116 32070 37130 32122
rect 37130 32070 37142 32122
rect 37142 32070 37172 32122
rect 37196 32070 37206 32122
rect 37206 32070 37252 32122
rect 36956 32068 37012 32070
rect 37036 32068 37092 32070
rect 37116 32068 37172 32070
rect 37196 32068 37252 32070
rect 36956 31034 37012 31036
rect 37036 31034 37092 31036
rect 37116 31034 37172 31036
rect 37196 31034 37252 31036
rect 36956 30982 37002 31034
rect 37002 30982 37012 31034
rect 37036 30982 37066 31034
rect 37066 30982 37078 31034
rect 37078 30982 37092 31034
rect 37116 30982 37130 31034
rect 37130 30982 37142 31034
rect 37142 30982 37172 31034
rect 37196 30982 37206 31034
rect 37206 30982 37252 31034
rect 36956 30980 37012 30982
rect 37036 30980 37092 30982
rect 37116 30980 37172 30982
rect 37196 30980 37252 30982
rect 36956 29946 37012 29948
rect 37036 29946 37092 29948
rect 37116 29946 37172 29948
rect 37196 29946 37252 29948
rect 36956 29894 37002 29946
rect 37002 29894 37012 29946
rect 37036 29894 37066 29946
rect 37066 29894 37078 29946
rect 37078 29894 37092 29946
rect 37116 29894 37130 29946
rect 37130 29894 37142 29946
rect 37142 29894 37172 29946
rect 37196 29894 37206 29946
rect 37206 29894 37252 29946
rect 36956 29892 37012 29894
rect 37036 29892 37092 29894
rect 37116 29892 37172 29894
rect 37196 29892 37252 29894
rect 36956 28858 37012 28860
rect 37036 28858 37092 28860
rect 37116 28858 37172 28860
rect 37196 28858 37252 28860
rect 36956 28806 37002 28858
rect 37002 28806 37012 28858
rect 37036 28806 37066 28858
rect 37066 28806 37078 28858
rect 37078 28806 37092 28858
rect 37116 28806 37130 28858
rect 37130 28806 37142 28858
rect 37142 28806 37172 28858
rect 37196 28806 37206 28858
rect 37206 28806 37252 28858
rect 36956 28804 37012 28806
rect 37036 28804 37092 28806
rect 37116 28804 37172 28806
rect 37196 28804 37252 28806
rect 36956 27770 37012 27772
rect 37036 27770 37092 27772
rect 37116 27770 37172 27772
rect 37196 27770 37252 27772
rect 36956 27718 37002 27770
rect 37002 27718 37012 27770
rect 37036 27718 37066 27770
rect 37066 27718 37078 27770
rect 37078 27718 37092 27770
rect 37116 27718 37130 27770
rect 37130 27718 37142 27770
rect 37142 27718 37172 27770
rect 37196 27718 37206 27770
rect 37206 27718 37252 27770
rect 36956 27716 37012 27718
rect 37036 27716 37092 27718
rect 37116 27716 37172 27718
rect 37196 27716 37252 27718
rect 36956 26682 37012 26684
rect 37036 26682 37092 26684
rect 37116 26682 37172 26684
rect 37196 26682 37252 26684
rect 36956 26630 37002 26682
rect 37002 26630 37012 26682
rect 37036 26630 37066 26682
rect 37066 26630 37078 26682
rect 37078 26630 37092 26682
rect 37116 26630 37130 26682
rect 37130 26630 37142 26682
rect 37142 26630 37172 26682
rect 37196 26630 37206 26682
rect 37206 26630 37252 26682
rect 36956 26628 37012 26630
rect 37036 26628 37092 26630
rect 37116 26628 37172 26630
rect 37196 26628 37252 26630
rect 36956 25594 37012 25596
rect 37036 25594 37092 25596
rect 37116 25594 37172 25596
rect 37196 25594 37252 25596
rect 36956 25542 37002 25594
rect 37002 25542 37012 25594
rect 37036 25542 37066 25594
rect 37066 25542 37078 25594
rect 37078 25542 37092 25594
rect 37116 25542 37130 25594
rect 37130 25542 37142 25594
rect 37142 25542 37172 25594
rect 37196 25542 37206 25594
rect 37206 25542 37252 25594
rect 36956 25540 37012 25542
rect 37036 25540 37092 25542
rect 37116 25540 37172 25542
rect 37196 25540 37252 25542
rect 36956 24506 37012 24508
rect 37036 24506 37092 24508
rect 37116 24506 37172 24508
rect 37196 24506 37252 24508
rect 36956 24454 37002 24506
rect 37002 24454 37012 24506
rect 37036 24454 37066 24506
rect 37066 24454 37078 24506
rect 37078 24454 37092 24506
rect 37116 24454 37130 24506
rect 37130 24454 37142 24506
rect 37142 24454 37172 24506
rect 37196 24454 37206 24506
rect 37206 24454 37252 24506
rect 36956 24452 37012 24454
rect 37036 24452 37092 24454
rect 37116 24452 37172 24454
rect 37196 24452 37252 24454
rect 36956 23418 37012 23420
rect 37036 23418 37092 23420
rect 37116 23418 37172 23420
rect 37196 23418 37252 23420
rect 36956 23366 37002 23418
rect 37002 23366 37012 23418
rect 37036 23366 37066 23418
rect 37066 23366 37078 23418
rect 37078 23366 37092 23418
rect 37116 23366 37130 23418
rect 37130 23366 37142 23418
rect 37142 23366 37172 23418
rect 37196 23366 37206 23418
rect 37206 23366 37252 23418
rect 36956 23364 37012 23366
rect 37036 23364 37092 23366
rect 37116 23364 37172 23366
rect 37196 23364 37252 23366
rect 36956 22330 37012 22332
rect 37036 22330 37092 22332
rect 37116 22330 37172 22332
rect 37196 22330 37252 22332
rect 36956 22278 37002 22330
rect 37002 22278 37012 22330
rect 37036 22278 37066 22330
rect 37066 22278 37078 22330
rect 37078 22278 37092 22330
rect 37116 22278 37130 22330
rect 37130 22278 37142 22330
rect 37142 22278 37172 22330
rect 37196 22278 37206 22330
rect 37206 22278 37252 22330
rect 36956 22276 37012 22278
rect 37036 22276 37092 22278
rect 37116 22276 37172 22278
rect 37196 22276 37252 22278
rect 36956 21242 37012 21244
rect 37036 21242 37092 21244
rect 37116 21242 37172 21244
rect 37196 21242 37252 21244
rect 36956 21190 37002 21242
rect 37002 21190 37012 21242
rect 37036 21190 37066 21242
rect 37066 21190 37078 21242
rect 37078 21190 37092 21242
rect 37116 21190 37130 21242
rect 37130 21190 37142 21242
rect 37142 21190 37172 21242
rect 37196 21190 37206 21242
rect 37206 21190 37252 21242
rect 36956 21188 37012 21190
rect 37036 21188 37092 21190
rect 37116 21188 37172 21190
rect 37196 21188 37252 21190
rect 36956 20154 37012 20156
rect 37036 20154 37092 20156
rect 37116 20154 37172 20156
rect 37196 20154 37252 20156
rect 36956 20102 37002 20154
rect 37002 20102 37012 20154
rect 37036 20102 37066 20154
rect 37066 20102 37078 20154
rect 37078 20102 37092 20154
rect 37116 20102 37130 20154
rect 37130 20102 37142 20154
rect 37142 20102 37172 20154
rect 37196 20102 37206 20154
rect 37206 20102 37252 20154
rect 36956 20100 37012 20102
rect 37036 20100 37092 20102
rect 37116 20100 37172 20102
rect 37196 20100 37252 20102
rect 36956 19066 37012 19068
rect 37036 19066 37092 19068
rect 37116 19066 37172 19068
rect 37196 19066 37252 19068
rect 36956 19014 37002 19066
rect 37002 19014 37012 19066
rect 37036 19014 37066 19066
rect 37066 19014 37078 19066
rect 37078 19014 37092 19066
rect 37116 19014 37130 19066
rect 37130 19014 37142 19066
rect 37142 19014 37172 19066
rect 37196 19014 37206 19066
rect 37206 19014 37252 19066
rect 36956 19012 37012 19014
rect 37036 19012 37092 19014
rect 37116 19012 37172 19014
rect 37196 19012 37252 19014
rect 36956 17978 37012 17980
rect 37036 17978 37092 17980
rect 37116 17978 37172 17980
rect 37196 17978 37252 17980
rect 36956 17926 37002 17978
rect 37002 17926 37012 17978
rect 37036 17926 37066 17978
rect 37066 17926 37078 17978
rect 37078 17926 37092 17978
rect 37116 17926 37130 17978
rect 37130 17926 37142 17978
rect 37142 17926 37172 17978
rect 37196 17926 37206 17978
rect 37206 17926 37252 17978
rect 36956 17924 37012 17926
rect 37036 17924 37092 17926
rect 37116 17924 37172 17926
rect 37196 17924 37252 17926
rect 36956 16890 37012 16892
rect 37036 16890 37092 16892
rect 37116 16890 37172 16892
rect 37196 16890 37252 16892
rect 36956 16838 37002 16890
rect 37002 16838 37012 16890
rect 37036 16838 37066 16890
rect 37066 16838 37078 16890
rect 37078 16838 37092 16890
rect 37116 16838 37130 16890
rect 37130 16838 37142 16890
rect 37142 16838 37172 16890
rect 37196 16838 37206 16890
rect 37206 16838 37252 16890
rect 36956 16836 37012 16838
rect 37036 16836 37092 16838
rect 37116 16836 37172 16838
rect 37196 16836 37252 16838
rect 36956 15802 37012 15804
rect 37036 15802 37092 15804
rect 37116 15802 37172 15804
rect 37196 15802 37252 15804
rect 36956 15750 37002 15802
rect 37002 15750 37012 15802
rect 37036 15750 37066 15802
rect 37066 15750 37078 15802
rect 37078 15750 37092 15802
rect 37116 15750 37130 15802
rect 37130 15750 37142 15802
rect 37142 15750 37172 15802
rect 37196 15750 37206 15802
rect 37206 15750 37252 15802
rect 36956 15748 37012 15750
rect 37036 15748 37092 15750
rect 37116 15748 37172 15750
rect 37196 15748 37252 15750
rect 36956 14714 37012 14716
rect 37036 14714 37092 14716
rect 37116 14714 37172 14716
rect 37196 14714 37252 14716
rect 36956 14662 37002 14714
rect 37002 14662 37012 14714
rect 37036 14662 37066 14714
rect 37066 14662 37078 14714
rect 37078 14662 37092 14714
rect 37116 14662 37130 14714
rect 37130 14662 37142 14714
rect 37142 14662 37172 14714
rect 37196 14662 37206 14714
rect 37206 14662 37252 14714
rect 36956 14660 37012 14662
rect 37036 14660 37092 14662
rect 37116 14660 37172 14662
rect 37196 14660 37252 14662
rect 36956 13626 37012 13628
rect 37036 13626 37092 13628
rect 37116 13626 37172 13628
rect 37196 13626 37252 13628
rect 36956 13574 37002 13626
rect 37002 13574 37012 13626
rect 37036 13574 37066 13626
rect 37066 13574 37078 13626
rect 37078 13574 37092 13626
rect 37116 13574 37130 13626
rect 37130 13574 37142 13626
rect 37142 13574 37172 13626
rect 37196 13574 37206 13626
rect 37206 13574 37252 13626
rect 36956 13572 37012 13574
rect 37036 13572 37092 13574
rect 37116 13572 37172 13574
rect 37196 13572 37252 13574
rect 36956 12538 37012 12540
rect 37036 12538 37092 12540
rect 37116 12538 37172 12540
rect 37196 12538 37252 12540
rect 36956 12486 37002 12538
rect 37002 12486 37012 12538
rect 37036 12486 37066 12538
rect 37066 12486 37078 12538
rect 37078 12486 37092 12538
rect 37116 12486 37130 12538
rect 37130 12486 37142 12538
rect 37142 12486 37172 12538
rect 37196 12486 37206 12538
rect 37206 12486 37252 12538
rect 36956 12484 37012 12486
rect 37036 12484 37092 12486
rect 37116 12484 37172 12486
rect 37196 12484 37252 12486
rect 36956 11450 37012 11452
rect 37036 11450 37092 11452
rect 37116 11450 37172 11452
rect 37196 11450 37252 11452
rect 36956 11398 37002 11450
rect 37002 11398 37012 11450
rect 37036 11398 37066 11450
rect 37066 11398 37078 11450
rect 37078 11398 37092 11450
rect 37116 11398 37130 11450
rect 37130 11398 37142 11450
rect 37142 11398 37172 11450
rect 37196 11398 37206 11450
rect 37206 11398 37252 11450
rect 36956 11396 37012 11398
rect 37036 11396 37092 11398
rect 37116 11396 37172 11398
rect 37196 11396 37252 11398
rect 36956 10362 37012 10364
rect 37036 10362 37092 10364
rect 37116 10362 37172 10364
rect 37196 10362 37252 10364
rect 36956 10310 37002 10362
rect 37002 10310 37012 10362
rect 37036 10310 37066 10362
rect 37066 10310 37078 10362
rect 37078 10310 37092 10362
rect 37116 10310 37130 10362
rect 37130 10310 37142 10362
rect 37142 10310 37172 10362
rect 37196 10310 37206 10362
rect 37206 10310 37252 10362
rect 36956 10308 37012 10310
rect 37036 10308 37092 10310
rect 37116 10308 37172 10310
rect 37196 10308 37252 10310
rect 36956 9274 37012 9276
rect 37036 9274 37092 9276
rect 37116 9274 37172 9276
rect 37196 9274 37252 9276
rect 36956 9222 37002 9274
rect 37002 9222 37012 9274
rect 37036 9222 37066 9274
rect 37066 9222 37078 9274
rect 37078 9222 37092 9274
rect 37116 9222 37130 9274
rect 37130 9222 37142 9274
rect 37142 9222 37172 9274
rect 37196 9222 37206 9274
rect 37206 9222 37252 9274
rect 36956 9220 37012 9222
rect 37036 9220 37092 9222
rect 37116 9220 37172 9222
rect 37196 9220 37252 9222
rect 36956 8186 37012 8188
rect 37036 8186 37092 8188
rect 37116 8186 37172 8188
rect 37196 8186 37252 8188
rect 36956 8134 37002 8186
rect 37002 8134 37012 8186
rect 37036 8134 37066 8186
rect 37066 8134 37078 8186
rect 37078 8134 37092 8186
rect 37116 8134 37130 8186
rect 37130 8134 37142 8186
rect 37142 8134 37172 8186
rect 37196 8134 37206 8186
rect 37206 8134 37252 8186
rect 36956 8132 37012 8134
rect 37036 8132 37092 8134
rect 37116 8132 37172 8134
rect 37196 8132 37252 8134
rect 36956 7098 37012 7100
rect 37036 7098 37092 7100
rect 37116 7098 37172 7100
rect 37196 7098 37252 7100
rect 36956 7046 37002 7098
rect 37002 7046 37012 7098
rect 37036 7046 37066 7098
rect 37066 7046 37078 7098
rect 37078 7046 37092 7098
rect 37116 7046 37130 7098
rect 37130 7046 37142 7098
rect 37142 7046 37172 7098
rect 37196 7046 37206 7098
rect 37206 7046 37252 7098
rect 36956 7044 37012 7046
rect 37036 7044 37092 7046
rect 37116 7044 37172 7046
rect 37196 7044 37252 7046
rect 37616 54426 37672 54428
rect 37696 54426 37752 54428
rect 37776 54426 37832 54428
rect 37856 54426 37912 54428
rect 37616 54374 37662 54426
rect 37662 54374 37672 54426
rect 37696 54374 37726 54426
rect 37726 54374 37738 54426
rect 37738 54374 37752 54426
rect 37776 54374 37790 54426
rect 37790 54374 37802 54426
rect 37802 54374 37832 54426
rect 37856 54374 37866 54426
rect 37866 54374 37912 54426
rect 37616 54372 37672 54374
rect 37696 54372 37752 54374
rect 37776 54372 37832 54374
rect 37856 54372 37912 54374
rect 37616 53338 37672 53340
rect 37696 53338 37752 53340
rect 37776 53338 37832 53340
rect 37856 53338 37912 53340
rect 37616 53286 37662 53338
rect 37662 53286 37672 53338
rect 37696 53286 37726 53338
rect 37726 53286 37738 53338
rect 37738 53286 37752 53338
rect 37776 53286 37790 53338
rect 37790 53286 37802 53338
rect 37802 53286 37832 53338
rect 37856 53286 37866 53338
rect 37866 53286 37912 53338
rect 37616 53284 37672 53286
rect 37696 53284 37752 53286
rect 37776 53284 37832 53286
rect 37856 53284 37912 53286
rect 37616 52250 37672 52252
rect 37696 52250 37752 52252
rect 37776 52250 37832 52252
rect 37856 52250 37912 52252
rect 37616 52198 37662 52250
rect 37662 52198 37672 52250
rect 37696 52198 37726 52250
rect 37726 52198 37738 52250
rect 37738 52198 37752 52250
rect 37776 52198 37790 52250
rect 37790 52198 37802 52250
rect 37802 52198 37832 52250
rect 37856 52198 37866 52250
rect 37866 52198 37912 52250
rect 37616 52196 37672 52198
rect 37696 52196 37752 52198
rect 37776 52196 37832 52198
rect 37856 52196 37912 52198
rect 37616 51162 37672 51164
rect 37696 51162 37752 51164
rect 37776 51162 37832 51164
rect 37856 51162 37912 51164
rect 37616 51110 37662 51162
rect 37662 51110 37672 51162
rect 37696 51110 37726 51162
rect 37726 51110 37738 51162
rect 37738 51110 37752 51162
rect 37776 51110 37790 51162
rect 37790 51110 37802 51162
rect 37802 51110 37832 51162
rect 37856 51110 37866 51162
rect 37866 51110 37912 51162
rect 37616 51108 37672 51110
rect 37696 51108 37752 51110
rect 37776 51108 37832 51110
rect 37856 51108 37912 51110
rect 37616 50074 37672 50076
rect 37696 50074 37752 50076
rect 37776 50074 37832 50076
rect 37856 50074 37912 50076
rect 37616 50022 37662 50074
rect 37662 50022 37672 50074
rect 37696 50022 37726 50074
rect 37726 50022 37738 50074
rect 37738 50022 37752 50074
rect 37776 50022 37790 50074
rect 37790 50022 37802 50074
rect 37802 50022 37832 50074
rect 37856 50022 37866 50074
rect 37866 50022 37912 50074
rect 37616 50020 37672 50022
rect 37696 50020 37752 50022
rect 37776 50020 37832 50022
rect 37856 50020 37912 50022
rect 37616 48986 37672 48988
rect 37696 48986 37752 48988
rect 37776 48986 37832 48988
rect 37856 48986 37912 48988
rect 37616 48934 37662 48986
rect 37662 48934 37672 48986
rect 37696 48934 37726 48986
rect 37726 48934 37738 48986
rect 37738 48934 37752 48986
rect 37776 48934 37790 48986
rect 37790 48934 37802 48986
rect 37802 48934 37832 48986
rect 37856 48934 37866 48986
rect 37866 48934 37912 48986
rect 37616 48932 37672 48934
rect 37696 48932 37752 48934
rect 37776 48932 37832 48934
rect 37856 48932 37912 48934
rect 37616 47898 37672 47900
rect 37696 47898 37752 47900
rect 37776 47898 37832 47900
rect 37856 47898 37912 47900
rect 37616 47846 37662 47898
rect 37662 47846 37672 47898
rect 37696 47846 37726 47898
rect 37726 47846 37738 47898
rect 37738 47846 37752 47898
rect 37776 47846 37790 47898
rect 37790 47846 37802 47898
rect 37802 47846 37832 47898
rect 37856 47846 37866 47898
rect 37866 47846 37912 47898
rect 37616 47844 37672 47846
rect 37696 47844 37752 47846
rect 37776 47844 37832 47846
rect 37856 47844 37912 47846
rect 37616 46810 37672 46812
rect 37696 46810 37752 46812
rect 37776 46810 37832 46812
rect 37856 46810 37912 46812
rect 37616 46758 37662 46810
rect 37662 46758 37672 46810
rect 37696 46758 37726 46810
rect 37726 46758 37738 46810
rect 37738 46758 37752 46810
rect 37776 46758 37790 46810
rect 37790 46758 37802 46810
rect 37802 46758 37832 46810
rect 37856 46758 37866 46810
rect 37866 46758 37912 46810
rect 37616 46756 37672 46758
rect 37696 46756 37752 46758
rect 37776 46756 37832 46758
rect 37856 46756 37912 46758
rect 37616 45722 37672 45724
rect 37696 45722 37752 45724
rect 37776 45722 37832 45724
rect 37856 45722 37912 45724
rect 37616 45670 37662 45722
rect 37662 45670 37672 45722
rect 37696 45670 37726 45722
rect 37726 45670 37738 45722
rect 37738 45670 37752 45722
rect 37776 45670 37790 45722
rect 37790 45670 37802 45722
rect 37802 45670 37832 45722
rect 37856 45670 37866 45722
rect 37866 45670 37912 45722
rect 37616 45668 37672 45670
rect 37696 45668 37752 45670
rect 37776 45668 37832 45670
rect 37856 45668 37912 45670
rect 37616 44634 37672 44636
rect 37696 44634 37752 44636
rect 37776 44634 37832 44636
rect 37856 44634 37912 44636
rect 37616 44582 37662 44634
rect 37662 44582 37672 44634
rect 37696 44582 37726 44634
rect 37726 44582 37738 44634
rect 37738 44582 37752 44634
rect 37776 44582 37790 44634
rect 37790 44582 37802 44634
rect 37802 44582 37832 44634
rect 37856 44582 37866 44634
rect 37866 44582 37912 44634
rect 37616 44580 37672 44582
rect 37696 44580 37752 44582
rect 37776 44580 37832 44582
rect 37856 44580 37912 44582
rect 37616 43546 37672 43548
rect 37696 43546 37752 43548
rect 37776 43546 37832 43548
rect 37856 43546 37912 43548
rect 37616 43494 37662 43546
rect 37662 43494 37672 43546
rect 37696 43494 37726 43546
rect 37726 43494 37738 43546
rect 37738 43494 37752 43546
rect 37776 43494 37790 43546
rect 37790 43494 37802 43546
rect 37802 43494 37832 43546
rect 37856 43494 37866 43546
rect 37866 43494 37912 43546
rect 37616 43492 37672 43494
rect 37696 43492 37752 43494
rect 37776 43492 37832 43494
rect 37856 43492 37912 43494
rect 37616 42458 37672 42460
rect 37696 42458 37752 42460
rect 37776 42458 37832 42460
rect 37856 42458 37912 42460
rect 37616 42406 37662 42458
rect 37662 42406 37672 42458
rect 37696 42406 37726 42458
rect 37726 42406 37738 42458
rect 37738 42406 37752 42458
rect 37776 42406 37790 42458
rect 37790 42406 37802 42458
rect 37802 42406 37832 42458
rect 37856 42406 37866 42458
rect 37866 42406 37912 42458
rect 37616 42404 37672 42406
rect 37696 42404 37752 42406
rect 37776 42404 37832 42406
rect 37856 42404 37912 42406
rect 37616 41370 37672 41372
rect 37696 41370 37752 41372
rect 37776 41370 37832 41372
rect 37856 41370 37912 41372
rect 37616 41318 37662 41370
rect 37662 41318 37672 41370
rect 37696 41318 37726 41370
rect 37726 41318 37738 41370
rect 37738 41318 37752 41370
rect 37776 41318 37790 41370
rect 37790 41318 37802 41370
rect 37802 41318 37832 41370
rect 37856 41318 37866 41370
rect 37866 41318 37912 41370
rect 37616 41316 37672 41318
rect 37696 41316 37752 41318
rect 37776 41316 37832 41318
rect 37856 41316 37912 41318
rect 37616 40282 37672 40284
rect 37696 40282 37752 40284
rect 37776 40282 37832 40284
rect 37856 40282 37912 40284
rect 37616 40230 37662 40282
rect 37662 40230 37672 40282
rect 37696 40230 37726 40282
rect 37726 40230 37738 40282
rect 37738 40230 37752 40282
rect 37776 40230 37790 40282
rect 37790 40230 37802 40282
rect 37802 40230 37832 40282
rect 37856 40230 37866 40282
rect 37866 40230 37912 40282
rect 37616 40228 37672 40230
rect 37696 40228 37752 40230
rect 37776 40228 37832 40230
rect 37856 40228 37912 40230
rect 37616 39194 37672 39196
rect 37696 39194 37752 39196
rect 37776 39194 37832 39196
rect 37856 39194 37912 39196
rect 37616 39142 37662 39194
rect 37662 39142 37672 39194
rect 37696 39142 37726 39194
rect 37726 39142 37738 39194
rect 37738 39142 37752 39194
rect 37776 39142 37790 39194
rect 37790 39142 37802 39194
rect 37802 39142 37832 39194
rect 37856 39142 37866 39194
rect 37866 39142 37912 39194
rect 37616 39140 37672 39142
rect 37696 39140 37752 39142
rect 37776 39140 37832 39142
rect 37856 39140 37912 39142
rect 37616 38106 37672 38108
rect 37696 38106 37752 38108
rect 37776 38106 37832 38108
rect 37856 38106 37912 38108
rect 37616 38054 37662 38106
rect 37662 38054 37672 38106
rect 37696 38054 37726 38106
rect 37726 38054 37738 38106
rect 37738 38054 37752 38106
rect 37776 38054 37790 38106
rect 37790 38054 37802 38106
rect 37802 38054 37832 38106
rect 37856 38054 37866 38106
rect 37866 38054 37912 38106
rect 37616 38052 37672 38054
rect 37696 38052 37752 38054
rect 37776 38052 37832 38054
rect 37856 38052 37912 38054
rect 37616 37018 37672 37020
rect 37696 37018 37752 37020
rect 37776 37018 37832 37020
rect 37856 37018 37912 37020
rect 37616 36966 37662 37018
rect 37662 36966 37672 37018
rect 37696 36966 37726 37018
rect 37726 36966 37738 37018
rect 37738 36966 37752 37018
rect 37776 36966 37790 37018
rect 37790 36966 37802 37018
rect 37802 36966 37832 37018
rect 37856 36966 37866 37018
rect 37866 36966 37912 37018
rect 37616 36964 37672 36966
rect 37696 36964 37752 36966
rect 37776 36964 37832 36966
rect 37856 36964 37912 36966
rect 40498 67244 40554 67280
rect 40498 67224 40500 67244
rect 40500 67224 40552 67244
rect 40552 67224 40554 67244
rect 37616 35930 37672 35932
rect 37696 35930 37752 35932
rect 37776 35930 37832 35932
rect 37856 35930 37912 35932
rect 37616 35878 37662 35930
rect 37662 35878 37672 35930
rect 37696 35878 37726 35930
rect 37726 35878 37738 35930
rect 37738 35878 37752 35930
rect 37776 35878 37790 35930
rect 37790 35878 37802 35930
rect 37802 35878 37832 35930
rect 37856 35878 37866 35930
rect 37866 35878 37912 35930
rect 37616 35876 37672 35878
rect 37696 35876 37752 35878
rect 37776 35876 37832 35878
rect 37856 35876 37912 35878
rect 37616 34842 37672 34844
rect 37696 34842 37752 34844
rect 37776 34842 37832 34844
rect 37856 34842 37912 34844
rect 37616 34790 37662 34842
rect 37662 34790 37672 34842
rect 37696 34790 37726 34842
rect 37726 34790 37738 34842
rect 37738 34790 37752 34842
rect 37776 34790 37790 34842
rect 37790 34790 37802 34842
rect 37802 34790 37832 34842
rect 37856 34790 37866 34842
rect 37866 34790 37912 34842
rect 37616 34788 37672 34790
rect 37696 34788 37752 34790
rect 37776 34788 37832 34790
rect 37856 34788 37912 34790
rect 37616 33754 37672 33756
rect 37696 33754 37752 33756
rect 37776 33754 37832 33756
rect 37856 33754 37912 33756
rect 37616 33702 37662 33754
rect 37662 33702 37672 33754
rect 37696 33702 37726 33754
rect 37726 33702 37738 33754
rect 37738 33702 37752 33754
rect 37776 33702 37790 33754
rect 37790 33702 37802 33754
rect 37802 33702 37832 33754
rect 37856 33702 37866 33754
rect 37866 33702 37912 33754
rect 37616 33700 37672 33702
rect 37696 33700 37752 33702
rect 37776 33700 37832 33702
rect 37856 33700 37912 33702
rect 37616 32666 37672 32668
rect 37696 32666 37752 32668
rect 37776 32666 37832 32668
rect 37856 32666 37912 32668
rect 37616 32614 37662 32666
rect 37662 32614 37672 32666
rect 37696 32614 37726 32666
rect 37726 32614 37738 32666
rect 37738 32614 37752 32666
rect 37776 32614 37790 32666
rect 37790 32614 37802 32666
rect 37802 32614 37832 32666
rect 37856 32614 37866 32666
rect 37866 32614 37912 32666
rect 37616 32612 37672 32614
rect 37696 32612 37752 32614
rect 37776 32612 37832 32614
rect 37856 32612 37912 32614
rect 37616 31578 37672 31580
rect 37696 31578 37752 31580
rect 37776 31578 37832 31580
rect 37856 31578 37912 31580
rect 37616 31526 37662 31578
rect 37662 31526 37672 31578
rect 37696 31526 37726 31578
rect 37726 31526 37738 31578
rect 37738 31526 37752 31578
rect 37776 31526 37790 31578
rect 37790 31526 37802 31578
rect 37802 31526 37832 31578
rect 37856 31526 37866 31578
rect 37866 31526 37912 31578
rect 37616 31524 37672 31526
rect 37696 31524 37752 31526
rect 37776 31524 37832 31526
rect 37856 31524 37912 31526
rect 37616 30490 37672 30492
rect 37696 30490 37752 30492
rect 37776 30490 37832 30492
rect 37856 30490 37912 30492
rect 37616 30438 37662 30490
rect 37662 30438 37672 30490
rect 37696 30438 37726 30490
rect 37726 30438 37738 30490
rect 37738 30438 37752 30490
rect 37776 30438 37790 30490
rect 37790 30438 37802 30490
rect 37802 30438 37832 30490
rect 37856 30438 37866 30490
rect 37866 30438 37912 30490
rect 37616 30436 37672 30438
rect 37696 30436 37752 30438
rect 37776 30436 37832 30438
rect 37856 30436 37912 30438
rect 37616 29402 37672 29404
rect 37696 29402 37752 29404
rect 37776 29402 37832 29404
rect 37856 29402 37912 29404
rect 37616 29350 37662 29402
rect 37662 29350 37672 29402
rect 37696 29350 37726 29402
rect 37726 29350 37738 29402
rect 37738 29350 37752 29402
rect 37776 29350 37790 29402
rect 37790 29350 37802 29402
rect 37802 29350 37832 29402
rect 37856 29350 37866 29402
rect 37866 29350 37912 29402
rect 37616 29348 37672 29350
rect 37696 29348 37752 29350
rect 37776 29348 37832 29350
rect 37856 29348 37912 29350
rect 37616 28314 37672 28316
rect 37696 28314 37752 28316
rect 37776 28314 37832 28316
rect 37856 28314 37912 28316
rect 37616 28262 37662 28314
rect 37662 28262 37672 28314
rect 37696 28262 37726 28314
rect 37726 28262 37738 28314
rect 37738 28262 37752 28314
rect 37776 28262 37790 28314
rect 37790 28262 37802 28314
rect 37802 28262 37832 28314
rect 37856 28262 37866 28314
rect 37866 28262 37912 28314
rect 37616 28260 37672 28262
rect 37696 28260 37752 28262
rect 37776 28260 37832 28262
rect 37856 28260 37912 28262
rect 37616 27226 37672 27228
rect 37696 27226 37752 27228
rect 37776 27226 37832 27228
rect 37856 27226 37912 27228
rect 37616 27174 37662 27226
rect 37662 27174 37672 27226
rect 37696 27174 37726 27226
rect 37726 27174 37738 27226
rect 37738 27174 37752 27226
rect 37776 27174 37790 27226
rect 37790 27174 37802 27226
rect 37802 27174 37832 27226
rect 37856 27174 37866 27226
rect 37866 27174 37912 27226
rect 37616 27172 37672 27174
rect 37696 27172 37752 27174
rect 37776 27172 37832 27174
rect 37856 27172 37912 27174
rect 37616 26138 37672 26140
rect 37696 26138 37752 26140
rect 37776 26138 37832 26140
rect 37856 26138 37912 26140
rect 37616 26086 37662 26138
rect 37662 26086 37672 26138
rect 37696 26086 37726 26138
rect 37726 26086 37738 26138
rect 37738 26086 37752 26138
rect 37776 26086 37790 26138
rect 37790 26086 37802 26138
rect 37802 26086 37832 26138
rect 37856 26086 37866 26138
rect 37866 26086 37912 26138
rect 37616 26084 37672 26086
rect 37696 26084 37752 26086
rect 37776 26084 37832 26086
rect 37856 26084 37912 26086
rect 37616 25050 37672 25052
rect 37696 25050 37752 25052
rect 37776 25050 37832 25052
rect 37856 25050 37912 25052
rect 37616 24998 37662 25050
rect 37662 24998 37672 25050
rect 37696 24998 37726 25050
rect 37726 24998 37738 25050
rect 37738 24998 37752 25050
rect 37776 24998 37790 25050
rect 37790 24998 37802 25050
rect 37802 24998 37832 25050
rect 37856 24998 37866 25050
rect 37866 24998 37912 25050
rect 37616 24996 37672 24998
rect 37696 24996 37752 24998
rect 37776 24996 37832 24998
rect 37856 24996 37912 24998
rect 37616 23962 37672 23964
rect 37696 23962 37752 23964
rect 37776 23962 37832 23964
rect 37856 23962 37912 23964
rect 37616 23910 37662 23962
rect 37662 23910 37672 23962
rect 37696 23910 37726 23962
rect 37726 23910 37738 23962
rect 37738 23910 37752 23962
rect 37776 23910 37790 23962
rect 37790 23910 37802 23962
rect 37802 23910 37832 23962
rect 37856 23910 37866 23962
rect 37866 23910 37912 23962
rect 37616 23908 37672 23910
rect 37696 23908 37752 23910
rect 37776 23908 37832 23910
rect 37856 23908 37912 23910
rect 37616 22874 37672 22876
rect 37696 22874 37752 22876
rect 37776 22874 37832 22876
rect 37856 22874 37912 22876
rect 37616 22822 37662 22874
rect 37662 22822 37672 22874
rect 37696 22822 37726 22874
rect 37726 22822 37738 22874
rect 37738 22822 37752 22874
rect 37776 22822 37790 22874
rect 37790 22822 37802 22874
rect 37802 22822 37832 22874
rect 37856 22822 37866 22874
rect 37866 22822 37912 22874
rect 37616 22820 37672 22822
rect 37696 22820 37752 22822
rect 37776 22820 37832 22822
rect 37856 22820 37912 22822
rect 37616 21786 37672 21788
rect 37696 21786 37752 21788
rect 37776 21786 37832 21788
rect 37856 21786 37912 21788
rect 37616 21734 37662 21786
rect 37662 21734 37672 21786
rect 37696 21734 37726 21786
rect 37726 21734 37738 21786
rect 37738 21734 37752 21786
rect 37776 21734 37790 21786
rect 37790 21734 37802 21786
rect 37802 21734 37832 21786
rect 37856 21734 37866 21786
rect 37866 21734 37912 21786
rect 37616 21732 37672 21734
rect 37696 21732 37752 21734
rect 37776 21732 37832 21734
rect 37856 21732 37912 21734
rect 37616 20698 37672 20700
rect 37696 20698 37752 20700
rect 37776 20698 37832 20700
rect 37856 20698 37912 20700
rect 37616 20646 37662 20698
rect 37662 20646 37672 20698
rect 37696 20646 37726 20698
rect 37726 20646 37738 20698
rect 37738 20646 37752 20698
rect 37776 20646 37790 20698
rect 37790 20646 37802 20698
rect 37802 20646 37832 20698
rect 37856 20646 37866 20698
rect 37866 20646 37912 20698
rect 37616 20644 37672 20646
rect 37696 20644 37752 20646
rect 37776 20644 37832 20646
rect 37856 20644 37912 20646
rect 37616 19610 37672 19612
rect 37696 19610 37752 19612
rect 37776 19610 37832 19612
rect 37856 19610 37912 19612
rect 37616 19558 37662 19610
rect 37662 19558 37672 19610
rect 37696 19558 37726 19610
rect 37726 19558 37738 19610
rect 37738 19558 37752 19610
rect 37776 19558 37790 19610
rect 37790 19558 37802 19610
rect 37802 19558 37832 19610
rect 37856 19558 37866 19610
rect 37866 19558 37912 19610
rect 37616 19556 37672 19558
rect 37696 19556 37752 19558
rect 37776 19556 37832 19558
rect 37856 19556 37912 19558
rect 37616 18522 37672 18524
rect 37696 18522 37752 18524
rect 37776 18522 37832 18524
rect 37856 18522 37912 18524
rect 37616 18470 37662 18522
rect 37662 18470 37672 18522
rect 37696 18470 37726 18522
rect 37726 18470 37738 18522
rect 37738 18470 37752 18522
rect 37776 18470 37790 18522
rect 37790 18470 37802 18522
rect 37802 18470 37832 18522
rect 37856 18470 37866 18522
rect 37866 18470 37912 18522
rect 37616 18468 37672 18470
rect 37696 18468 37752 18470
rect 37776 18468 37832 18470
rect 37856 18468 37912 18470
rect 37616 17434 37672 17436
rect 37696 17434 37752 17436
rect 37776 17434 37832 17436
rect 37856 17434 37912 17436
rect 37616 17382 37662 17434
rect 37662 17382 37672 17434
rect 37696 17382 37726 17434
rect 37726 17382 37738 17434
rect 37738 17382 37752 17434
rect 37776 17382 37790 17434
rect 37790 17382 37802 17434
rect 37802 17382 37832 17434
rect 37856 17382 37866 17434
rect 37866 17382 37912 17434
rect 37616 17380 37672 17382
rect 37696 17380 37752 17382
rect 37776 17380 37832 17382
rect 37856 17380 37912 17382
rect 37616 16346 37672 16348
rect 37696 16346 37752 16348
rect 37776 16346 37832 16348
rect 37856 16346 37912 16348
rect 37616 16294 37662 16346
rect 37662 16294 37672 16346
rect 37696 16294 37726 16346
rect 37726 16294 37738 16346
rect 37738 16294 37752 16346
rect 37776 16294 37790 16346
rect 37790 16294 37802 16346
rect 37802 16294 37832 16346
rect 37856 16294 37866 16346
rect 37866 16294 37912 16346
rect 37616 16292 37672 16294
rect 37696 16292 37752 16294
rect 37776 16292 37832 16294
rect 37856 16292 37912 16294
rect 37616 15258 37672 15260
rect 37696 15258 37752 15260
rect 37776 15258 37832 15260
rect 37856 15258 37912 15260
rect 37616 15206 37662 15258
rect 37662 15206 37672 15258
rect 37696 15206 37726 15258
rect 37726 15206 37738 15258
rect 37738 15206 37752 15258
rect 37776 15206 37790 15258
rect 37790 15206 37802 15258
rect 37802 15206 37832 15258
rect 37856 15206 37866 15258
rect 37866 15206 37912 15258
rect 37616 15204 37672 15206
rect 37696 15204 37752 15206
rect 37776 15204 37832 15206
rect 37856 15204 37912 15206
rect 37616 14170 37672 14172
rect 37696 14170 37752 14172
rect 37776 14170 37832 14172
rect 37856 14170 37912 14172
rect 37616 14118 37662 14170
rect 37662 14118 37672 14170
rect 37696 14118 37726 14170
rect 37726 14118 37738 14170
rect 37738 14118 37752 14170
rect 37776 14118 37790 14170
rect 37790 14118 37802 14170
rect 37802 14118 37832 14170
rect 37856 14118 37866 14170
rect 37866 14118 37912 14170
rect 37616 14116 37672 14118
rect 37696 14116 37752 14118
rect 37776 14116 37832 14118
rect 37856 14116 37912 14118
rect 37616 13082 37672 13084
rect 37696 13082 37752 13084
rect 37776 13082 37832 13084
rect 37856 13082 37912 13084
rect 37616 13030 37662 13082
rect 37662 13030 37672 13082
rect 37696 13030 37726 13082
rect 37726 13030 37738 13082
rect 37738 13030 37752 13082
rect 37776 13030 37790 13082
rect 37790 13030 37802 13082
rect 37802 13030 37832 13082
rect 37856 13030 37866 13082
rect 37866 13030 37912 13082
rect 37616 13028 37672 13030
rect 37696 13028 37752 13030
rect 37776 13028 37832 13030
rect 37856 13028 37912 13030
rect 37616 11994 37672 11996
rect 37696 11994 37752 11996
rect 37776 11994 37832 11996
rect 37856 11994 37912 11996
rect 37616 11942 37662 11994
rect 37662 11942 37672 11994
rect 37696 11942 37726 11994
rect 37726 11942 37738 11994
rect 37738 11942 37752 11994
rect 37776 11942 37790 11994
rect 37790 11942 37802 11994
rect 37802 11942 37832 11994
rect 37856 11942 37866 11994
rect 37866 11942 37912 11994
rect 37616 11940 37672 11942
rect 37696 11940 37752 11942
rect 37776 11940 37832 11942
rect 37856 11940 37912 11942
rect 37616 10906 37672 10908
rect 37696 10906 37752 10908
rect 37776 10906 37832 10908
rect 37856 10906 37912 10908
rect 37616 10854 37662 10906
rect 37662 10854 37672 10906
rect 37696 10854 37726 10906
rect 37726 10854 37738 10906
rect 37738 10854 37752 10906
rect 37776 10854 37790 10906
rect 37790 10854 37802 10906
rect 37802 10854 37832 10906
rect 37856 10854 37866 10906
rect 37866 10854 37912 10906
rect 37616 10852 37672 10854
rect 37696 10852 37752 10854
rect 37776 10852 37832 10854
rect 37856 10852 37912 10854
rect 37616 9818 37672 9820
rect 37696 9818 37752 9820
rect 37776 9818 37832 9820
rect 37856 9818 37912 9820
rect 37616 9766 37662 9818
rect 37662 9766 37672 9818
rect 37696 9766 37726 9818
rect 37726 9766 37738 9818
rect 37738 9766 37752 9818
rect 37776 9766 37790 9818
rect 37790 9766 37802 9818
rect 37802 9766 37832 9818
rect 37856 9766 37866 9818
rect 37866 9766 37912 9818
rect 37616 9764 37672 9766
rect 37696 9764 37752 9766
rect 37776 9764 37832 9766
rect 37856 9764 37912 9766
rect 37616 8730 37672 8732
rect 37696 8730 37752 8732
rect 37776 8730 37832 8732
rect 37856 8730 37912 8732
rect 37616 8678 37662 8730
rect 37662 8678 37672 8730
rect 37696 8678 37726 8730
rect 37726 8678 37738 8730
rect 37738 8678 37752 8730
rect 37776 8678 37790 8730
rect 37790 8678 37802 8730
rect 37802 8678 37832 8730
rect 37856 8678 37866 8730
rect 37866 8678 37912 8730
rect 37616 8676 37672 8678
rect 37696 8676 37752 8678
rect 37776 8676 37832 8678
rect 37856 8676 37912 8678
rect 37616 7642 37672 7644
rect 37696 7642 37752 7644
rect 37776 7642 37832 7644
rect 37856 7642 37912 7644
rect 37616 7590 37662 7642
rect 37662 7590 37672 7642
rect 37696 7590 37726 7642
rect 37726 7590 37738 7642
rect 37738 7590 37752 7642
rect 37776 7590 37790 7642
rect 37790 7590 37802 7642
rect 37802 7590 37832 7642
rect 37856 7590 37866 7642
rect 37866 7590 37912 7642
rect 37616 7588 37672 7590
rect 37696 7588 37752 7590
rect 37776 7588 37832 7590
rect 37856 7588 37912 7590
rect 36956 6010 37012 6012
rect 37036 6010 37092 6012
rect 37116 6010 37172 6012
rect 37196 6010 37252 6012
rect 36956 5958 37002 6010
rect 37002 5958 37012 6010
rect 37036 5958 37066 6010
rect 37066 5958 37078 6010
rect 37078 5958 37092 6010
rect 37116 5958 37130 6010
rect 37130 5958 37142 6010
rect 37142 5958 37172 6010
rect 37196 5958 37206 6010
rect 37206 5958 37252 6010
rect 36956 5956 37012 5958
rect 37036 5956 37092 5958
rect 37116 5956 37172 5958
rect 37196 5956 37252 5958
rect 36956 4922 37012 4924
rect 37036 4922 37092 4924
rect 37116 4922 37172 4924
rect 37196 4922 37252 4924
rect 36956 4870 37002 4922
rect 37002 4870 37012 4922
rect 37036 4870 37066 4922
rect 37066 4870 37078 4922
rect 37078 4870 37092 4922
rect 37116 4870 37130 4922
rect 37130 4870 37142 4922
rect 37142 4870 37172 4922
rect 37196 4870 37206 4922
rect 37206 4870 37252 4922
rect 36956 4868 37012 4870
rect 37036 4868 37092 4870
rect 37116 4868 37172 4870
rect 37196 4868 37252 4870
rect 37616 6554 37672 6556
rect 37696 6554 37752 6556
rect 37776 6554 37832 6556
rect 37856 6554 37912 6556
rect 37616 6502 37662 6554
rect 37662 6502 37672 6554
rect 37696 6502 37726 6554
rect 37726 6502 37738 6554
rect 37738 6502 37752 6554
rect 37776 6502 37790 6554
rect 37790 6502 37802 6554
rect 37802 6502 37832 6554
rect 37856 6502 37866 6554
rect 37866 6502 37912 6554
rect 37616 6500 37672 6502
rect 37696 6500 37752 6502
rect 37776 6500 37832 6502
rect 37856 6500 37912 6502
rect 37616 5466 37672 5468
rect 37696 5466 37752 5468
rect 37776 5466 37832 5468
rect 37856 5466 37912 5468
rect 37616 5414 37662 5466
rect 37662 5414 37672 5466
rect 37696 5414 37726 5466
rect 37726 5414 37738 5466
rect 37738 5414 37752 5466
rect 37776 5414 37790 5466
rect 37790 5414 37802 5466
rect 37802 5414 37832 5466
rect 37856 5414 37866 5466
rect 37866 5414 37912 5466
rect 37616 5412 37672 5414
rect 37696 5412 37752 5414
rect 37776 5412 37832 5414
rect 37856 5412 37912 5414
rect 39946 58248 40002 58304
rect 40498 49272 40554 49328
rect 40866 40296 40922 40352
rect 40498 31340 40554 31376
rect 40498 31320 40500 31340
rect 40500 31320 40552 31340
rect 40552 31320 40554 31340
rect 40498 22344 40554 22400
rect 39946 13368 40002 13424
rect 40498 4392 40554 4448
rect 37616 4378 37672 4380
rect 37696 4378 37752 4380
rect 37776 4378 37832 4380
rect 37856 4378 37912 4380
rect 37616 4326 37662 4378
rect 37662 4326 37672 4378
rect 37696 4326 37726 4378
rect 37726 4326 37738 4378
rect 37738 4326 37752 4378
rect 37776 4326 37790 4378
rect 37790 4326 37802 4378
rect 37802 4326 37832 4378
rect 37856 4326 37866 4378
rect 37866 4326 37912 4378
rect 37616 4324 37672 4326
rect 37696 4324 37752 4326
rect 37776 4324 37832 4326
rect 37856 4324 37912 4326
rect 36956 3834 37012 3836
rect 37036 3834 37092 3836
rect 37116 3834 37172 3836
rect 37196 3834 37252 3836
rect 36956 3782 37002 3834
rect 37002 3782 37012 3834
rect 37036 3782 37066 3834
rect 37066 3782 37078 3834
rect 37078 3782 37092 3834
rect 37116 3782 37130 3834
rect 37130 3782 37142 3834
rect 37142 3782 37172 3834
rect 37196 3782 37206 3834
rect 37206 3782 37252 3834
rect 36956 3780 37012 3782
rect 37036 3780 37092 3782
rect 37116 3780 37172 3782
rect 37196 3780 37252 3782
rect 37616 3290 37672 3292
rect 37696 3290 37752 3292
rect 37776 3290 37832 3292
rect 37856 3290 37912 3292
rect 37616 3238 37662 3290
rect 37662 3238 37672 3290
rect 37696 3238 37726 3290
rect 37726 3238 37738 3290
rect 37738 3238 37752 3290
rect 37776 3238 37790 3290
rect 37790 3238 37802 3290
rect 37802 3238 37832 3290
rect 37856 3238 37866 3290
rect 37866 3238 37912 3290
rect 37616 3236 37672 3238
rect 37696 3236 37752 3238
rect 37776 3236 37832 3238
rect 37856 3236 37912 3238
rect 36956 2746 37012 2748
rect 37036 2746 37092 2748
rect 37116 2746 37172 2748
rect 37196 2746 37252 2748
rect 36956 2694 37002 2746
rect 37002 2694 37012 2746
rect 37036 2694 37066 2746
rect 37066 2694 37078 2746
rect 37078 2694 37092 2746
rect 37116 2694 37130 2746
rect 37130 2694 37142 2746
rect 37142 2694 37172 2746
rect 37196 2694 37206 2746
rect 37206 2694 37252 2746
rect 36956 2692 37012 2694
rect 37036 2692 37092 2694
rect 37116 2692 37172 2694
rect 37196 2692 37252 2694
rect 28630 2372 28686 2408
rect 28630 2352 28632 2372
rect 28632 2352 28684 2372
rect 28684 2352 28686 2372
rect 2616 2202 2672 2204
rect 2696 2202 2752 2204
rect 2776 2202 2832 2204
rect 2856 2202 2912 2204
rect 2616 2150 2662 2202
rect 2662 2150 2672 2202
rect 2696 2150 2726 2202
rect 2726 2150 2738 2202
rect 2738 2150 2752 2202
rect 2776 2150 2790 2202
rect 2790 2150 2802 2202
rect 2802 2150 2832 2202
rect 2856 2150 2866 2202
rect 2866 2150 2912 2202
rect 2616 2148 2672 2150
rect 2696 2148 2752 2150
rect 2776 2148 2832 2150
rect 2856 2148 2912 2150
rect 7616 2202 7672 2204
rect 7696 2202 7752 2204
rect 7776 2202 7832 2204
rect 7856 2202 7912 2204
rect 7616 2150 7662 2202
rect 7662 2150 7672 2202
rect 7696 2150 7726 2202
rect 7726 2150 7738 2202
rect 7738 2150 7752 2202
rect 7776 2150 7790 2202
rect 7790 2150 7802 2202
rect 7802 2150 7832 2202
rect 7856 2150 7866 2202
rect 7866 2150 7912 2202
rect 7616 2148 7672 2150
rect 7696 2148 7752 2150
rect 7776 2148 7832 2150
rect 7856 2148 7912 2150
rect 12616 2202 12672 2204
rect 12696 2202 12752 2204
rect 12776 2202 12832 2204
rect 12856 2202 12912 2204
rect 12616 2150 12662 2202
rect 12662 2150 12672 2202
rect 12696 2150 12726 2202
rect 12726 2150 12738 2202
rect 12738 2150 12752 2202
rect 12776 2150 12790 2202
rect 12790 2150 12802 2202
rect 12802 2150 12832 2202
rect 12856 2150 12866 2202
rect 12866 2150 12912 2202
rect 12616 2148 12672 2150
rect 12696 2148 12752 2150
rect 12776 2148 12832 2150
rect 12856 2148 12912 2150
rect 17616 2202 17672 2204
rect 17696 2202 17752 2204
rect 17776 2202 17832 2204
rect 17856 2202 17912 2204
rect 17616 2150 17662 2202
rect 17662 2150 17672 2202
rect 17696 2150 17726 2202
rect 17726 2150 17738 2202
rect 17738 2150 17752 2202
rect 17776 2150 17790 2202
rect 17790 2150 17802 2202
rect 17802 2150 17832 2202
rect 17856 2150 17866 2202
rect 17866 2150 17912 2202
rect 17616 2148 17672 2150
rect 17696 2148 17752 2150
rect 17776 2148 17832 2150
rect 17856 2148 17912 2150
rect 22616 2202 22672 2204
rect 22696 2202 22752 2204
rect 22776 2202 22832 2204
rect 22856 2202 22912 2204
rect 22616 2150 22662 2202
rect 22662 2150 22672 2202
rect 22696 2150 22726 2202
rect 22726 2150 22738 2202
rect 22738 2150 22752 2202
rect 22776 2150 22790 2202
rect 22790 2150 22802 2202
rect 22802 2150 22832 2202
rect 22856 2150 22866 2202
rect 22866 2150 22912 2202
rect 22616 2148 22672 2150
rect 22696 2148 22752 2150
rect 22776 2148 22832 2150
rect 22856 2148 22912 2150
rect 27616 2202 27672 2204
rect 27696 2202 27752 2204
rect 27776 2202 27832 2204
rect 27856 2202 27912 2204
rect 27616 2150 27662 2202
rect 27662 2150 27672 2202
rect 27696 2150 27726 2202
rect 27726 2150 27738 2202
rect 27738 2150 27752 2202
rect 27776 2150 27790 2202
rect 27790 2150 27802 2202
rect 27802 2150 27832 2202
rect 27856 2150 27866 2202
rect 27866 2150 27912 2202
rect 27616 2148 27672 2150
rect 27696 2148 27752 2150
rect 27776 2148 27832 2150
rect 27856 2148 27912 2150
rect 32616 2202 32672 2204
rect 32696 2202 32752 2204
rect 32776 2202 32832 2204
rect 32856 2202 32912 2204
rect 32616 2150 32662 2202
rect 32662 2150 32672 2202
rect 32696 2150 32726 2202
rect 32726 2150 32738 2202
rect 32738 2150 32752 2202
rect 32776 2150 32790 2202
rect 32790 2150 32802 2202
rect 32802 2150 32832 2202
rect 32856 2150 32866 2202
rect 32866 2150 32912 2202
rect 32616 2148 32672 2150
rect 32696 2148 32752 2150
rect 32776 2148 32832 2150
rect 32856 2148 32912 2150
rect 37616 2202 37672 2204
rect 37696 2202 37752 2204
rect 37776 2202 37832 2204
rect 37856 2202 37912 2204
rect 37616 2150 37662 2202
rect 37662 2150 37672 2202
rect 37696 2150 37726 2202
rect 37726 2150 37738 2202
rect 37738 2150 37752 2202
rect 37776 2150 37790 2202
rect 37790 2150 37802 2202
rect 37802 2150 37832 2202
rect 37856 2150 37866 2202
rect 37866 2150 37912 2202
rect 37616 2148 37672 2150
rect 37696 2148 37752 2150
rect 37776 2148 37832 2150
rect 37856 2148 37912 2150
<< metal3 >>
rect 2606 69664 2922 69665
rect 2606 69600 2612 69664
rect 2676 69600 2692 69664
rect 2756 69600 2772 69664
rect 2836 69600 2852 69664
rect 2916 69600 2922 69664
rect 2606 69599 2922 69600
rect 7606 69664 7922 69665
rect 7606 69600 7612 69664
rect 7676 69600 7692 69664
rect 7756 69600 7772 69664
rect 7836 69600 7852 69664
rect 7916 69600 7922 69664
rect 7606 69599 7922 69600
rect 12606 69664 12922 69665
rect 12606 69600 12612 69664
rect 12676 69600 12692 69664
rect 12756 69600 12772 69664
rect 12836 69600 12852 69664
rect 12916 69600 12922 69664
rect 12606 69599 12922 69600
rect 17606 69664 17922 69665
rect 17606 69600 17612 69664
rect 17676 69600 17692 69664
rect 17756 69600 17772 69664
rect 17836 69600 17852 69664
rect 17916 69600 17922 69664
rect 17606 69599 17922 69600
rect 22606 69664 22922 69665
rect 22606 69600 22612 69664
rect 22676 69600 22692 69664
rect 22756 69600 22772 69664
rect 22836 69600 22852 69664
rect 22916 69600 22922 69664
rect 22606 69599 22922 69600
rect 27606 69664 27922 69665
rect 27606 69600 27612 69664
rect 27676 69600 27692 69664
rect 27756 69600 27772 69664
rect 27836 69600 27852 69664
rect 27916 69600 27922 69664
rect 27606 69599 27922 69600
rect 32606 69664 32922 69665
rect 32606 69600 32612 69664
rect 32676 69600 32692 69664
rect 32756 69600 32772 69664
rect 32836 69600 32852 69664
rect 32916 69600 32922 69664
rect 32606 69599 32922 69600
rect 37606 69664 37922 69665
rect 37606 69600 37612 69664
rect 37676 69600 37692 69664
rect 37756 69600 37772 69664
rect 37836 69600 37852 69664
rect 37916 69600 37922 69664
rect 37606 69599 37922 69600
rect 1946 69120 2262 69121
rect 1946 69056 1952 69120
rect 2016 69056 2032 69120
rect 2096 69056 2112 69120
rect 2176 69056 2192 69120
rect 2256 69056 2262 69120
rect 1946 69055 2262 69056
rect 6946 69120 7262 69121
rect 6946 69056 6952 69120
rect 7016 69056 7032 69120
rect 7096 69056 7112 69120
rect 7176 69056 7192 69120
rect 7256 69056 7262 69120
rect 6946 69055 7262 69056
rect 11946 69120 12262 69121
rect 11946 69056 11952 69120
rect 12016 69056 12032 69120
rect 12096 69056 12112 69120
rect 12176 69056 12192 69120
rect 12256 69056 12262 69120
rect 11946 69055 12262 69056
rect 16946 69120 17262 69121
rect 16946 69056 16952 69120
rect 17016 69056 17032 69120
rect 17096 69056 17112 69120
rect 17176 69056 17192 69120
rect 17256 69056 17262 69120
rect 16946 69055 17262 69056
rect 21946 69120 22262 69121
rect 21946 69056 21952 69120
rect 22016 69056 22032 69120
rect 22096 69056 22112 69120
rect 22176 69056 22192 69120
rect 22256 69056 22262 69120
rect 21946 69055 22262 69056
rect 26946 69120 27262 69121
rect 26946 69056 26952 69120
rect 27016 69056 27032 69120
rect 27096 69056 27112 69120
rect 27176 69056 27192 69120
rect 27256 69056 27262 69120
rect 26946 69055 27262 69056
rect 31946 69120 32262 69121
rect 31946 69056 31952 69120
rect 32016 69056 32032 69120
rect 32096 69056 32112 69120
rect 32176 69056 32192 69120
rect 32256 69056 32262 69120
rect 31946 69055 32262 69056
rect 36946 69120 37262 69121
rect 36946 69056 36952 69120
rect 37016 69056 37032 69120
rect 37096 69056 37112 69120
rect 37176 69056 37192 69120
rect 37256 69056 37262 69120
rect 36946 69055 37262 69056
rect 2606 68576 2922 68577
rect 2606 68512 2612 68576
rect 2676 68512 2692 68576
rect 2756 68512 2772 68576
rect 2836 68512 2852 68576
rect 2916 68512 2922 68576
rect 2606 68511 2922 68512
rect 7606 68576 7922 68577
rect 7606 68512 7612 68576
rect 7676 68512 7692 68576
rect 7756 68512 7772 68576
rect 7836 68512 7852 68576
rect 7916 68512 7922 68576
rect 7606 68511 7922 68512
rect 12606 68576 12922 68577
rect 12606 68512 12612 68576
rect 12676 68512 12692 68576
rect 12756 68512 12772 68576
rect 12836 68512 12852 68576
rect 12916 68512 12922 68576
rect 12606 68511 12922 68512
rect 17606 68576 17922 68577
rect 17606 68512 17612 68576
rect 17676 68512 17692 68576
rect 17756 68512 17772 68576
rect 17836 68512 17852 68576
rect 17916 68512 17922 68576
rect 17606 68511 17922 68512
rect 22606 68576 22922 68577
rect 22606 68512 22612 68576
rect 22676 68512 22692 68576
rect 22756 68512 22772 68576
rect 22836 68512 22852 68576
rect 22916 68512 22922 68576
rect 22606 68511 22922 68512
rect 27606 68576 27922 68577
rect 27606 68512 27612 68576
rect 27676 68512 27692 68576
rect 27756 68512 27772 68576
rect 27836 68512 27852 68576
rect 27916 68512 27922 68576
rect 27606 68511 27922 68512
rect 32606 68576 32922 68577
rect 32606 68512 32612 68576
rect 32676 68512 32692 68576
rect 32756 68512 32772 68576
rect 32836 68512 32852 68576
rect 32916 68512 32922 68576
rect 32606 68511 32922 68512
rect 37606 68576 37922 68577
rect 37606 68512 37612 68576
rect 37676 68512 37692 68576
rect 37756 68512 37772 68576
rect 37836 68512 37852 68576
rect 37916 68512 37922 68576
rect 37606 68511 37922 68512
rect 1946 68032 2262 68033
rect 1946 67968 1952 68032
rect 2016 67968 2032 68032
rect 2096 67968 2112 68032
rect 2176 67968 2192 68032
rect 2256 67968 2262 68032
rect 1946 67967 2262 67968
rect 6946 68032 7262 68033
rect 6946 67968 6952 68032
rect 7016 67968 7032 68032
rect 7096 67968 7112 68032
rect 7176 67968 7192 68032
rect 7256 67968 7262 68032
rect 6946 67967 7262 67968
rect 11946 68032 12262 68033
rect 11946 67968 11952 68032
rect 12016 67968 12032 68032
rect 12096 67968 12112 68032
rect 12176 67968 12192 68032
rect 12256 67968 12262 68032
rect 11946 67967 12262 67968
rect 16946 68032 17262 68033
rect 16946 67968 16952 68032
rect 17016 67968 17032 68032
rect 17096 67968 17112 68032
rect 17176 67968 17192 68032
rect 17256 67968 17262 68032
rect 16946 67967 17262 67968
rect 21946 68032 22262 68033
rect 21946 67968 21952 68032
rect 22016 67968 22032 68032
rect 22096 67968 22112 68032
rect 22176 67968 22192 68032
rect 22256 67968 22262 68032
rect 21946 67967 22262 67968
rect 26946 68032 27262 68033
rect 26946 67968 26952 68032
rect 27016 67968 27032 68032
rect 27096 67968 27112 68032
rect 27176 67968 27192 68032
rect 27256 67968 27262 68032
rect 26946 67967 27262 67968
rect 31946 68032 32262 68033
rect 31946 67968 31952 68032
rect 32016 67968 32032 68032
rect 32096 67968 32112 68032
rect 32176 67968 32192 68032
rect 32256 67968 32262 68032
rect 31946 67967 32262 67968
rect 36946 68032 37262 68033
rect 36946 67968 36952 68032
rect 37016 67968 37032 68032
rect 37096 67968 37112 68032
rect 37176 67968 37192 68032
rect 37256 67968 37262 68032
rect 36946 67967 37262 67968
rect 14958 67764 14964 67828
rect 15028 67826 15034 67828
rect 38009 67826 38075 67829
rect 15028 67824 38075 67826
rect 15028 67768 38014 67824
rect 38070 67768 38075 67824
rect 15028 67766 38075 67768
rect 15028 67764 15034 67766
rect 38009 67763 38075 67766
rect 3366 67628 3372 67692
rect 3436 67690 3442 67692
rect 37089 67690 37155 67693
rect 3436 67688 37155 67690
rect 3436 67632 37094 67688
rect 37150 67632 37155 67688
rect 3436 67630 37155 67632
rect 3436 67628 3442 67630
rect 37089 67627 37155 67630
rect 2606 67488 2922 67489
rect 2606 67424 2612 67488
rect 2676 67424 2692 67488
rect 2756 67424 2772 67488
rect 2836 67424 2852 67488
rect 2916 67424 2922 67488
rect 2606 67423 2922 67424
rect 7606 67488 7922 67489
rect 7606 67424 7612 67488
rect 7676 67424 7692 67488
rect 7756 67424 7772 67488
rect 7836 67424 7852 67488
rect 7916 67424 7922 67488
rect 7606 67423 7922 67424
rect 12606 67488 12922 67489
rect 12606 67424 12612 67488
rect 12676 67424 12692 67488
rect 12756 67424 12772 67488
rect 12836 67424 12852 67488
rect 12916 67424 12922 67488
rect 12606 67423 12922 67424
rect 17606 67488 17922 67489
rect 17606 67424 17612 67488
rect 17676 67424 17692 67488
rect 17756 67424 17772 67488
rect 17836 67424 17852 67488
rect 17916 67424 17922 67488
rect 17606 67423 17922 67424
rect 22606 67488 22922 67489
rect 22606 67424 22612 67488
rect 22676 67424 22692 67488
rect 22756 67424 22772 67488
rect 22836 67424 22852 67488
rect 22916 67424 22922 67488
rect 22606 67423 22922 67424
rect 27606 67488 27922 67489
rect 27606 67424 27612 67488
rect 27676 67424 27692 67488
rect 27756 67424 27772 67488
rect 27836 67424 27852 67488
rect 27916 67424 27922 67488
rect 27606 67423 27922 67424
rect 32606 67488 32922 67489
rect 32606 67424 32612 67488
rect 32676 67424 32692 67488
rect 32756 67424 32772 67488
rect 32836 67424 32852 67488
rect 32916 67424 32922 67488
rect 32606 67423 32922 67424
rect 37606 67488 37922 67489
rect 37606 67424 37612 67488
rect 37676 67424 37692 67488
rect 37756 67424 37772 67488
rect 37836 67424 37852 67488
rect 37916 67424 37922 67488
rect 37606 67423 37922 67424
rect 0 67282 800 67312
rect 1393 67282 1459 67285
rect 0 67280 1459 67282
rect 0 67224 1398 67280
rect 1454 67224 1459 67280
rect 0 67222 1459 67224
rect 0 67192 800 67222
rect 1393 67219 1459 67222
rect 40493 67282 40559 67285
rect 41200 67282 42000 67312
rect 40493 67280 42000 67282
rect 40493 67224 40498 67280
rect 40554 67224 42000 67280
rect 40493 67222 42000 67224
rect 40493 67219 40559 67222
rect 41200 67192 42000 67222
rect 1946 66944 2262 66945
rect 1946 66880 1952 66944
rect 2016 66880 2032 66944
rect 2096 66880 2112 66944
rect 2176 66880 2192 66944
rect 2256 66880 2262 66944
rect 1946 66879 2262 66880
rect 6946 66944 7262 66945
rect 6946 66880 6952 66944
rect 7016 66880 7032 66944
rect 7096 66880 7112 66944
rect 7176 66880 7192 66944
rect 7256 66880 7262 66944
rect 6946 66879 7262 66880
rect 11946 66944 12262 66945
rect 11946 66880 11952 66944
rect 12016 66880 12032 66944
rect 12096 66880 12112 66944
rect 12176 66880 12192 66944
rect 12256 66880 12262 66944
rect 11946 66879 12262 66880
rect 16946 66944 17262 66945
rect 16946 66880 16952 66944
rect 17016 66880 17032 66944
rect 17096 66880 17112 66944
rect 17176 66880 17192 66944
rect 17256 66880 17262 66944
rect 16946 66879 17262 66880
rect 21946 66944 22262 66945
rect 21946 66880 21952 66944
rect 22016 66880 22032 66944
rect 22096 66880 22112 66944
rect 22176 66880 22192 66944
rect 22256 66880 22262 66944
rect 21946 66879 22262 66880
rect 26946 66944 27262 66945
rect 26946 66880 26952 66944
rect 27016 66880 27032 66944
rect 27096 66880 27112 66944
rect 27176 66880 27192 66944
rect 27256 66880 27262 66944
rect 26946 66879 27262 66880
rect 31946 66944 32262 66945
rect 31946 66880 31952 66944
rect 32016 66880 32032 66944
rect 32096 66880 32112 66944
rect 32176 66880 32192 66944
rect 32256 66880 32262 66944
rect 31946 66879 32262 66880
rect 36946 66944 37262 66945
rect 36946 66880 36952 66944
rect 37016 66880 37032 66944
rect 37096 66880 37112 66944
rect 37176 66880 37192 66944
rect 37256 66880 37262 66944
rect 36946 66879 37262 66880
rect 2606 66400 2922 66401
rect 2606 66336 2612 66400
rect 2676 66336 2692 66400
rect 2756 66336 2772 66400
rect 2836 66336 2852 66400
rect 2916 66336 2922 66400
rect 2606 66335 2922 66336
rect 7606 66400 7922 66401
rect 7606 66336 7612 66400
rect 7676 66336 7692 66400
rect 7756 66336 7772 66400
rect 7836 66336 7852 66400
rect 7916 66336 7922 66400
rect 7606 66335 7922 66336
rect 12606 66400 12922 66401
rect 12606 66336 12612 66400
rect 12676 66336 12692 66400
rect 12756 66336 12772 66400
rect 12836 66336 12852 66400
rect 12916 66336 12922 66400
rect 12606 66335 12922 66336
rect 17606 66400 17922 66401
rect 17606 66336 17612 66400
rect 17676 66336 17692 66400
rect 17756 66336 17772 66400
rect 17836 66336 17852 66400
rect 17916 66336 17922 66400
rect 17606 66335 17922 66336
rect 22606 66400 22922 66401
rect 22606 66336 22612 66400
rect 22676 66336 22692 66400
rect 22756 66336 22772 66400
rect 22836 66336 22852 66400
rect 22916 66336 22922 66400
rect 22606 66335 22922 66336
rect 27606 66400 27922 66401
rect 27606 66336 27612 66400
rect 27676 66336 27692 66400
rect 27756 66336 27772 66400
rect 27836 66336 27852 66400
rect 27916 66336 27922 66400
rect 27606 66335 27922 66336
rect 32606 66400 32922 66401
rect 32606 66336 32612 66400
rect 32676 66336 32692 66400
rect 32756 66336 32772 66400
rect 32836 66336 32852 66400
rect 32916 66336 32922 66400
rect 32606 66335 32922 66336
rect 37606 66400 37922 66401
rect 37606 66336 37612 66400
rect 37676 66336 37692 66400
rect 37756 66336 37772 66400
rect 37836 66336 37852 66400
rect 37916 66336 37922 66400
rect 37606 66335 37922 66336
rect 1946 65856 2262 65857
rect 1946 65792 1952 65856
rect 2016 65792 2032 65856
rect 2096 65792 2112 65856
rect 2176 65792 2192 65856
rect 2256 65792 2262 65856
rect 1946 65791 2262 65792
rect 6946 65856 7262 65857
rect 6946 65792 6952 65856
rect 7016 65792 7032 65856
rect 7096 65792 7112 65856
rect 7176 65792 7192 65856
rect 7256 65792 7262 65856
rect 6946 65791 7262 65792
rect 11946 65856 12262 65857
rect 11946 65792 11952 65856
rect 12016 65792 12032 65856
rect 12096 65792 12112 65856
rect 12176 65792 12192 65856
rect 12256 65792 12262 65856
rect 11946 65791 12262 65792
rect 16946 65856 17262 65857
rect 16946 65792 16952 65856
rect 17016 65792 17032 65856
rect 17096 65792 17112 65856
rect 17176 65792 17192 65856
rect 17256 65792 17262 65856
rect 16946 65791 17262 65792
rect 21946 65856 22262 65857
rect 21946 65792 21952 65856
rect 22016 65792 22032 65856
rect 22096 65792 22112 65856
rect 22176 65792 22192 65856
rect 22256 65792 22262 65856
rect 21946 65791 22262 65792
rect 26946 65856 27262 65857
rect 26946 65792 26952 65856
rect 27016 65792 27032 65856
rect 27096 65792 27112 65856
rect 27176 65792 27192 65856
rect 27256 65792 27262 65856
rect 26946 65791 27262 65792
rect 31946 65856 32262 65857
rect 31946 65792 31952 65856
rect 32016 65792 32032 65856
rect 32096 65792 32112 65856
rect 32176 65792 32192 65856
rect 32256 65792 32262 65856
rect 31946 65791 32262 65792
rect 36946 65856 37262 65857
rect 36946 65792 36952 65856
rect 37016 65792 37032 65856
rect 37096 65792 37112 65856
rect 37176 65792 37192 65856
rect 37256 65792 37262 65856
rect 36946 65791 37262 65792
rect 8109 65514 8175 65517
rect 23606 65514 23612 65516
rect 8109 65512 23612 65514
rect 8109 65456 8114 65512
rect 8170 65456 23612 65512
rect 8109 65454 23612 65456
rect 8109 65451 8175 65454
rect 23606 65452 23612 65454
rect 23676 65452 23682 65516
rect 2606 65312 2922 65313
rect 2606 65248 2612 65312
rect 2676 65248 2692 65312
rect 2756 65248 2772 65312
rect 2836 65248 2852 65312
rect 2916 65248 2922 65312
rect 2606 65247 2922 65248
rect 7606 65312 7922 65313
rect 7606 65248 7612 65312
rect 7676 65248 7692 65312
rect 7756 65248 7772 65312
rect 7836 65248 7852 65312
rect 7916 65248 7922 65312
rect 7606 65247 7922 65248
rect 12606 65312 12922 65313
rect 12606 65248 12612 65312
rect 12676 65248 12692 65312
rect 12756 65248 12772 65312
rect 12836 65248 12852 65312
rect 12916 65248 12922 65312
rect 12606 65247 12922 65248
rect 17606 65312 17922 65313
rect 17606 65248 17612 65312
rect 17676 65248 17692 65312
rect 17756 65248 17772 65312
rect 17836 65248 17852 65312
rect 17916 65248 17922 65312
rect 17606 65247 17922 65248
rect 22606 65312 22922 65313
rect 22606 65248 22612 65312
rect 22676 65248 22692 65312
rect 22756 65248 22772 65312
rect 22836 65248 22852 65312
rect 22916 65248 22922 65312
rect 22606 65247 22922 65248
rect 27606 65312 27922 65313
rect 27606 65248 27612 65312
rect 27676 65248 27692 65312
rect 27756 65248 27772 65312
rect 27836 65248 27852 65312
rect 27916 65248 27922 65312
rect 27606 65247 27922 65248
rect 32606 65312 32922 65313
rect 32606 65248 32612 65312
rect 32676 65248 32692 65312
rect 32756 65248 32772 65312
rect 32836 65248 32852 65312
rect 32916 65248 32922 65312
rect 32606 65247 32922 65248
rect 37606 65312 37922 65313
rect 37606 65248 37612 65312
rect 37676 65248 37692 65312
rect 37756 65248 37772 65312
rect 37836 65248 37852 65312
rect 37916 65248 37922 65312
rect 37606 65247 37922 65248
rect 1946 64768 2262 64769
rect 1946 64704 1952 64768
rect 2016 64704 2032 64768
rect 2096 64704 2112 64768
rect 2176 64704 2192 64768
rect 2256 64704 2262 64768
rect 1946 64703 2262 64704
rect 6946 64768 7262 64769
rect 6946 64704 6952 64768
rect 7016 64704 7032 64768
rect 7096 64704 7112 64768
rect 7176 64704 7192 64768
rect 7256 64704 7262 64768
rect 6946 64703 7262 64704
rect 11946 64768 12262 64769
rect 11946 64704 11952 64768
rect 12016 64704 12032 64768
rect 12096 64704 12112 64768
rect 12176 64704 12192 64768
rect 12256 64704 12262 64768
rect 11946 64703 12262 64704
rect 16946 64768 17262 64769
rect 16946 64704 16952 64768
rect 17016 64704 17032 64768
rect 17096 64704 17112 64768
rect 17176 64704 17192 64768
rect 17256 64704 17262 64768
rect 16946 64703 17262 64704
rect 21946 64768 22262 64769
rect 21946 64704 21952 64768
rect 22016 64704 22032 64768
rect 22096 64704 22112 64768
rect 22176 64704 22192 64768
rect 22256 64704 22262 64768
rect 21946 64703 22262 64704
rect 26946 64768 27262 64769
rect 26946 64704 26952 64768
rect 27016 64704 27032 64768
rect 27096 64704 27112 64768
rect 27176 64704 27192 64768
rect 27256 64704 27262 64768
rect 26946 64703 27262 64704
rect 31946 64768 32262 64769
rect 31946 64704 31952 64768
rect 32016 64704 32032 64768
rect 32096 64704 32112 64768
rect 32176 64704 32192 64768
rect 32256 64704 32262 64768
rect 31946 64703 32262 64704
rect 36946 64768 37262 64769
rect 36946 64704 36952 64768
rect 37016 64704 37032 64768
rect 37096 64704 37112 64768
rect 37176 64704 37192 64768
rect 37256 64704 37262 64768
rect 36946 64703 37262 64704
rect 2606 64224 2922 64225
rect 2606 64160 2612 64224
rect 2676 64160 2692 64224
rect 2756 64160 2772 64224
rect 2836 64160 2852 64224
rect 2916 64160 2922 64224
rect 2606 64159 2922 64160
rect 7606 64224 7922 64225
rect 7606 64160 7612 64224
rect 7676 64160 7692 64224
rect 7756 64160 7772 64224
rect 7836 64160 7852 64224
rect 7916 64160 7922 64224
rect 7606 64159 7922 64160
rect 12606 64224 12922 64225
rect 12606 64160 12612 64224
rect 12676 64160 12692 64224
rect 12756 64160 12772 64224
rect 12836 64160 12852 64224
rect 12916 64160 12922 64224
rect 12606 64159 12922 64160
rect 17606 64224 17922 64225
rect 17606 64160 17612 64224
rect 17676 64160 17692 64224
rect 17756 64160 17772 64224
rect 17836 64160 17852 64224
rect 17916 64160 17922 64224
rect 17606 64159 17922 64160
rect 22606 64224 22922 64225
rect 22606 64160 22612 64224
rect 22676 64160 22692 64224
rect 22756 64160 22772 64224
rect 22836 64160 22852 64224
rect 22916 64160 22922 64224
rect 22606 64159 22922 64160
rect 27606 64224 27922 64225
rect 27606 64160 27612 64224
rect 27676 64160 27692 64224
rect 27756 64160 27772 64224
rect 27836 64160 27852 64224
rect 27916 64160 27922 64224
rect 27606 64159 27922 64160
rect 32606 64224 32922 64225
rect 32606 64160 32612 64224
rect 32676 64160 32692 64224
rect 32756 64160 32772 64224
rect 32836 64160 32852 64224
rect 32916 64160 32922 64224
rect 32606 64159 32922 64160
rect 37606 64224 37922 64225
rect 37606 64160 37612 64224
rect 37676 64160 37692 64224
rect 37756 64160 37772 64224
rect 37836 64160 37852 64224
rect 37916 64160 37922 64224
rect 37606 64159 37922 64160
rect 1946 63680 2262 63681
rect 1946 63616 1952 63680
rect 2016 63616 2032 63680
rect 2096 63616 2112 63680
rect 2176 63616 2192 63680
rect 2256 63616 2262 63680
rect 1946 63615 2262 63616
rect 6946 63680 7262 63681
rect 6946 63616 6952 63680
rect 7016 63616 7032 63680
rect 7096 63616 7112 63680
rect 7176 63616 7192 63680
rect 7256 63616 7262 63680
rect 6946 63615 7262 63616
rect 11946 63680 12262 63681
rect 11946 63616 11952 63680
rect 12016 63616 12032 63680
rect 12096 63616 12112 63680
rect 12176 63616 12192 63680
rect 12256 63616 12262 63680
rect 11946 63615 12262 63616
rect 16946 63680 17262 63681
rect 16946 63616 16952 63680
rect 17016 63616 17032 63680
rect 17096 63616 17112 63680
rect 17176 63616 17192 63680
rect 17256 63616 17262 63680
rect 16946 63615 17262 63616
rect 21946 63680 22262 63681
rect 21946 63616 21952 63680
rect 22016 63616 22032 63680
rect 22096 63616 22112 63680
rect 22176 63616 22192 63680
rect 22256 63616 22262 63680
rect 21946 63615 22262 63616
rect 26946 63680 27262 63681
rect 26946 63616 26952 63680
rect 27016 63616 27032 63680
rect 27096 63616 27112 63680
rect 27176 63616 27192 63680
rect 27256 63616 27262 63680
rect 26946 63615 27262 63616
rect 31946 63680 32262 63681
rect 31946 63616 31952 63680
rect 32016 63616 32032 63680
rect 32096 63616 32112 63680
rect 32176 63616 32192 63680
rect 32256 63616 32262 63680
rect 31946 63615 32262 63616
rect 36946 63680 37262 63681
rect 36946 63616 36952 63680
rect 37016 63616 37032 63680
rect 37096 63616 37112 63680
rect 37176 63616 37192 63680
rect 37256 63616 37262 63680
rect 36946 63615 37262 63616
rect 20345 63610 20411 63613
rect 20478 63610 20484 63612
rect 20345 63608 20484 63610
rect 20345 63552 20350 63608
rect 20406 63552 20484 63608
rect 20345 63550 20484 63552
rect 20345 63547 20411 63550
rect 20478 63548 20484 63550
rect 20548 63548 20554 63612
rect 21582 63548 21588 63612
rect 21652 63610 21658 63612
rect 21725 63610 21791 63613
rect 21652 63608 21791 63610
rect 21652 63552 21730 63608
rect 21786 63552 21791 63608
rect 21652 63550 21791 63552
rect 21652 63548 21658 63550
rect 21725 63547 21791 63550
rect 2606 63136 2922 63137
rect 2606 63072 2612 63136
rect 2676 63072 2692 63136
rect 2756 63072 2772 63136
rect 2836 63072 2852 63136
rect 2916 63072 2922 63136
rect 2606 63071 2922 63072
rect 7606 63136 7922 63137
rect 7606 63072 7612 63136
rect 7676 63072 7692 63136
rect 7756 63072 7772 63136
rect 7836 63072 7852 63136
rect 7916 63072 7922 63136
rect 7606 63071 7922 63072
rect 12606 63136 12922 63137
rect 12606 63072 12612 63136
rect 12676 63072 12692 63136
rect 12756 63072 12772 63136
rect 12836 63072 12852 63136
rect 12916 63072 12922 63136
rect 12606 63071 12922 63072
rect 17606 63136 17922 63137
rect 17606 63072 17612 63136
rect 17676 63072 17692 63136
rect 17756 63072 17772 63136
rect 17836 63072 17852 63136
rect 17916 63072 17922 63136
rect 17606 63071 17922 63072
rect 22606 63136 22922 63137
rect 22606 63072 22612 63136
rect 22676 63072 22692 63136
rect 22756 63072 22772 63136
rect 22836 63072 22852 63136
rect 22916 63072 22922 63136
rect 22606 63071 22922 63072
rect 27606 63136 27922 63137
rect 27606 63072 27612 63136
rect 27676 63072 27692 63136
rect 27756 63072 27772 63136
rect 27836 63072 27852 63136
rect 27916 63072 27922 63136
rect 27606 63071 27922 63072
rect 32606 63136 32922 63137
rect 32606 63072 32612 63136
rect 32676 63072 32692 63136
rect 32756 63072 32772 63136
rect 32836 63072 32852 63136
rect 32916 63072 32922 63136
rect 32606 63071 32922 63072
rect 37606 63136 37922 63137
rect 37606 63072 37612 63136
rect 37676 63072 37692 63136
rect 37756 63072 37772 63136
rect 37836 63072 37852 63136
rect 37916 63072 37922 63136
rect 37606 63071 37922 63072
rect 24710 62732 24716 62796
rect 24780 62794 24786 62796
rect 33593 62794 33659 62797
rect 24780 62792 33659 62794
rect 24780 62736 33598 62792
rect 33654 62736 33659 62792
rect 24780 62734 33659 62736
rect 24780 62732 24786 62734
rect 33593 62731 33659 62734
rect 1946 62592 2262 62593
rect 1946 62528 1952 62592
rect 2016 62528 2032 62592
rect 2096 62528 2112 62592
rect 2176 62528 2192 62592
rect 2256 62528 2262 62592
rect 1946 62527 2262 62528
rect 6946 62592 7262 62593
rect 6946 62528 6952 62592
rect 7016 62528 7032 62592
rect 7096 62528 7112 62592
rect 7176 62528 7192 62592
rect 7256 62528 7262 62592
rect 6946 62527 7262 62528
rect 11946 62592 12262 62593
rect 11946 62528 11952 62592
rect 12016 62528 12032 62592
rect 12096 62528 12112 62592
rect 12176 62528 12192 62592
rect 12256 62528 12262 62592
rect 11946 62527 12262 62528
rect 16946 62592 17262 62593
rect 16946 62528 16952 62592
rect 17016 62528 17032 62592
rect 17096 62528 17112 62592
rect 17176 62528 17192 62592
rect 17256 62528 17262 62592
rect 16946 62527 17262 62528
rect 21946 62592 22262 62593
rect 21946 62528 21952 62592
rect 22016 62528 22032 62592
rect 22096 62528 22112 62592
rect 22176 62528 22192 62592
rect 22256 62528 22262 62592
rect 21946 62527 22262 62528
rect 26946 62592 27262 62593
rect 26946 62528 26952 62592
rect 27016 62528 27032 62592
rect 27096 62528 27112 62592
rect 27176 62528 27192 62592
rect 27256 62528 27262 62592
rect 26946 62527 27262 62528
rect 31946 62592 32262 62593
rect 31946 62528 31952 62592
rect 32016 62528 32032 62592
rect 32096 62528 32112 62592
rect 32176 62528 32192 62592
rect 32256 62528 32262 62592
rect 31946 62527 32262 62528
rect 36946 62592 37262 62593
rect 36946 62528 36952 62592
rect 37016 62528 37032 62592
rect 37096 62528 37112 62592
rect 37176 62528 37192 62592
rect 37256 62528 37262 62592
rect 36946 62527 37262 62528
rect 2606 62048 2922 62049
rect 2606 61984 2612 62048
rect 2676 61984 2692 62048
rect 2756 61984 2772 62048
rect 2836 61984 2852 62048
rect 2916 61984 2922 62048
rect 2606 61983 2922 61984
rect 7606 62048 7922 62049
rect 7606 61984 7612 62048
rect 7676 61984 7692 62048
rect 7756 61984 7772 62048
rect 7836 61984 7852 62048
rect 7916 61984 7922 62048
rect 7606 61983 7922 61984
rect 12606 62048 12922 62049
rect 12606 61984 12612 62048
rect 12676 61984 12692 62048
rect 12756 61984 12772 62048
rect 12836 61984 12852 62048
rect 12916 61984 12922 62048
rect 12606 61983 12922 61984
rect 17606 62048 17922 62049
rect 17606 61984 17612 62048
rect 17676 61984 17692 62048
rect 17756 61984 17772 62048
rect 17836 61984 17852 62048
rect 17916 61984 17922 62048
rect 17606 61983 17922 61984
rect 22606 62048 22922 62049
rect 22606 61984 22612 62048
rect 22676 61984 22692 62048
rect 22756 61984 22772 62048
rect 22836 61984 22852 62048
rect 22916 61984 22922 62048
rect 22606 61983 22922 61984
rect 27606 62048 27922 62049
rect 27606 61984 27612 62048
rect 27676 61984 27692 62048
rect 27756 61984 27772 62048
rect 27836 61984 27852 62048
rect 27916 61984 27922 62048
rect 27606 61983 27922 61984
rect 32606 62048 32922 62049
rect 32606 61984 32612 62048
rect 32676 61984 32692 62048
rect 32756 61984 32772 62048
rect 32836 61984 32852 62048
rect 32916 61984 32922 62048
rect 32606 61983 32922 61984
rect 37606 62048 37922 62049
rect 37606 61984 37612 62048
rect 37676 61984 37692 62048
rect 37756 61984 37772 62048
rect 37836 61984 37852 62048
rect 37916 61984 37922 62048
rect 37606 61983 37922 61984
rect 25262 61644 25268 61708
rect 25332 61706 25338 61708
rect 35249 61706 35315 61709
rect 25332 61704 35315 61706
rect 25332 61648 35254 61704
rect 35310 61648 35315 61704
rect 25332 61646 35315 61648
rect 25332 61644 25338 61646
rect 35249 61643 35315 61646
rect 1946 61504 2262 61505
rect 1946 61440 1952 61504
rect 2016 61440 2032 61504
rect 2096 61440 2112 61504
rect 2176 61440 2192 61504
rect 2256 61440 2262 61504
rect 1946 61439 2262 61440
rect 6946 61504 7262 61505
rect 6946 61440 6952 61504
rect 7016 61440 7032 61504
rect 7096 61440 7112 61504
rect 7176 61440 7192 61504
rect 7256 61440 7262 61504
rect 6946 61439 7262 61440
rect 11946 61504 12262 61505
rect 11946 61440 11952 61504
rect 12016 61440 12032 61504
rect 12096 61440 12112 61504
rect 12176 61440 12192 61504
rect 12256 61440 12262 61504
rect 11946 61439 12262 61440
rect 16946 61504 17262 61505
rect 16946 61440 16952 61504
rect 17016 61440 17032 61504
rect 17096 61440 17112 61504
rect 17176 61440 17192 61504
rect 17256 61440 17262 61504
rect 16946 61439 17262 61440
rect 21946 61504 22262 61505
rect 21946 61440 21952 61504
rect 22016 61440 22032 61504
rect 22096 61440 22112 61504
rect 22176 61440 22192 61504
rect 22256 61440 22262 61504
rect 21946 61439 22262 61440
rect 26946 61504 27262 61505
rect 26946 61440 26952 61504
rect 27016 61440 27032 61504
rect 27096 61440 27112 61504
rect 27176 61440 27192 61504
rect 27256 61440 27262 61504
rect 26946 61439 27262 61440
rect 31946 61504 32262 61505
rect 31946 61440 31952 61504
rect 32016 61440 32032 61504
rect 32096 61440 32112 61504
rect 32176 61440 32192 61504
rect 32256 61440 32262 61504
rect 31946 61439 32262 61440
rect 36946 61504 37262 61505
rect 36946 61440 36952 61504
rect 37016 61440 37032 61504
rect 37096 61440 37112 61504
rect 37176 61440 37192 61504
rect 37256 61440 37262 61504
rect 36946 61439 37262 61440
rect 2606 60960 2922 60961
rect 2606 60896 2612 60960
rect 2676 60896 2692 60960
rect 2756 60896 2772 60960
rect 2836 60896 2852 60960
rect 2916 60896 2922 60960
rect 2606 60895 2922 60896
rect 7606 60960 7922 60961
rect 7606 60896 7612 60960
rect 7676 60896 7692 60960
rect 7756 60896 7772 60960
rect 7836 60896 7852 60960
rect 7916 60896 7922 60960
rect 7606 60895 7922 60896
rect 12606 60960 12922 60961
rect 12606 60896 12612 60960
rect 12676 60896 12692 60960
rect 12756 60896 12772 60960
rect 12836 60896 12852 60960
rect 12916 60896 12922 60960
rect 12606 60895 12922 60896
rect 17606 60960 17922 60961
rect 17606 60896 17612 60960
rect 17676 60896 17692 60960
rect 17756 60896 17772 60960
rect 17836 60896 17852 60960
rect 17916 60896 17922 60960
rect 17606 60895 17922 60896
rect 22606 60960 22922 60961
rect 22606 60896 22612 60960
rect 22676 60896 22692 60960
rect 22756 60896 22772 60960
rect 22836 60896 22852 60960
rect 22916 60896 22922 60960
rect 22606 60895 22922 60896
rect 27606 60960 27922 60961
rect 27606 60896 27612 60960
rect 27676 60896 27692 60960
rect 27756 60896 27772 60960
rect 27836 60896 27852 60960
rect 27916 60896 27922 60960
rect 27606 60895 27922 60896
rect 32606 60960 32922 60961
rect 32606 60896 32612 60960
rect 32676 60896 32692 60960
rect 32756 60896 32772 60960
rect 32836 60896 32852 60960
rect 32916 60896 32922 60960
rect 32606 60895 32922 60896
rect 37606 60960 37922 60961
rect 37606 60896 37612 60960
rect 37676 60896 37692 60960
rect 37756 60896 37772 60960
rect 37836 60896 37852 60960
rect 37916 60896 37922 60960
rect 37606 60895 37922 60896
rect 1946 60416 2262 60417
rect 1946 60352 1952 60416
rect 2016 60352 2032 60416
rect 2096 60352 2112 60416
rect 2176 60352 2192 60416
rect 2256 60352 2262 60416
rect 1946 60351 2262 60352
rect 6946 60416 7262 60417
rect 6946 60352 6952 60416
rect 7016 60352 7032 60416
rect 7096 60352 7112 60416
rect 7176 60352 7192 60416
rect 7256 60352 7262 60416
rect 6946 60351 7262 60352
rect 11946 60416 12262 60417
rect 11946 60352 11952 60416
rect 12016 60352 12032 60416
rect 12096 60352 12112 60416
rect 12176 60352 12192 60416
rect 12256 60352 12262 60416
rect 11946 60351 12262 60352
rect 16946 60416 17262 60417
rect 16946 60352 16952 60416
rect 17016 60352 17032 60416
rect 17096 60352 17112 60416
rect 17176 60352 17192 60416
rect 17256 60352 17262 60416
rect 16946 60351 17262 60352
rect 21946 60416 22262 60417
rect 21946 60352 21952 60416
rect 22016 60352 22032 60416
rect 22096 60352 22112 60416
rect 22176 60352 22192 60416
rect 22256 60352 22262 60416
rect 21946 60351 22262 60352
rect 26946 60416 27262 60417
rect 26946 60352 26952 60416
rect 27016 60352 27032 60416
rect 27096 60352 27112 60416
rect 27176 60352 27192 60416
rect 27256 60352 27262 60416
rect 26946 60351 27262 60352
rect 31946 60416 32262 60417
rect 31946 60352 31952 60416
rect 32016 60352 32032 60416
rect 32096 60352 32112 60416
rect 32176 60352 32192 60416
rect 32256 60352 32262 60416
rect 31946 60351 32262 60352
rect 36946 60416 37262 60417
rect 36946 60352 36952 60416
rect 37016 60352 37032 60416
rect 37096 60352 37112 60416
rect 37176 60352 37192 60416
rect 37256 60352 37262 60416
rect 36946 60351 37262 60352
rect 2606 59872 2922 59873
rect 2606 59808 2612 59872
rect 2676 59808 2692 59872
rect 2756 59808 2772 59872
rect 2836 59808 2852 59872
rect 2916 59808 2922 59872
rect 2606 59807 2922 59808
rect 7606 59872 7922 59873
rect 7606 59808 7612 59872
rect 7676 59808 7692 59872
rect 7756 59808 7772 59872
rect 7836 59808 7852 59872
rect 7916 59808 7922 59872
rect 7606 59807 7922 59808
rect 12606 59872 12922 59873
rect 12606 59808 12612 59872
rect 12676 59808 12692 59872
rect 12756 59808 12772 59872
rect 12836 59808 12852 59872
rect 12916 59808 12922 59872
rect 12606 59807 12922 59808
rect 17606 59872 17922 59873
rect 17606 59808 17612 59872
rect 17676 59808 17692 59872
rect 17756 59808 17772 59872
rect 17836 59808 17852 59872
rect 17916 59808 17922 59872
rect 17606 59807 17922 59808
rect 22606 59872 22922 59873
rect 22606 59808 22612 59872
rect 22676 59808 22692 59872
rect 22756 59808 22772 59872
rect 22836 59808 22852 59872
rect 22916 59808 22922 59872
rect 22606 59807 22922 59808
rect 27606 59872 27922 59873
rect 27606 59808 27612 59872
rect 27676 59808 27692 59872
rect 27756 59808 27772 59872
rect 27836 59808 27852 59872
rect 27916 59808 27922 59872
rect 27606 59807 27922 59808
rect 32606 59872 32922 59873
rect 32606 59808 32612 59872
rect 32676 59808 32692 59872
rect 32756 59808 32772 59872
rect 32836 59808 32852 59872
rect 32916 59808 32922 59872
rect 32606 59807 32922 59808
rect 37606 59872 37922 59873
rect 37606 59808 37612 59872
rect 37676 59808 37692 59872
rect 37756 59808 37772 59872
rect 37836 59808 37852 59872
rect 37916 59808 37922 59872
rect 37606 59807 37922 59808
rect 22093 59530 22159 59533
rect 24894 59530 24900 59532
rect 22093 59528 24900 59530
rect 22093 59472 22098 59528
rect 22154 59472 24900 59528
rect 22093 59470 24900 59472
rect 22093 59467 22159 59470
rect 24894 59468 24900 59470
rect 24964 59468 24970 59532
rect 1946 59328 2262 59329
rect 1946 59264 1952 59328
rect 2016 59264 2032 59328
rect 2096 59264 2112 59328
rect 2176 59264 2192 59328
rect 2256 59264 2262 59328
rect 1946 59263 2262 59264
rect 6946 59328 7262 59329
rect 6946 59264 6952 59328
rect 7016 59264 7032 59328
rect 7096 59264 7112 59328
rect 7176 59264 7192 59328
rect 7256 59264 7262 59328
rect 6946 59263 7262 59264
rect 11946 59328 12262 59329
rect 11946 59264 11952 59328
rect 12016 59264 12032 59328
rect 12096 59264 12112 59328
rect 12176 59264 12192 59328
rect 12256 59264 12262 59328
rect 11946 59263 12262 59264
rect 16946 59328 17262 59329
rect 16946 59264 16952 59328
rect 17016 59264 17032 59328
rect 17096 59264 17112 59328
rect 17176 59264 17192 59328
rect 17256 59264 17262 59328
rect 16946 59263 17262 59264
rect 21946 59328 22262 59329
rect 21946 59264 21952 59328
rect 22016 59264 22032 59328
rect 22096 59264 22112 59328
rect 22176 59264 22192 59328
rect 22256 59264 22262 59328
rect 21946 59263 22262 59264
rect 26946 59328 27262 59329
rect 26946 59264 26952 59328
rect 27016 59264 27032 59328
rect 27096 59264 27112 59328
rect 27176 59264 27192 59328
rect 27256 59264 27262 59328
rect 26946 59263 27262 59264
rect 31946 59328 32262 59329
rect 31946 59264 31952 59328
rect 32016 59264 32032 59328
rect 32096 59264 32112 59328
rect 32176 59264 32192 59328
rect 32256 59264 32262 59328
rect 31946 59263 32262 59264
rect 36946 59328 37262 59329
rect 36946 59264 36952 59328
rect 37016 59264 37032 59328
rect 37096 59264 37112 59328
rect 37176 59264 37192 59328
rect 37256 59264 37262 59328
rect 36946 59263 37262 59264
rect 2606 58784 2922 58785
rect 2606 58720 2612 58784
rect 2676 58720 2692 58784
rect 2756 58720 2772 58784
rect 2836 58720 2852 58784
rect 2916 58720 2922 58784
rect 2606 58719 2922 58720
rect 7606 58784 7922 58785
rect 7606 58720 7612 58784
rect 7676 58720 7692 58784
rect 7756 58720 7772 58784
rect 7836 58720 7852 58784
rect 7916 58720 7922 58784
rect 7606 58719 7922 58720
rect 12606 58784 12922 58785
rect 12606 58720 12612 58784
rect 12676 58720 12692 58784
rect 12756 58720 12772 58784
rect 12836 58720 12852 58784
rect 12916 58720 12922 58784
rect 12606 58719 12922 58720
rect 17606 58784 17922 58785
rect 17606 58720 17612 58784
rect 17676 58720 17692 58784
rect 17756 58720 17772 58784
rect 17836 58720 17852 58784
rect 17916 58720 17922 58784
rect 17606 58719 17922 58720
rect 22606 58784 22922 58785
rect 22606 58720 22612 58784
rect 22676 58720 22692 58784
rect 22756 58720 22772 58784
rect 22836 58720 22852 58784
rect 22916 58720 22922 58784
rect 22606 58719 22922 58720
rect 27606 58784 27922 58785
rect 27606 58720 27612 58784
rect 27676 58720 27692 58784
rect 27756 58720 27772 58784
rect 27836 58720 27852 58784
rect 27916 58720 27922 58784
rect 27606 58719 27922 58720
rect 32606 58784 32922 58785
rect 32606 58720 32612 58784
rect 32676 58720 32692 58784
rect 32756 58720 32772 58784
rect 32836 58720 32852 58784
rect 32916 58720 32922 58784
rect 32606 58719 32922 58720
rect 37606 58784 37922 58785
rect 37606 58720 37612 58784
rect 37676 58720 37692 58784
rect 37756 58720 37772 58784
rect 37836 58720 37852 58784
rect 37916 58720 37922 58784
rect 37606 58719 37922 58720
rect 841 58442 907 58445
rect 798 58440 907 58442
rect 798 58384 846 58440
rect 902 58384 907 58440
rect 798 58379 907 58384
rect 798 58336 858 58379
rect 0 58246 858 58336
rect 39941 58306 40007 58309
rect 41200 58306 42000 58336
rect 39941 58304 42000 58306
rect 39941 58248 39946 58304
rect 40002 58248 42000 58304
rect 39941 58246 42000 58248
rect 0 58216 800 58246
rect 39941 58243 40007 58246
rect 1946 58240 2262 58241
rect 1946 58176 1952 58240
rect 2016 58176 2032 58240
rect 2096 58176 2112 58240
rect 2176 58176 2192 58240
rect 2256 58176 2262 58240
rect 1946 58175 2262 58176
rect 6946 58240 7262 58241
rect 6946 58176 6952 58240
rect 7016 58176 7032 58240
rect 7096 58176 7112 58240
rect 7176 58176 7192 58240
rect 7256 58176 7262 58240
rect 6946 58175 7262 58176
rect 11946 58240 12262 58241
rect 11946 58176 11952 58240
rect 12016 58176 12032 58240
rect 12096 58176 12112 58240
rect 12176 58176 12192 58240
rect 12256 58176 12262 58240
rect 11946 58175 12262 58176
rect 16946 58240 17262 58241
rect 16946 58176 16952 58240
rect 17016 58176 17032 58240
rect 17096 58176 17112 58240
rect 17176 58176 17192 58240
rect 17256 58176 17262 58240
rect 16946 58175 17262 58176
rect 21946 58240 22262 58241
rect 21946 58176 21952 58240
rect 22016 58176 22032 58240
rect 22096 58176 22112 58240
rect 22176 58176 22192 58240
rect 22256 58176 22262 58240
rect 21946 58175 22262 58176
rect 26946 58240 27262 58241
rect 26946 58176 26952 58240
rect 27016 58176 27032 58240
rect 27096 58176 27112 58240
rect 27176 58176 27192 58240
rect 27256 58176 27262 58240
rect 26946 58175 27262 58176
rect 31946 58240 32262 58241
rect 31946 58176 31952 58240
rect 32016 58176 32032 58240
rect 32096 58176 32112 58240
rect 32176 58176 32192 58240
rect 32256 58176 32262 58240
rect 31946 58175 32262 58176
rect 36946 58240 37262 58241
rect 36946 58176 36952 58240
rect 37016 58176 37032 58240
rect 37096 58176 37112 58240
rect 37176 58176 37192 58240
rect 37256 58176 37262 58240
rect 41200 58216 42000 58246
rect 36946 58175 37262 58176
rect 2606 57696 2922 57697
rect 2606 57632 2612 57696
rect 2676 57632 2692 57696
rect 2756 57632 2772 57696
rect 2836 57632 2852 57696
rect 2916 57632 2922 57696
rect 2606 57631 2922 57632
rect 7606 57696 7922 57697
rect 7606 57632 7612 57696
rect 7676 57632 7692 57696
rect 7756 57632 7772 57696
rect 7836 57632 7852 57696
rect 7916 57632 7922 57696
rect 7606 57631 7922 57632
rect 12606 57696 12922 57697
rect 12606 57632 12612 57696
rect 12676 57632 12692 57696
rect 12756 57632 12772 57696
rect 12836 57632 12852 57696
rect 12916 57632 12922 57696
rect 12606 57631 12922 57632
rect 17606 57696 17922 57697
rect 17606 57632 17612 57696
rect 17676 57632 17692 57696
rect 17756 57632 17772 57696
rect 17836 57632 17852 57696
rect 17916 57632 17922 57696
rect 17606 57631 17922 57632
rect 22606 57696 22922 57697
rect 22606 57632 22612 57696
rect 22676 57632 22692 57696
rect 22756 57632 22772 57696
rect 22836 57632 22852 57696
rect 22916 57632 22922 57696
rect 22606 57631 22922 57632
rect 27606 57696 27922 57697
rect 27606 57632 27612 57696
rect 27676 57632 27692 57696
rect 27756 57632 27772 57696
rect 27836 57632 27852 57696
rect 27916 57632 27922 57696
rect 27606 57631 27922 57632
rect 32606 57696 32922 57697
rect 32606 57632 32612 57696
rect 32676 57632 32692 57696
rect 32756 57632 32772 57696
rect 32836 57632 32852 57696
rect 32916 57632 32922 57696
rect 32606 57631 32922 57632
rect 37606 57696 37922 57697
rect 37606 57632 37612 57696
rect 37676 57632 37692 57696
rect 37756 57632 37772 57696
rect 37836 57632 37852 57696
rect 37916 57632 37922 57696
rect 37606 57631 37922 57632
rect 1946 57152 2262 57153
rect 1946 57088 1952 57152
rect 2016 57088 2032 57152
rect 2096 57088 2112 57152
rect 2176 57088 2192 57152
rect 2256 57088 2262 57152
rect 1946 57087 2262 57088
rect 6946 57152 7262 57153
rect 6946 57088 6952 57152
rect 7016 57088 7032 57152
rect 7096 57088 7112 57152
rect 7176 57088 7192 57152
rect 7256 57088 7262 57152
rect 6946 57087 7262 57088
rect 11946 57152 12262 57153
rect 11946 57088 11952 57152
rect 12016 57088 12032 57152
rect 12096 57088 12112 57152
rect 12176 57088 12192 57152
rect 12256 57088 12262 57152
rect 11946 57087 12262 57088
rect 16946 57152 17262 57153
rect 16946 57088 16952 57152
rect 17016 57088 17032 57152
rect 17096 57088 17112 57152
rect 17176 57088 17192 57152
rect 17256 57088 17262 57152
rect 16946 57087 17262 57088
rect 21946 57152 22262 57153
rect 21946 57088 21952 57152
rect 22016 57088 22032 57152
rect 22096 57088 22112 57152
rect 22176 57088 22192 57152
rect 22256 57088 22262 57152
rect 21946 57087 22262 57088
rect 26946 57152 27262 57153
rect 26946 57088 26952 57152
rect 27016 57088 27032 57152
rect 27096 57088 27112 57152
rect 27176 57088 27192 57152
rect 27256 57088 27262 57152
rect 26946 57087 27262 57088
rect 31946 57152 32262 57153
rect 31946 57088 31952 57152
rect 32016 57088 32032 57152
rect 32096 57088 32112 57152
rect 32176 57088 32192 57152
rect 32256 57088 32262 57152
rect 31946 57087 32262 57088
rect 36946 57152 37262 57153
rect 36946 57088 36952 57152
rect 37016 57088 37032 57152
rect 37096 57088 37112 57152
rect 37176 57088 37192 57152
rect 37256 57088 37262 57152
rect 36946 57087 37262 57088
rect 10777 56810 10843 56813
rect 18454 56810 18460 56812
rect 10777 56808 18460 56810
rect 10777 56752 10782 56808
rect 10838 56752 18460 56808
rect 10777 56750 18460 56752
rect 10777 56747 10843 56750
rect 18454 56748 18460 56750
rect 18524 56748 18530 56812
rect 2606 56608 2922 56609
rect 2606 56544 2612 56608
rect 2676 56544 2692 56608
rect 2756 56544 2772 56608
rect 2836 56544 2852 56608
rect 2916 56544 2922 56608
rect 2606 56543 2922 56544
rect 7606 56608 7922 56609
rect 7606 56544 7612 56608
rect 7676 56544 7692 56608
rect 7756 56544 7772 56608
rect 7836 56544 7852 56608
rect 7916 56544 7922 56608
rect 7606 56543 7922 56544
rect 12606 56608 12922 56609
rect 12606 56544 12612 56608
rect 12676 56544 12692 56608
rect 12756 56544 12772 56608
rect 12836 56544 12852 56608
rect 12916 56544 12922 56608
rect 12606 56543 12922 56544
rect 17606 56608 17922 56609
rect 17606 56544 17612 56608
rect 17676 56544 17692 56608
rect 17756 56544 17772 56608
rect 17836 56544 17852 56608
rect 17916 56544 17922 56608
rect 17606 56543 17922 56544
rect 22606 56608 22922 56609
rect 22606 56544 22612 56608
rect 22676 56544 22692 56608
rect 22756 56544 22772 56608
rect 22836 56544 22852 56608
rect 22916 56544 22922 56608
rect 22606 56543 22922 56544
rect 27606 56608 27922 56609
rect 27606 56544 27612 56608
rect 27676 56544 27692 56608
rect 27756 56544 27772 56608
rect 27836 56544 27852 56608
rect 27916 56544 27922 56608
rect 27606 56543 27922 56544
rect 32606 56608 32922 56609
rect 32606 56544 32612 56608
rect 32676 56544 32692 56608
rect 32756 56544 32772 56608
rect 32836 56544 32852 56608
rect 32916 56544 32922 56608
rect 32606 56543 32922 56544
rect 37606 56608 37922 56609
rect 37606 56544 37612 56608
rect 37676 56544 37692 56608
rect 37756 56544 37772 56608
rect 37836 56544 37852 56608
rect 37916 56544 37922 56608
rect 37606 56543 37922 56544
rect 1946 56064 2262 56065
rect 1946 56000 1952 56064
rect 2016 56000 2032 56064
rect 2096 56000 2112 56064
rect 2176 56000 2192 56064
rect 2256 56000 2262 56064
rect 1946 55999 2262 56000
rect 6946 56064 7262 56065
rect 6946 56000 6952 56064
rect 7016 56000 7032 56064
rect 7096 56000 7112 56064
rect 7176 56000 7192 56064
rect 7256 56000 7262 56064
rect 6946 55999 7262 56000
rect 11946 56064 12262 56065
rect 11946 56000 11952 56064
rect 12016 56000 12032 56064
rect 12096 56000 12112 56064
rect 12176 56000 12192 56064
rect 12256 56000 12262 56064
rect 11946 55999 12262 56000
rect 16946 56064 17262 56065
rect 16946 56000 16952 56064
rect 17016 56000 17032 56064
rect 17096 56000 17112 56064
rect 17176 56000 17192 56064
rect 17256 56000 17262 56064
rect 16946 55999 17262 56000
rect 21946 56064 22262 56065
rect 21946 56000 21952 56064
rect 22016 56000 22032 56064
rect 22096 56000 22112 56064
rect 22176 56000 22192 56064
rect 22256 56000 22262 56064
rect 21946 55999 22262 56000
rect 26946 56064 27262 56065
rect 26946 56000 26952 56064
rect 27016 56000 27032 56064
rect 27096 56000 27112 56064
rect 27176 56000 27192 56064
rect 27256 56000 27262 56064
rect 26946 55999 27262 56000
rect 31946 56064 32262 56065
rect 31946 56000 31952 56064
rect 32016 56000 32032 56064
rect 32096 56000 32112 56064
rect 32176 56000 32192 56064
rect 32256 56000 32262 56064
rect 31946 55999 32262 56000
rect 36946 56064 37262 56065
rect 36946 56000 36952 56064
rect 37016 56000 37032 56064
rect 37096 56000 37112 56064
rect 37176 56000 37192 56064
rect 37256 56000 37262 56064
rect 36946 55999 37262 56000
rect 2606 55520 2922 55521
rect 2606 55456 2612 55520
rect 2676 55456 2692 55520
rect 2756 55456 2772 55520
rect 2836 55456 2852 55520
rect 2916 55456 2922 55520
rect 2606 55455 2922 55456
rect 7606 55520 7922 55521
rect 7606 55456 7612 55520
rect 7676 55456 7692 55520
rect 7756 55456 7772 55520
rect 7836 55456 7852 55520
rect 7916 55456 7922 55520
rect 7606 55455 7922 55456
rect 12606 55520 12922 55521
rect 12606 55456 12612 55520
rect 12676 55456 12692 55520
rect 12756 55456 12772 55520
rect 12836 55456 12852 55520
rect 12916 55456 12922 55520
rect 12606 55455 12922 55456
rect 17606 55520 17922 55521
rect 17606 55456 17612 55520
rect 17676 55456 17692 55520
rect 17756 55456 17772 55520
rect 17836 55456 17852 55520
rect 17916 55456 17922 55520
rect 17606 55455 17922 55456
rect 22606 55520 22922 55521
rect 22606 55456 22612 55520
rect 22676 55456 22692 55520
rect 22756 55456 22772 55520
rect 22836 55456 22852 55520
rect 22916 55456 22922 55520
rect 22606 55455 22922 55456
rect 27606 55520 27922 55521
rect 27606 55456 27612 55520
rect 27676 55456 27692 55520
rect 27756 55456 27772 55520
rect 27836 55456 27852 55520
rect 27916 55456 27922 55520
rect 27606 55455 27922 55456
rect 32606 55520 32922 55521
rect 32606 55456 32612 55520
rect 32676 55456 32692 55520
rect 32756 55456 32772 55520
rect 32836 55456 32852 55520
rect 32916 55456 32922 55520
rect 32606 55455 32922 55456
rect 37606 55520 37922 55521
rect 37606 55456 37612 55520
rect 37676 55456 37692 55520
rect 37756 55456 37772 55520
rect 37836 55456 37852 55520
rect 37916 55456 37922 55520
rect 37606 55455 37922 55456
rect 16481 55316 16547 55317
rect 16430 55314 16436 55316
rect 16390 55254 16436 55314
rect 16500 55312 16547 55316
rect 16542 55256 16547 55312
rect 16430 55252 16436 55254
rect 16500 55252 16547 55256
rect 16481 55251 16547 55252
rect 1946 54976 2262 54977
rect 1946 54912 1952 54976
rect 2016 54912 2032 54976
rect 2096 54912 2112 54976
rect 2176 54912 2192 54976
rect 2256 54912 2262 54976
rect 1946 54911 2262 54912
rect 6946 54976 7262 54977
rect 6946 54912 6952 54976
rect 7016 54912 7032 54976
rect 7096 54912 7112 54976
rect 7176 54912 7192 54976
rect 7256 54912 7262 54976
rect 6946 54911 7262 54912
rect 11946 54976 12262 54977
rect 11946 54912 11952 54976
rect 12016 54912 12032 54976
rect 12096 54912 12112 54976
rect 12176 54912 12192 54976
rect 12256 54912 12262 54976
rect 11946 54911 12262 54912
rect 16946 54976 17262 54977
rect 16946 54912 16952 54976
rect 17016 54912 17032 54976
rect 17096 54912 17112 54976
rect 17176 54912 17192 54976
rect 17256 54912 17262 54976
rect 16946 54911 17262 54912
rect 21946 54976 22262 54977
rect 21946 54912 21952 54976
rect 22016 54912 22032 54976
rect 22096 54912 22112 54976
rect 22176 54912 22192 54976
rect 22256 54912 22262 54976
rect 21946 54911 22262 54912
rect 26946 54976 27262 54977
rect 26946 54912 26952 54976
rect 27016 54912 27032 54976
rect 27096 54912 27112 54976
rect 27176 54912 27192 54976
rect 27256 54912 27262 54976
rect 26946 54911 27262 54912
rect 31946 54976 32262 54977
rect 31946 54912 31952 54976
rect 32016 54912 32032 54976
rect 32096 54912 32112 54976
rect 32176 54912 32192 54976
rect 32256 54912 32262 54976
rect 31946 54911 32262 54912
rect 36946 54976 37262 54977
rect 36946 54912 36952 54976
rect 37016 54912 37032 54976
rect 37096 54912 37112 54976
rect 37176 54912 37192 54976
rect 37256 54912 37262 54976
rect 36946 54911 37262 54912
rect 2606 54432 2922 54433
rect 2606 54368 2612 54432
rect 2676 54368 2692 54432
rect 2756 54368 2772 54432
rect 2836 54368 2852 54432
rect 2916 54368 2922 54432
rect 2606 54367 2922 54368
rect 7606 54432 7922 54433
rect 7606 54368 7612 54432
rect 7676 54368 7692 54432
rect 7756 54368 7772 54432
rect 7836 54368 7852 54432
rect 7916 54368 7922 54432
rect 7606 54367 7922 54368
rect 12606 54432 12922 54433
rect 12606 54368 12612 54432
rect 12676 54368 12692 54432
rect 12756 54368 12772 54432
rect 12836 54368 12852 54432
rect 12916 54368 12922 54432
rect 12606 54367 12922 54368
rect 17606 54432 17922 54433
rect 17606 54368 17612 54432
rect 17676 54368 17692 54432
rect 17756 54368 17772 54432
rect 17836 54368 17852 54432
rect 17916 54368 17922 54432
rect 17606 54367 17922 54368
rect 22606 54432 22922 54433
rect 22606 54368 22612 54432
rect 22676 54368 22692 54432
rect 22756 54368 22772 54432
rect 22836 54368 22852 54432
rect 22916 54368 22922 54432
rect 22606 54367 22922 54368
rect 27606 54432 27922 54433
rect 27606 54368 27612 54432
rect 27676 54368 27692 54432
rect 27756 54368 27772 54432
rect 27836 54368 27852 54432
rect 27916 54368 27922 54432
rect 27606 54367 27922 54368
rect 32606 54432 32922 54433
rect 32606 54368 32612 54432
rect 32676 54368 32692 54432
rect 32756 54368 32772 54432
rect 32836 54368 32852 54432
rect 32916 54368 32922 54432
rect 32606 54367 32922 54368
rect 37606 54432 37922 54433
rect 37606 54368 37612 54432
rect 37676 54368 37692 54432
rect 37756 54368 37772 54432
rect 37836 54368 37852 54432
rect 37916 54368 37922 54432
rect 37606 54367 37922 54368
rect 1946 53888 2262 53889
rect 1946 53824 1952 53888
rect 2016 53824 2032 53888
rect 2096 53824 2112 53888
rect 2176 53824 2192 53888
rect 2256 53824 2262 53888
rect 1946 53823 2262 53824
rect 6946 53888 7262 53889
rect 6946 53824 6952 53888
rect 7016 53824 7032 53888
rect 7096 53824 7112 53888
rect 7176 53824 7192 53888
rect 7256 53824 7262 53888
rect 6946 53823 7262 53824
rect 11946 53888 12262 53889
rect 11946 53824 11952 53888
rect 12016 53824 12032 53888
rect 12096 53824 12112 53888
rect 12176 53824 12192 53888
rect 12256 53824 12262 53888
rect 11946 53823 12262 53824
rect 16946 53888 17262 53889
rect 16946 53824 16952 53888
rect 17016 53824 17032 53888
rect 17096 53824 17112 53888
rect 17176 53824 17192 53888
rect 17256 53824 17262 53888
rect 16946 53823 17262 53824
rect 21946 53888 22262 53889
rect 21946 53824 21952 53888
rect 22016 53824 22032 53888
rect 22096 53824 22112 53888
rect 22176 53824 22192 53888
rect 22256 53824 22262 53888
rect 21946 53823 22262 53824
rect 26946 53888 27262 53889
rect 26946 53824 26952 53888
rect 27016 53824 27032 53888
rect 27096 53824 27112 53888
rect 27176 53824 27192 53888
rect 27256 53824 27262 53888
rect 26946 53823 27262 53824
rect 31946 53888 32262 53889
rect 31946 53824 31952 53888
rect 32016 53824 32032 53888
rect 32096 53824 32112 53888
rect 32176 53824 32192 53888
rect 32256 53824 32262 53888
rect 31946 53823 32262 53824
rect 36946 53888 37262 53889
rect 36946 53824 36952 53888
rect 37016 53824 37032 53888
rect 37096 53824 37112 53888
rect 37176 53824 37192 53888
rect 37256 53824 37262 53888
rect 36946 53823 37262 53824
rect 2606 53344 2922 53345
rect 2606 53280 2612 53344
rect 2676 53280 2692 53344
rect 2756 53280 2772 53344
rect 2836 53280 2852 53344
rect 2916 53280 2922 53344
rect 2606 53279 2922 53280
rect 7606 53344 7922 53345
rect 7606 53280 7612 53344
rect 7676 53280 7692 53344
rect 7756 53280 7772 53344
rect 7836 53280 7852 53344
rect 7916 53280 7922 53344
rect 7606 53279 7922 53280
rect 12606 53344 12922 53345
rect 12606 53280 12612 53344
rect 12676 53280 12692 53344
rect 12756 53280 12772 53344
rect 12836 53280 12852 53344
rect 12916 53280 12922 53344
rect 12606 53279 12922 53280
rect 17606 53344 17922 53345
rect 17606 53280 17612 53344
rect 17676 53280 17692 53344
rect 17756 53280 17772 53344
rect 17836 53280 17852 53344
rect 17916 53280 17922 53344
rect 17606 53279 17922 53280
rect 22606 53344 22922 53345
rect 22606 53280 22612 53344
rect 22676 53280 22692 53344
rect 22756 53280 22772 53344
rect 22836 53280 22852 53344
rect 22916 53280 22922 53344
rect 22606 53279 22922 53280
rect 27606 53344 27922 53345
rect 27606 53280 27612 53344
rect 27676 53280 27692 53344
rect 27756 53280 27772 53344
rect 27836 53280 27852 53344
rect 27916 53280 27922 53344
rect 27606 53279 27922 53280
rect 32606 53344 32922 53345
rect 32606 53280 32612 53344
rect 32676 53280 32692 53344
rect 32756 53280 32772 53344
rect 32836 53280 32852 53344
rect 32916 53280 32922 53344
rect 32606 53279 32922 53280
rect 37606 53344 37922 53345
rect 37606 53280 37612 53344
rect 37676 53280 37692 53344
rect 37756 53280 37772 53344
rect 37836 53280 37852 53344
rect 37916 53280 37922 53344
rect 37606 53279 37922 53280
rect 1946 52800 2262 52801
rect 1946 52736 1952 52800
rect 2016 52736 2032 52800
rect 2096 52736 2112 52800
rect 2176 52736 2192 52800
rect 2256 52736 2262 52800
rect 1946 52735 2262 52736
rect 6946 52800 7262 52801
rect 6946 52736 6952 52800
rect 7016 52736 7032 52800
rect 7096 52736 7112 52800
rect 7176 52736 7192 52800
rect 7256 52736 7262 52800
rect 6946 52735 7262 52736
rect 11946 52800 12262 52801
rect 11946 52736 11952 52800
rect 12016 52736 12032 52800
rect 12096 52736 12112 52800
rect 12176 52736 12192 52800
rect 12256 52736 12262 52800
rect 11946 52735 12262 52736
rect 16946 52800 17262 52801
rect 16946 52736 16952 52800
rect 17016 52736 17032 52800
rect 17096 52736 17112 52800
rect 17176 52736 17192 52800
rect 17256 52736 17262 52800
rect 16946 52735 17262 52736
rect 21946 52800 22262 52801
rect 21946 52736 21952 52800
rect 22016 52736 22032 52800
rect 22096 52736 22112 52800
rect 22176 52736 22192 52800
rect 22256 52736 22262 52800
rect 21946 52735 22262 52736
rect 26946 52800 27262 52801
rect 26946 52736 26952 52800
rect 27016 52736 27032 52800
rect 27096 52736 27112 52800
rect 27176 52736 27192 52800
rect 27256 52736 27262 52800
rect 26946 52735 27262 52736
rect 31946 52800 32262 52801
rect 31946 52736 31952 52800
rect 32016 52736 32032 52800
rect 32096 52736 32112 52800
rect 32176 52736 32192 52800
rect 32256 52736 32262 52800
rect 31946 52735 32262 52736
rect 36946 52800 37262 52801
rect 36946 52736 36952 52800
rect 37016 52736 37032 52800
rect 37096 52736 37112 52800
rect 37176 52736 37192 52800
rect 37256 52736 37262 52800
rect 36946 52735 37262 52736
rect 2606 52256 2922 52257
rect 2606 52192 2612 52256
rect 2676 52192 2692 52256
rect 2756 52192 2772 52256
rect 2836 52192 2852 52256
rect 2916 52192 2922 52256
rect 2606 52191 2922 52192
rect 7606 52256 7922 52257
rect 7606 52192 7612 52256
rect 7676 52192 7692 52256
rect 7756 52192 7772 52256
rect 7836 52192 7852 52256
rect 7916 52192 7922 52256
rect 7606 52191 7922 52192
rect 12606 52256 12922 52257
rect 12606 52192 12612 52256
rect 12676 52192 12692 52256
rect 12756 52192 12772 52256
rect 12836 52192 12852 52256
rect 12916 52192 12922 52256
rect 12606 52191 12922 52192
rect 17606 52256 17922 52257
rect 17606 52192 17612 52256
rect 17676 52192 17692 52256
rect 17756 52192 17772 52256
rect 17836 52192 17852 52256
rect 17916 52192 17922 52256
rect 17606 52191 17922 52192
rect 22606 52256 22922 52257
rect 22606 52192 22612 52256
rect 22676 52192 22692 52256
rect 22756 52192 22772 52256
rect 22836 52192 22852 52256
rect 22916 52192 22922 52256
rect 22606 52191 22922 52192
rect 27606 52256 27922 52257
rect 27606 52192 27612 52256
rect 27676 52192 27692 52256
rect 27756 52192 27772 52256
rect 27836 52192 27852 52256
rect 27916 52192 27922 52256
rect 27606 52191 27922 52192
rect 32606 52256 32922 52257
rect 32606 52192 32612 52256
rect 32676 52192 32692 52256
rect 32756 52192 32772 52256
rect 32836 52192 32852 52256
rect 32916 52192 32922 52256
rect 32606 52191 32922 52192
rect 37606 52256 37922 52257
rect 37606 52192 37612 52256
rect 37676 52192 37692 52256
rect 37756 52192 37772 52256
rect 37836 52192 37852 52256
rect 37916 52192 37922 52256
rect 37606 52191 37922 52192
rect 20621 52050 20687 52053
rect 21449 52050 21515 52053
rect 20621 52048 21515 52050
rect 20621 51992 20626 52048
rect 20682 51992 21454 52048
rect 21510 51992 21515 52048
rect 20621 51990 21515 51992
rect 20621 51987 20687 51990
rect 21449 51987 21515 51990
rect 1946 51712 2262 51713
rect 1946 51648 1952 51712
rect 2016 51648 2032 51712
rect 2096 51648 2112 51712
rect 2176 51648 2192 51712
rect 2256 51648 2262 51712
rect 1946 51647 2262 51648
rect 6946 51712 7262 51713
rect 6946 51648 6952 51712
rect 7016 51648 7032 51712
rect 7096 51648 7112 51712
rect 7176 51648 7192 51712
rect 7256 51648 7262 51712
rect 6946 51647 7262 51648
rect 11946 51712 12262 51713
rect 11946 51648 11952 51712
rect 12016 51648 12032 51712
rect 12096 51648 12112 51712
rect 12176 51648 12192 51712
rect 12256 51648 12262 51712
rect 11946 51647 12262 51648
rect 16946 51712 17262 51713
rect 16946 51648 16952 51712
rect 17016 51648 17032 51712
rect 17096 51648 17112 51712
rect 17176 51648 17192 51712
rect 17256 51648 17262 51712
rect 16946 51647 17262 51648
rect 21946 51712 22262 51713
rect 21946 51648 21952 51712
rect 22016 51648 22032 51712
rect 22096 51648 22112 51712
rect 22176 51648 22192 51712
rect 22256 51648 22262 51712
rect 21946 51647 22262 51648
rect 26946 51712 27262 51713
rect 26946 51648 26952 51712
rect 27016 51648 27032 51712
rect 27096 51648 27112 51712
rect 27176 51648 27192 51712
rect 27256 51648 27262 51712
rect 26946 51647 27262 51648
rect 31946 51712 32262 51713
rect 31946 51648 31952 51712
rect 32016 51648 32032 51712
rect 32096 51648 32112 51712
rect 32176 51648 32192 51712
rect 32256 51648 32262 51712
rect 31946 51647 32262 51648
rect 36946 51712 37262 51713
rect 36946 51648 36952 51712
rect 37016 51648 37032 51712
rect 37096 51648 37112 51712
rect 37176 51648 37192 51712
rect 37256 51648 37262 51712
rect 36946 51647 37262 51648
rect 2606 51168 2922 51169
rect 2606 51104 2612 51168
rect 2676 51104 2692 51168
rect 2756 51104 2772 51168
rect 2836 51104 2852 51168
rect 2916 51104 2922 51168
rect 2606 51103 2922 51104
rect 7606 51168 7922 51169
rect 7606 51104 7612 51168
rect 7676 51104 7692 51168
rect 7756 51104 7772 51168
rect 7836 51104 7852 51168
rect 7916 51104 7922 51168
rect 7606 51103 7922 51104
rect 12606 51168 12922 51169
rect 12606 51104 12612 51168
rect 12676 51104 12692 51168
rect 12756 51104 12772 51168
rect 12836 51104 12852 51168
rect 12916 51104 12922 51168
rect 12606 51103 12922 51104
rect 17606 51168 17922 51169
rect 17606 51104 17612 51168
rect 17676 51104 17692 51168
rect 17756 51104 17772 51168
rect 17836 51104 17852 51168
rect 17916 51104 17922 51168
rect 17606 51103 17922 51104
rect 22606 51168 22922 51169
rect 22606 51104 22612 51168
rect 22676 51104 22692 51168
rect 22756 51104 22772 51168
rect 22836 51104 22852 51168
rect 22916 51104 22922 51168
rect 22606 51103 22922 51104
rect 27606 51168 27922 51169
rect 27606 51104 27612 51168
rect 27676 51104 27692 51168
rect 27756 51104 27772 51168
rect 27836 51104 27852 51168
rect 27916 51104 27922 51168
rect 27606 51103 27922 51104
rect 32606 51168 32922 51169
rect 32606 51104 32612 51168
rect 32676 51104 32692 51168
rect 32756 51104 32772 51168
rect 32836 51104 32852 51168
rect 32916 51104 32922 51168
rect 32606 51103 32922 51104
rect 37606 51168 37922 51169
rect 37606 51104 37612 51168
rect 37676 51104 37692 51168
rect 37756 51104 37772 51168
rect 37836 51104 37852 51168
rect 37916 51104 37922 51168
rect 37606 51103 37922 51104
rect 34697 51098 34763 51101
rect 34830 51098 34836 51100
rect 34697 51096 34836 51098
rect 34697 51040 34702 51096
rect 34758 51040 34836 51096
rect 34697 51038 34836 51040
rect 34697 51035 34763 51038
rect 34830 51036 34836 51038
rect 34900 51036 34906 51100
rect 1946 50624 2262 50625
rect 1946 50560 1952 50624
rect 2016 50560 2032 50624
rect 2096 50560 2112 50624
rect 2176 50560 2192 50624
rect 2256 50560 2262 50624
rect 1946 50559 2262 50560
rect 6946 50624 7262 50625
rect 6946 50560 6952 50624
rect 7016 50560 7032 50624
rect 7096 50560 7112 50624
rect 7176 50560 7192 50624
rect 7256 50560 7262 50624
rect 6946 50559 7262 50560
rect 11946 50624 12262 50625
rect 11946 50560 11952 50624
rect 12016 50560 12032 50624
rect 12096 50560 12112 50624
rect 12176 50560 12192 50624
rect 12256 50560 12262 50624
rect 11946 50559 12262 50560
rect 16946 50624 17262 50625
rect 16946 50560 16952 50624
rect 17016 50560 17032 50624
rect 17096 50560 17112 50624
rect 17176 50560 17192 50624
rect 17256 50560 17262 50624
rect 16946 50559 17262 50560
rect 21946 50624 22262 50625
rect 21946 50560 21952 50624
rect 22016 50560 22032 50624
rect 22096 50560 22112 50624
rect 22176 50560 22192 50624
rect 22256 50560 22262 50624
rect 21946 50559 22262 50560
rect 26946 50624 27262 50625
rect 26946 50560 26952 50624
rect 27016 50560 27032 50624
rect 27096 50560 27112 50624
rect 27176 50560 27192 50624
rect 27256 50560 27262 50624
rect 26946 50559 27262 50560
rect 31946 50624 32262 50625
rect 31946 50560 31952 50624
rect 32016 50560 32032 50624
rect 32096 50560 32112 50624
rect 32176 50560 32192 50624
rect 32256 50560 32262 50624
rect 31946 50559 32262 50560
rect 36946 50624 37262 50625
rect 36946 50560 36952 50624
rect 37016 50560 37032 50624
rect 37096 50560 37112 50624
rect 37176 50560 37192 50624
rect 37256 50560 37262 50624
rect 36946 50559 37262 50560
rect 2606 50080 2922 50081
rect 2606 50016 2612 50080
rect 2676 50016 2692 50080
rect 2756 50016 2772 50080
rect 2836 50016 2852 50080
rect 2916 50016 2922 50080
rect 2606 50015 2922 50016
rect 7606 50080 7922 50081
rect 7606 50016 7612 50080
rect 7676 50016 7692 50080
rect 7756 50016 7772 50080
rect 7836 50016 7852 50080
rect 7916 50016 7922 50080
rect 7606 50015 7922 50016
rect 12606 50080 12922 50081
rect 12606 50016 12612 50080
rect 12676 50016 12692 50080
rect 12756 50016 12772 50080
rect 12836 50016 12852 50080
rect 12916 50016 12922 50080
rect 12606 50015 12922 50016
rect 17606 50080 17922 50081
rect 17606 50016 17612 50080
rect 17676 50016 17692 50080
rect 17756 50016 17772 50080
rect 17836 50016 17852 50080
rect 17916 50016 17922 50080
rect 17606 50015 17922 50016
rect 22606 50080 22922 50081
rect 22606 50016 22612 50080
rect 22676 50016 22692 50080
rect 22756 50016 22772 50080
rect 22836 50016 22852 50080
rect 22916 50016 22922 50080
rect 22606 50015 22922 50016
rect 27606 50080 27922 50081
rect 27606 50016 27612 50080
rect 27676 50016 27692 50080
rect 27756 50016 27772 50080
rect 27836 50016 27852 50080
rect 27916 50016 27922 50080
rect 27606 50015 27922 50016
rect 32606 50080 32922 50081
rect 32606 50016 32612 50080
rect 32676 50016 32692 50080
rect 32756 50016 32772 50080
rect 32836 50016 32852 50080
rect 32916 50016 32922 50080
rect 32606 50015 32922 50016
rect 37606 50080 37922 50081
rect 37606 50016 37612 50080
rect 37676 50016 37692 50080
rect 37756 50016 37772 50080
rect 37836 50016 37852 50080
rect 37916 50016 37922 50080
rect 37606 50015 37922 50016
rect 1946 49536 2262 49537
rect 1946 49472 1952 49536
rect 2016 49472 2032 49536
rect 2096 49472 2112 49536
rect 2176 49472 2192 49536
rect 2256 49472 2262 49536
rect 1946 49471 2262 49472
rect 6946 49536 7262 49537
rect 6946 49472 6952 49536
rect 7016 49472 7032 49536
rect 7096 49472 7112 49536
rect 7176 49472 7192 49536
rect 7256 49472 7262 49536
rect 6946 49471 7262 49472
rect 11946 49536 12262 49537
rect 11946 49472 11952 49536
rect 12016 49472 12032 49536
rect 12096 49472 12112 49536
rect 12176 49472 12192 49536
rect 12256 49472 12262 49536
rect 11946 49471 12262 49472
rect 16946 49536 17262 49537
rect 16946 49472 16952 49536
rect 17016 49472 17032 49536
rect 17096 49472 17112 49536
rect 17176 49472 17192 49536
rect 17256 49472 17262 49536
rect 16946 49471 17262 49472
rect 21946 49536 22262 49537
rect 21946 49472 21952 49536
rect 22016 49472 22032 49536
rect 22096 49472 22112 49536
rect 22176 49472 22192 49536
rect 22256 49472 22262 49536
rect 21946 49471 22262 49472
rect 26946 49536 27262 49537
rect 26946 49472 26952 49536
rect 27016 49472 27032 49536
rect 27096 49472 27112 49536
rect 27176 49472 27192 49536
rect 27256 49472 27262 49536
rect 26946 49471 27262 49472
rect 31946 49536 32262 49537
rect 31946 49472 31952 49536
rect 32016 49472 32032 49536
rect 32096 49472 32112 49536
rect 32176 49472 32192 49536
rect 32256 49472 32262 49536
rect 31946 49471 32262 49472
rect 36946 49536 37262 49537
rect 36946 49472 36952 49536
rect 37016 49472 37032 49536
rect 37096 49472 37112 49536
rect 37176 49472 37192 49536
rect 37256 49472 37262 49536
rect 36946 49471 37262 49472
rect 0 49330 800 49360
rect 1393 49330 1459 49333
rect 0 49328 1459 49330
rect 0 49272 1398 49328
rect 1454 49272 1459 49328
rect 0 49270 1459 49272
rect 0 49240 800 49270
rect 1393 49267 1459 49270
rect 40493 49330 40559 49333
rect 41200 49330 42000 49360
rect 40493 49328 42000 49330
rect 40493 49272 40498 49328
rect 40554 49272 42000 49328
rect 40493 49270 42000 49272
rect 40493 49267 40559 49270
rect 41200 49240 42000 49270
rect 2606 48992 2922 48993
rect 2606 48928 2612 48992
rect 2676 48928 2692 48992
rect 2756 48928 2772 48992
rect 2836 48928 2852 48992
rect 2916 48928 2922 48992
rect 2606 48927 2922 48928
rect 7606 48992 7922 48993
rect 7606 48928 7612 48992
rect 7676 48928 7692 48992
rect 7756 48928 7772 48992
rect 7836 48928 7852 48992
rect 7916 48928 7922 48992
rect 7606 48927 7922 48928
rect 12606 48992 12922 48993
rect 12606 48928 12612 48992
rect 12676 48928 12692 48992
rect 12756 48928 12772 48992
rect 12836 48928 12852 48992
rect 12916 48928 12922 48992
rect 12606 48927 12922 48928
rect 17606 48992 17922 48993
rect 17606 48928 17612 48992
rect 17676 48928 17692 48992
rect 17756 48928 17772 48992
rect 17836 48928 17852 48992
rect 17916 48928 17922 48992
rect 17606 48927 17922 48928
rect 22606 48992 22922 48993
rect 22606 48928 22612 48992
rect 22676 48928 22692 48992
rect 22756 48928 22772 48992
rect 22836 48928 22852 48992
rect 22916 48928 22922 48992
rect 22606 48927 22922 48928
rect 27606 48992 27922 48993
rect 27606 48928 27612 48992
rect 27676 48928 27692 48992
rect 27756 48928 27772 48992
rect 27836 48928 27852 48992
rect 27916 48928 27922 48992
rect 27606 48927 27922 48928
rect 32606 48992 32922 48993
rect 32606 48928 32612 48992
rect 32676 48928 32692 48992
rect 32756 48928 32772 48992
rect 32836 48928 32852 48992
rect 32916 48928 32922 48992
rect 32606 48927 32922 48928
rect 37606 48992 37922 48993
rect 37606 48928 37612 48992
rect 37676 48928 37692 48992
rect 37756 48928 37772 48992
rect 37836 48928 37852 48992
rect 37916 48928 37922 48992
rect 37606 48927 37922 48928
rect 1946 48448 2262 48449
rect 1946 48384 1952 48448
rect 2016 48384 2032 48448
rect 2096 48384 2112 48448
rect 2176 48384 2192 48448
rect 2256 48384 2262 48448
rect 1946 48383 2262 48384
rect 6946 48448 7262 48449
rect 6946 48384 6952 48448
rect 7016 48384 7032 48448
rect 7096 48384 7112 48448
rect 7176 48384 7192 48448
rect 7256 48384 7262 48448
rect 6946 48383 7262 48384
rect 11946 48448 12262 48449
rect 11946 48384 11952 48448
rect 12016 48384 12032 48448
rect 12096 48384 12112 48448
rect 12176 48384 12192 48448
rect 12256 48384 12262 48448
rect 11946 48383 12262 48384
rect 16946 48448 17262 48449
rect 16946 48384 16952 48448
rect 17016 48384 17032 48448
rect 17096 48384 17112 48448
rect 17176 48384 17192 48448
rect 17256 48384 17262 48448
rect 16946 48383 17262 48384
rect 21946 48448 22262 48449
rect 21946 48384 21952 48448
rect 22016 48384 22032 48448
rect 22096 48384 22112 48448
rect 22176 48384 22192 48448
rect 22256 48384 22262 48448
rect 21946 48383 22262 48384
rect 26946 48448 27262 48449
rect 26946 48384 26952 48448
rect 27016 48384 27032 48448
rect 27096 48384 27112 48448
rect 27176 48384 27192 48448
rect 27256 48384 27262 48448
rect 26946 48383 27262 48384
rect 31946 48448 32262 48449
rect 31946 48384 31952 48448
rect 32016 48384 32032 48448
rect 32096 48384 32112 48448
rect 32176 48384 32192 48448
rect 32256 48384 32262 48448
rect 31946 48383 32262 48384
rect 36946 48448 37262 48449
rect 36946 48384 36952 48448
rect 37016 48384 37032 48448
rect 37096 48384 37112 48448
rect 37176 48384 37192 48448
rect 37256 48384 37262 48448
rect 36946 48383 37262 48384
rect 2606 47904 2922 47905
rect 2606 47840 2612 47904
rect 2676 47840 2692 47904
rect 2756 47840 2772 47904
rect 2836 47840 2852 47904
rect 2916 47840 2922 47904
rect 2606 47839 2922 47840
rect 7606 47904 7922 47905
rect 7606 47840 7612 47904
rect 7676 47840 7692 47904
rect 7756 47840 7772 47904
rect 7836 47840 7852 47904
rect 7916 47840 7922 47904
rect 7606 47839 7922 47840
rect 12606 47904 12922 47905
rect 12606 47840 12612 47904
rect 12676 47840 12692 47904
rect 12756 47840 12772 47904
rect 12836 47840 12852 47904
rect 12916 47840 12922 47904
rect 12606 47839 12922 47840
rect 17606 47904 17922 47905
rect 17606 47840 17612 47904
rect 17676 47840 17692 47904
rect 17756 47840 17772 47904
rect 17836 47840 17852 47904
rect 17916 47840 17922 47904
rect 17606 47839 17922 47840
rect 22606 47904 22922 47905
rect 22606 47840 22612 47904
rect 22676 47840 22692 47904
rect 22756 47840 22772 47904
rect 22836 47840 22852 47904
rect 22916 47840 22922 47904
rect 22606 47839 22922 47840
rect 27606 47904 27922 47905
rect 27606 47840 27612 47904
rect 27676 47840 27692 47904
rect 27756 47840 27772 47904
rect 27836 47840 27852 47904
rect 27916 47840 27922 47904
rect 27606 47839 27922 47840
rect 32606 47904 32922 47905
rect 32606 47840 32612 47904
rect 32676 47840 32692 47904
rect 32756 47840 32772 47904
rect 32836 47840 32852 47904
rect 32916 47840 32922 47904
rect 32606 47839 32922 47840
rect 37606 47904 37922 47905
rect 37606 47840 37612 47904
rect 37676 47840 37692 47904
rect 37756 47840 37772 47904
rect 37836 47840 37852 47904
rect 37916 47840 37922 47904
rect 37606 47839 37922 47840
rect 1946 47360 2262 47361
rect 1946 47296 1952 47360
rect 2016 47296 2032 47360
rect 2096 47296 2112 47360
rect 2176 47296 2192 47360
rect 2256 47296 2262 47360
rect 1946 47295 2262 47296
rect 6946 47360 7262 47361
rect 6946 47296 6952 47360
rect 7016 47296 7032 47360
rect 7096 47296 7112 47360
rect 7176 47296 7192 47360
rect 7256 47296 7262 47360
rect 6946 47295 7262 47296
rect 11946 47360 12262 47361
rect 11946 47296 11952 47360
rect 12016 47296 12032 47360
rect 12096 47296 12112 47360
rect 12176 47296 12192 47360
rect 12256 47296 12262 47360
rect 11946 47295 12262 47296
rect 16946 47360 17262 47361
rect 16946 47296 16952 47360
rect 17016 47296 17032 47360
rect 17096 47296 17112 47360
rect 17176 47296 17192 47360
rect 17256 47296 17262 47360
rect 16946 47295 17262 47296
rect 21946 47360 22262 47361
rect 21946 47296 21952 47360
rect 22016 47296 22032 47360
rect 22096 47296 22112 47360
rect 22176 47296 22192 47360
rect 22256 47296 22262 47360
rect 21946 47295 22262 47296
rect 26946 47360 27262 47361
rect 26946 47296 26952 47360
rect 27016 47296 27032 47360
rect 27096 47296 27112 47360
rect 27176 47296 27192 47360
rect 27256 47296 27262 47360
rect 26946 47295 27262 47296
rect 31946 47360 32262 47361
rect 31946 47296 31952 47360
rect 32016 47296 32032 47360
rect 32096 47296 32112 47360
rect 32176 47296 32192 47360
rect 32256 47296 32262 47360
rect 31946 47295 32262 47296
rect 36946 47360 37262 47361
rect 36946 47296 36952 47360
rect 37016 47296 37032 47360
rect 37096 47296 37112 47360
rect 37176 47296 37192 47360
rect 37256 47296 37262 47360
rect 36946 47295 37262 47296
rect 2606 46816 2922 46817
rect 2606 46752 2612 46816
rect 2676 46752 2692 46816
rect 2756 46752 2772 46816
rect 2836 46752 2852 46816
rect 2916 46752 2922 46816
rect 2606 46751 2922 46752
rect 7606 46816 7922 46817
rect 7606 46752 7612 46816
rect 7676 46752 7692 46816
rect 7756 46752 7772 46816
rect 7836 46752 7852 46816
rect 7916 46752 7922 46816
rect 7606 46751 7922 46752
rect 12606 46816 12922 46817
rect 12606 46752 12612 46816
rect 12676 46752 12692 46816
rect 12756 46752 12772 46816
rect 12836 46752 12852 46816
rect 12916 46752 12922 46816
rect 12606 46751 12922 46752
rect 17606 46816 17922 46817
rect 17606 46752 17612 46816
rect 17676 46752 17692 46816
rect 17756 46752 17772 46816
rect 17836 46752 17852 46816
rect 17916 46752 17922 46816
rect 17606 46751 17922 46752
rect 22606 46816 22922 46817
rect 22606 46752 22612 46816
rect 22676 46752 22692 46816
rect 22756 46752 22772 46816
rect 22836 46752 22852 46816
rect 22916 46752 22922 46816
rect 22606 46751 22922 46752
rect 27606 46816 27922 46817
rect 27606 46752 27612 46816
rect 27676 46752 27692 46816
rect 27756 46752 27772 46816
rect 27836 46752 27852 46816
rect 27916 46752 27922 46816
rect 27606 46751 27922 46752
rect 32606 46816 32922 46817
rect 32606 46752 32612 46816
rect 32676 46752 32692 46816
rect 32756 46752 32772 46816
rect 32836 46752 32852 46816
rect 32916 46752 32922 46816
rect 32606 46751 32922 46752
rect 37606 46816 37922 46817
rect 37606 46752 37612 46816
rect 37676 46752 37692 46816
rect 37756 46752 37772 46816
rect 37836 46752 37852 46816
rect 37916 46752 37922 46816
rect 37606 46751 37922 46752
rect 1946 46272 2262 46273
rect 1946 46208 1952 46272
rect 2016 46208 2032 46272
rect 2096 46208 2112 46272
rect 2176 46208 2192 46272
rect 2256 46208 2262 46272
rect 1946 46207 2262 46208
rect 6946 46272 7262 46273
rect 6946 46208 6952 46272
rect 7016 46208 7032 46272
rect 7096 46208 7112 46272
rect 7176 46208 7192 46272
rect 7256 46208 7262 46272
rect 6946 46207 7262 46208
rect 11946 46272 12262 46273
rect 11946 46208 11952 46272
rect 12016 46208 12032 46272
rect 12096 46208 12112 46272
rect 12176 46208 12192 46272
rect 12256 46208 12262 46272
rect 11946 46207 12262 46208
rect 16946 46272 17262 46273
rect 16946 46208 16952 46272
rect 17016 46208 17032 46272
rect 17096 46208 17112 46272
rect 17176 46208 17192 46272
rect 17256 46208 17262 46272
rect 16946 46207 17262 46208
rect 21946 46272 22262 46273
rect 21946 46208 21952 46272
rect 22016 46208 22032 46272
rect 22096 46208 22112 46272
rect 22176 46208 22192 46272
rect 22256 46208 22262 46272
rect 21946 46207 22262 46208
rect 26946 46272 27262 46273
rect 26946 46208 26952 46272
rect 27016 46208 27032 46272
rect 27096 46208 27112 46272
rect 27176 46208 27192 46272
rect 27256 46208 27262 46272
rect 26946 46207 27262 46208
rect 31946 46272 32262 46273
rect 31946 46208 31952 46272
rect 32016 46208 32032 46272
rect 32096 46208 32112 46272
rect 32176 46208 32192 46272
rect 32256 46208 32262 46272
rect 31946 46207 32262 46208
rect 36946 46272 37262 46273
rect 36946 46208 36952 46272
rect 37016 46208 37032 46272
rect 37096 46208 37112 46272
rect 37176 46208 37192 46272
rect 37256 46208 37262 46272
rect 36946 46207 37262 46208
rect 2606 45728 2922 45729
rect 2606 45664 2612 45728
rect 2676 45664 2692 45728
rect 2756 45664 2772 45728
rect 2836 45664 2852 45728
rect 2916 45664 2922 45728
rect 2606 45663 2922 45664
rect 7606 45728 7922 45729
rect 7606 45664 7612 45728
rect 7676 45664 7692 45728
rect 7756 45664 7772 45728
rect 7836 45664 7852 45728
rect 7916 45664 7922 45728
rect 7606 45663 7922 45664
rect 12606 45728 12922 45729
rect 12606 45664 12612 45728
rect 12676 45664 12692 45728
rect 12756 45664 12772 45728
rect 12836 45664 12852 45728
rect 12916 45664 12922 45728
rect 12606 45663 12922 45664
rect 17606 45728 17922 45729
rect 17606 45664 17612 45728
rect 17676 45664 17692 45728
rect 17756 45664 17772 45728
rect 17836 45664 17852 45728
rect 17916 45664 17922 45728
rect 17606 45663 17922 45664
rect 22606 45728 22922 45729
rect 22606 45664 22612 45728
rect 22676 45664 22692 45728
rect 22756 45664 22772 45728
rect 22836 45664 22852 45728
rect 22916 45664 22922 45728
rect 22606 45663 22922 45664
rect 27606 45728 27922 45729
rect 27606 45664 27612 45728
rect 27676 45664 27692 45728
rect 27756 45664 27772 45728
rect 27836 45664 27852 45728
rect 27916 45664 27922 45728
rect 27606 45663 27922 45664
rect 32606 45728 32922 45729
rect 32606 45664 32612 45728
rect 32676 45664 32692 45728
rect 32756 45664 32772 45728
rect 32836 45664 32852 45728
rect 32916 45664 32922 45728
rect 32606 45663 32922 45664
rect 37606 45728 37922 45729
rect 37606 45664 37612 45728
rect 37676 45664 37692 45728
rect 37756 45664 37772 45728
rect 37836 45664 37852 45728
rect 37916 45664 37922 45728
rect 37606 45663 37922 45664
rect 1946 45184 2262 45185
rect 1946 45120 1952 45184
rect 2016 45120 2032 45184
rect 2096 45120 2112 45184
rect 2176 45120 2192 45184
rect 2256 45120 2262 45184
rect 1946 45119 2262 45120
rect 6946 45184 7262 45185
rect 6946 45120 6952 45184
rect 7016 45120 7032 45184
rect 7096 45120 7112 45184
rect 7176 45120 7192 45184
rect 7256 45120 7262 45184
rect 6946 45119 7262 45120
rect 11946 45184 12262 45185
rect 11946 45120 11952 45184
rect 12016 45120 12032 45184
rect 12096 45120 12112 45184
rect 12176 45120 12192 45184
rect 12256 45120 12262 45184
rect 11946 45119 12262 45120
rect 16946 45184 17262 45185
rect 16946 45120 16952 45184
rect 17016 45120 17032 45184
rect 17096 45120 17112 45184
rect 17176 45120 17192 45184
rect 17256 45120 17262 45184
rect 16946 45119 17262 45120
rect 21946 45184 22262 45185
rect 21946 45120 21952 45184
rect 22016 45120 22032 45184
rect 22096 45120 22112 45184
rect 22176 45120 22192 45184
rect 22256 45120 22262 45184
rect 21946 45119 22262 45120
rect 26946 45184 27262 45185
rect 26946 45120 26952 45184
rect 27016 45120 27032 45184
rect 27096 45120 27112 45184
rect 27176 45120 27192 45184
rect 27256 45120 27262 45184
rect 26946 45119 27262 45120
rect 31946 45184 32262 45185
rect 31946 45120 31952 45184
rect 32016 45120 32032 45184
rect 32096 45120 32112 45184
rect 32176 45120 32192 45184
rect 32256 45120 32262 45184
rect 31946 45119 32262 45120
rect 36946 45184 37262 45185
rect 36946 45120 36952 45184
rect 37016 45120 37032 45184
rect 37096 45120 37112 45184
rect 37176 45120 37192 45184
rect 37256 45120 37262 45184
rect 36946 45119 37262 45120
rect 2606 44640 2922 44641
rect 2606 44576 2612 44640
rect 2676 44576 2692 44640
rect 2756 44576 2772 44640
rect 2836 44576 2852 44640
rect 2916 44576 2922 44640
rect 2606 44575 2922 44576
rect 7606 44640 7922 44641
rect 7606 44576 7612 44640
rect 7676 44576 7692 44640
rect 7756 44576 7772 44640
rect 7836 44576 7852 44640
rect 7916 44576 7922 44640
rect 7606 44575 7922 44576
rect 12606 44640 12922 44641
rect 12606 44576 12612 44640
rect 12676 44576 12692 44640
rect 12756 44576 12772 44640
rect 12836 44576 12852 44640
rect 12916 44576 12922 44640
rect 12606 44575 12922 44576
rect 17606 44640 17922 44641
rect 17606 44576 17612 44640
rect 17676 44576 17692 44640
rect 17756 44576 17772 44640
rect 17836 44576 17852 44640
rect 17916 44576 17922 44640
rect 17606 44575 17922 44576
rect 22606 44640 22922 44641
rect 22606 44576 22612 44640
rect 22676 44576 22692 44640
rect 22756 44576 22772 44640
rect 22836 44576 22852 44640
rect 22916 44576 22922 44640
rect 22606 44575 22922 44576
rect 27606 44640 27922 44641
rect 27606 44576 27612 44640
rect 27676 44576 27692 44640
rect 27756 44576 27772 44640
rect 27836 44576 27852 44640
rect 27916 44576 27922 44640
rect 27606 44575 27922 44576
rect 32606 44640 32922 44641
rect 32606 44576 32612 44640
rect 32676 44576 32692 44640
rect 32756 44576 32772 44640
rect 32836 44576 32852 44640
rect 32916 44576 32922 44640
rect 32606 44575 32922 44576
rect 37606 44640 37922 44641
rect 37606 44576 37612 44640
rect 37676 44576 37692 44640
rect 37756 44576 37772 44640
rect 37836 44576 37852 44640
rect 37916 44576 37922 44640
rect 37606 44575 37922 44576
rect 1946 44096 2262 44097
rect 1946 44032 1952 44096
rect 2016 44032 2032 44096
rect 2096 44032 2112 44096
rect 2176 44032 2192 44096
rect 2256 44032 2262 44096
rect 1946 44031 2262 44032
rect 6946 44096 7262 44097
rect 6946 44032 6952 44096
rect 7016 44032 7032 44096
rect 7096 44032 7112 44096
rect 7176 44032 7192 44096
rect 7256 44032 7262 44096
rect 6946 44031 7262 44032
rect 11946 44096 12262 44097
rect 11946 44032 11952 44096
rect 12016 44032 12032 44096
rect 12096 44032 12112 44096
rect 12176 44032 12192 44096
rect 12256 44032 12262 44096
rect 11946 44031 12262 44032
rect 16946 44096 17262 44097
rect 16946 44032 16952 44096
rect 17016 44032 17032 44096
rect 17096 44032 17112 44096
rect 17176 44032 17192 44096
rect 17256 44032 17262 44096
rect 16946 44031 17262 44032
rect 21946 44096 22262 44097
rect 21946 44032 21952 44096
rect 22016 44032 22032 44096
rect 22096 44032 22112 44096
rect 22176 44032 22192 44096
rect 22256 44032 22262 44096
rect 21946 44031 22262 44032
rect 26946 44096 27262 44097
rect 26946 44032 26952 44096
rect 27016 44032 27032 44096
rect 27096 44032 27112 44096
rect 27176 44032 27192 44096
rect 27256 44032 27262 44096
rect 26946 44031 27262 44032
rect 31946 44096 32262 44097
rect 31946 44032 31952 44096
rect 32016 44032 32032 44096
rect 32096 44032 32112 44096
rect 32176 44032 32192 44096
rect 32256 44032 32262 44096
rect 31946 44031 32262 44032
rect 36946 44096 37262 44097
rect 36946 44032 36952 44096
rect 37016 44032 37032 44096
rect 37096 44032 37112 44096
rect 37176 44032 37192 44096
rect 37256 44032 37262 44096
rect 36946 44031 37262 44032
rect 2606 43552 2922 43553
rect 2606 43488 2612 43552
rect 2676 43488 2692 43552
rect 2756 43488 2772 43552
rect 2836 43488 2852 43552
rect 2916 43488 2922 43552
rect 2606 43487 2922 43488
rect 7606 43552 7922 43553
rect 7606 43488 7612 43552
rect 7676 43488 7692 43552
rect 7756 43488 7772 43552
rect 7836 43488 7852 43552
rect 7916 43488 7922 43552
rect 7606 43487 7922 43488
rect 12606 43552 12922 43553
rect 12606 43488 12612 43552
rect 12676 43488 12692 43552
rect 12756 43488 12772 43552
rect 12836 43488 12852 43552
rect 12916 43488 12922 43552
rect 12606 43487 12922 43488
rect 17606 43552 17922 43553
rect 17606 43488 17612 43552
rect 17676 43488 17692 43552
rect 17756 43488 17772 43552
rect 17836 43488 17852 43552
rect 17916 43488 17922 43552
rect 17606 43487 17922 43488
rect 22606 43552 22922 43553
rect 22606 43488 22612 43552
rect 22676 43488 22692 43552
rect 22756 43488 22772 43552
rect 22836 43488 22852 43552
rect 22916 43488 22922 43552
rect 22606 43487 22922 43488
rect 27606 43552 27922 43553
rect 27606 43488 27612 43552
rect 27676 43488 27692 43552
rect 27756 43488 27772 43552
rect 27836 43488 27852 43552
rect 27916 43488 27922 43552
rect 27606 43487 27922 43488
rect 32606 43552 32922 43553
rect 32606 43488 32612 43552
rect 32676 43488 32692 43552
rect 32756 43488 32772 43552
rect 32836 43488 32852 43552
rect 32916 43488 32922 43552
rect 32606 43487 32922 43488
rect 37606 43552 37922 43553
rect 37606 43488 37612 43552
rect 37676 43488 37692 43552
rect 37756 43488 37772 43552
rect 37836 43488 37852 43552
rect 37916 43488 37922 43552
rect 37606 43487 37922 43488
rect 1946 43008 2262 43009
rect 1946 42944 1952 43008
rect 2016 42944 2032 43008
rect 2096 42944 2112 43008
rect 2176 42944 2192 43008
rect 2256 42944 2262 43008
rect 1946 42943 2262 42944
rect 6946 43008 7262 43009
rect 6946 42944 6952 43008
rect 7016 42944 7032 43008
rect 7096 42944 7112 43008
rect 7176 42944 7192 43008
rect 7256 42944 7262 43008
rect 6946 42943 7262 42944
rect 11946 43008 12262 43009
rect 11946 42944 11952 43008
rect 12016 42944 12032 43008
rect 12096 42944 12112 43008
rect 12176 42944 12192 43008
rect 12256 42944 12262 43008
rect 11946 42943 12262 42944
rect 16946 43008 17262 43009
rect 16946 42944 16952 43008
rect 17016 42944 17032 43008
rect 17096 42944 17112 43008
rect 17176 42944 17192 43008
rect 17256 42944 17262 43008
rect 16946 42943 17262 42944
rect 21946 43008 22262 43009
rect 21946 42944 21952 43008
rect 22016 42944 22032 43008
rect 22096 42944 22112 43008
rect 22176 42944 22192 43008
rect 22256 42944 22262 43008
rect 21946 42943 22262 42944
rect 26946 43008 27262 43009
rect 26946 42944 26952 43008
rect 27016 42944 27032 43008
rect 27096 42944 27112 43008
rect 27176 42944 27192 43008
rect 27256 42944 27262 43008
rect 26946 42943 27262 42944
rect 31946 43008 32262 43009
rect 31946 42944 31952 43008
rect 32016 42944 32032 43008
rect 32096 42944 32112 43008
rect 32176 42944 32192 43008
rect 32256 42944 32262 43008
rect 31946 42943 32262 42944
rect 36946 43008 37262 43009
rect 36946 42944 36952 43008
rect 37016 42944 37032 43008
rect 37096 42944 37112 43008
rect 37176 42944 37192 43008
rect 37256 42944 37262 43008
rect 36946 42943 37262 42944
rect 22093 42802 22159 42805
rect 22461 42802 22527 42805
rect 22093 42800 22527 42802
rect 22093 42744 22098 42800
rect 22154 42744 22466 42800
rect 22522 42744 22527 42800
rect 22093 42742 22527 42744
rect 22093 42739 22159 42742
rect 22461 42739 22527 42742
rect 2606 42464 2922 42465
rect 2606 42400 2612 42464
rect 2676 42400 2692 42464
rect 2756 42400 2772 42464
rect 2836 42400 2852 42464
rect 2916 42400 2922 42464
rect 2606 42399 2922 42400
rect 7606 42464 7922 42465
rect 7606 42400 7612 42464
rect 7676 42400 7692 42464
rect 7756 42400 7772 42464
rect 7836 42400 7852 42464
rect 7916 42400 7922 42464
rect 7606 42399 7922 42400
rect 12606 42464 12922 42465
rect 12606 42400 12612 42464
rect 12676 42400 12692 42464
rect 12756 42400 12772 42464
rect 12836 42400 12852 42464
rect 12916 42400 12922 42464
rect 12606 42399 12922 42400
rect 17606 42464 17922 42465
rect 17606 42400 17612 42464
rect 17676 42400 17692 42464
rect 17756 42400 17772 42464
rect 17836 42400 17852 42464
rect 17916 42400 17922 42464
rect 17606 42399 17922 42400
rect 22606 42464 22922 42465
rect 22606 42400 22612 42464
rect 22676 42400 22692 42464
rect 22756 42400 22772 42464
rect 22836 42400 22852 42464
rect 22916 42400 22922 42464
rect 22606 42399 22922 42400
rect 27606 42464 27922 42465
rect 27606 42400 27612 42464
rect 27676 42400 27692 42464
rect 27756 42400 27772 42464
rect 27836 42400 27852 42464
rect 27916 42400 27922 42464
rect 27606 42399 27922 42400
rect 32606 42464 32922 42465
rect 32606 42400 32612 42464
rect 32676 42400 32692 42464
rect 32756 42400 32772 42464
rect 32836 42400 32852 42464
rect 32916 42400 32922 42464
rect 32606 42399 32922 42400
rect 37606 42464 37922 42465
rect 37606 42400 37612 42464
rect 37676 42400 37692 42464
rect 37756 42400 37772 42464
rect 37836 42400 37852 42464
rect 37916 42400 37922 42464
rect 37606 42399 37922 42400
rect 1946 41920 2262 41921
rect 1946 41856 1952 41920
rect 2016 41856 2032 41920
rect 2096 41856 2112 41920
rect 2176 41856 2192 41920
rect 2256 41856 2262 41920
rect 1946 41855 2262 41856
rect 6946 41920 7262 41921
rect 6946 41856 6952 41920
rect 7016 41856 7032 41920
rect 7096 41856 7112 41920
rect 7176 41856 7192 41920
rect 7256 41856 7262 41920
rect 6946 41855 7262 41856
rect 11946 41920 12262 41921
rect 11946 41856 11952 41920
rect 12016 41856 12032 41920
rect 12096 41856 12112 41920
rect 12176 41856 12192 41920
rect 12256 41856 12262 41920
rect 11946 41855 12262 41856
rect 16946 41920 17262 41921
rect 16946 41856 16952 41920
rect 17016 41856 17032 41920
rect 17096 41856 17112 41920
rect 17176 41856 17192 41920
rect 17256 41856 17262 41920
rect 16946 41855 17262 41856
rect 21946 41920 22262 41921
rect 21946 41856 21952 41920
rect 22016 41856 22032 41920
rect 22096 41856 22112 41920
rect 22176 41856 22192 41920
rect 22256 41856 22262 41920
rect 21946 41855 22262 41856
rect 26946 41920 27262 41921
rect 26946 41856 26952 41920
rect 27016 41856 27032 41920
rect 27096 41856 27112 41920
rect 27176 41856 27192 41920
rect 27256 41856 27262 41920
rect 26946 41855 27262 41856
rect 31946 41920 32262 41921
rect 31946 41856 31952 41920
rect 32016 41856 32032 41920
rect 32096 41856 32112 41920
rect 32176 41856 32192 41920
rect 32256 41856 32262 41920
rect 31946 41855 32262 41856
rect 36946 41920 37262 41921
rect 36946 41856 36952 41920
rect 37016 41856 37032 41920
rect 37096 41856 37112 41920
rect 37176 41856 37192 41920
rect 37256 41856 37262 41920
rect 36946 41855 37262 41856
rect 2606 41376 2922 41377
rect 2606 41312 2612 41376
rect 2676 41312 2692 41376
rect 2756 41312 2772 41376
rect 2836 41312 2852 41376
rect 2916 41312 2922 41376
rect 2606 41311 2922 41312
rect 7606 41376 7922 41377
rect 7606 41312 7612 41376
rect 7676 41312 7692 41376
rect 7756 41312 7772 41376
rect 7836 41312 7852 41376
rect 7916 41312 7922 41376
rect 7606 41311 7922 41312
rect 12606 41376 12922 41377
rect 12606 41312 12612 41376
rect 12676 41312 12692 41376
rect 12756 41312 12772 41376
rect 12836 41312 12852 41376
rect 12916 41312 12922 41376
rect 12606 41311 12922 41312
rect 17606 41376 17922 41377
rect 17606 41312 17612 41376
rect 17676 41312 17692 41376
rect 17756 41312 17772 41376
rect 17836 41312 17852 41376
rect 17916 41312 17922 41376
rect 17606 41311 17922 41312
rect 22606 41376 22922 41377
rect 22606 41312 22612 41376
rect 22676 41312 22692 41376
rect 22756 41312 22772 41376
rect 22836 41312 22852 41376
rect 22916 41312 22922 41376
rect 22606 41311 22922 41312
rect 27606 41376 27922 41377
rect 27606 41312 27612 41376
rect 27676 41312 27692 41376
rect 27756 41312 27772 41376
rect 27836 41312 27852 41376
rect 27916 41312 27922 41376
rect 27606 41311 27922 41312
rect 32606 41376 32922 41377
rect 32606 41312 32612 41376
rect 32676 41312 32692 41376
rect 32756 41312 32772 41376
rect 32836 41312 32852 41376
rect 32916 41312 32922 41376
rect 32606 41311 32922 41312
rect 37606 41376 37922 41377
rect 37606 41312 37612 41376
rect 37676 41312 37692 41376
rect 37756 41312 37772 41376
rect 37836 41312 37852 41376
rect 37916 41312 37922 41376
rect 37606 41311 37922 41312
rect 1946 40832 2262 40833
rect 1946 40768 1952 40832
rect 2016 40768 2032 40832
rect 2096 40768 2112 40832
rect 2176 40768 2192 40832
rect 2256 40768 2262 40832
rect 1946 40767 2262 40768
rect 6946 40832 7262 40833
rect 6946 40768 6952 40832
rect 7016 40768 7032 40832
rect 7096 40768 7112 40832
rect 7176 40768 7192 40832
rect 7256 40768 7262 40832
rect 6946 40767 7262 40768
rect 11946 40832 12262 40833
rect 11946 40768 11952 40832
rect 12016 40768 12032 40832
rect 12096 40768 12112 40832
rect 12176 40768 12192 40832
rect 12256 40768 12262 40832
rect 11946 40767 12262 40768
rect 16946 40832 17262 40833
rect 16946 40768 16952 40832
rect 17016 40768 17032 40832
rect 17096 40768 17112 40832
rect 17176 40768 17192 40832
rect 17256 40768 17262 40832
rect 16946 40767 17262 40768
rect 21946 40832 22262 40833
rect 21946 40768 21952 40832
rect 22016 40768 22032 40832
rect 22096 40768 22112 40832
rect 22176 40768 22192 40832
rect 22256 40768 22262 40832
rect 21946 40767 22262 40768
rect 26946 40832 27262 40833
rect 26946 40768 26952 40832
rect 27016 40768 27032 40832
rect 27096 40768 27112 40832
rect 27176 40768 27192 40832
rect 27256 40768 27262 40832
rect 26946 40767 27262 40768
rect 31946 40832 32262 40833
rect 31946 40768 31952 40832
rect 32016 40768 32032 40832
rect 32096 40768 32112 40832
rect 32176 40768 32192 40832
rect 32256 40768 32262 40832
rect 31946 40767 32262 40768
rect 36946 40832 37262 40833
rect 36946 40768 36952 40832
rect 37016 40768 37032 40832
rect 37096 40768 37112 40832
rect 37176 40768 37192 40832
rect 37256 40768 37262 40832
rect 36946 40767 37262 40768
rect 23565 40628 23631 40629
rect 23565 40624 23612 40628
rect 23676 40626 23682 40628
rect 23565 40568 23570 40624
rect 23565 40564 23612 40568
rect 23676 40566 23722 40626
rect 23676 40564 23682 40566
rect 23565 40563 23631 40564
rect 0 40354 800 40384
rect 40861 40354 40927 40357
rect 41200 40354 42000 40384
rect 0 40264 858 40354
rect 40861 40352 42000 40354
rect 40861 40296 40866 40352
rect 40922 40296 42000 40352
rect 40861 40294 42000 40296
rect 40861 40291 40927 40294
rect 798 40221 858 40264
rect 2606 40288 2922 40289
rect 2606 40224 2612 40288
rect 2676 40224 2692 40288
rect 2756 40224 2772 40288
rect 2836 40224 2852 40288
rect 2916 40224 2922 40288
rect 2606 40223 2922 40224
rect 7606 40288 7922 40289
rect 7606 40224 7612 40288
rect 7676 40224 7692 40288
rect 7756 40224 7772 40288
rect 7836 40224 7852 40288
rect 7916 40224 7922 40288
rect 7606 40223 7922 40224
rect 12606 40288 12922 40289
rect 12606 40224 12612 40288
rect 12676 40224 12692 40288
rect 12756 40224 12772 40288
rect 12836 40224 12852 40288
rect 12916 40224 12922 40288
rect 12606 40223 12922 40224
rect 17606 40288 17922 40289
rect 17606 40224 17612 40288
rect 17676 40224 17692 40288
rect 17756 40224 17772 40288
rect 17836 40224 17852 40288
rect 17916 40224 17922 40288
rect 17606 40223 17922 40224
rect 22606 40288 22922 40289
rect 22606 40224 22612 40288
rect 22676 40224 22692 40288
rect 22756 40224 22772 40288
rect 22836 40224 22852 40288
rect 22916 40224 22922 40288
rect 22606 40223 22922 40224
rect 27606 40288 27922 40289
rect 27606 40224 27612 40288
rect 27676 40224 27692 40288
rect 27756 40224 27772 40288
rect 27836 40224 27852 40288
rect 27916 40224 27922 40288
rect 27606 40223 27922 40224
rect 32606 40288 32922 40289
rect 32606 40224 32612 40288
rect 32676 40224 32692 40288
rect 32756 40224 32772 40288
rect 32836 40224 32852 40288
rect 32916 40224 32922 40288
rect 32606 40223 32922 40224
rect 37606 40288 37922 40289
rect 37606 40224 37612 40288
rect 37676 40224 37692 40288
rect 37756 40224 37772 40288
rect 37836 40224 37852 40288
rect 37916 40224 37922 40288
rect 41200 40264 42000 40294
rect 37606 40223 37922 40224
rect 798 40216 907 40221
rect 798 40160 846 40216
rect 902 40160 907 40216
rect 798 40158 907 40160
rect 841 40155 907 40158
rect 30557 40084 30623 40085
rect 30557 40082 30604 40084
rect 30512 40080 30604 40082
rect 30512 40024 30562 40080
rect 30512 40022 30604 40024
rect 30557 40020 30604 40022
rect 30668 40020 30674 40084
rect 30557 40019 30623 40020
rect 1946 39744 2262 39745
rect 1946 39680 1952 39744
rect 2016 39680 2032 39744
rect 2096 39680 2112 39744
rect 2176 39680 2192 39744
rect 2256 39680 2262 39744
rect 1946 39679 2262 39680
rect 6946 39744 7262 39745
rect 6946 39680 6952 39744
rect 7016 39680 7032 39744
rect 7096 39680 7112 39744
rect 7176 39680 7192 39744
rect 7256 39680 7262 39744
rect 6946 39679 7262 39680
rect 11946 39744 12262 39745
rect 11946 39680 11952 39744
rect 12016 39680 12032 39744
rect 12096 39680 12112 39744
rect 12176 39680 12192 39744
rect 12256 39680 12262 39744
rect 11946 39679 12262 39680
rect 16946 39744 17262 39745
rect 16946 39680 16952 39744
rect 17016 39680 17032 39744
rect 17096 39680 17112 39744
rect 17176 39680 17192 39744
rect 17256 39680 17262 39744
rect 16946 39679 17262 39680
rect 21946 39744 22262 39745
rect 21946 39680 21952 39744
rect 22016 39680 22032 39744
rect 22096 39680 22112 39744
rect 22176 39680 22192 39744
rect 22256 39680 22262 39744
rect 21946 39679 22262 39680
rect 26946 39744 27262 39745
rect 26946 39680 26952 39744
rect 27016 39680 27032 39744
rect 27096 39680 27112 39744
rect 27176 39680 27192 39744
rect 27256 39680 27262 39744
rect 26946 39679 27262 39680
rect 31946 39744 32262 39745
rect 31946 39680 31952 39744
rect 32016 39680 32032 39744
rect 32096 39680 32112 39744
rect 32176 39680 32192 39744
rect 32256 39680 32262 39744
rect 31946 39679 32262 39680
rect 36946 39744 37262 39745
rect 36946 39680 36952 39744
rect 37016 39680 37032 39744
rect 37096 39680 37112 39744
rect 37176 39680 37192 39744
rect 37256 39680 37262 39744
rect 36946 39679 37262 39680
rect 22185 39402 22251 39405
rect 23841 39402 23907 39405
rect 22185 39400 23907 39402
rect 22185 39344 22190 39400
rect 22246 39344 23846 39400
rect 23902 39344 23907 39400
rect 22185 39342 23907 39344
rect 22185 39339 22251 39342
rect 23841 39339 23907 39342
rect 2606 39200 2922 39201
rect 2606 39136 2612 39200
rect 2676 39136 2692 39200
rect 2756 39136 2772 39200
rect 2836 39136 2852 39200
rect 2916 39136 2922 39200
rect 2606 39135 2922 39136
rect 7606 39200 7922 39201
rect 7606 39136 7612 39200
rect 7676 39136 7692 39200
rect 7756 39136 7772 39200
rect 7836 39136 7852 39200
rect 7916 39136 7922 39200
rect 7606 39135 7922 39136
rect 12606 39200 12922 39201
rect 12606 39136 12612 39200
rect 12676 39136 12692 39200
rect 12756 39136 12772 39200
rect 12836 39136 12852 39200
rect 12916 39136 12922 39200
rect 12606 39135 12922 39136
rect 17606 39200 17922 39201
rect 17606 39136 17612 39200
rect 17676 39136 17692 39200
rect 17756 39136 17772 39200
rect 17836 39136 17852 39200
rect 17916 39136 17922 39200
rect 17606 39135 17922 39136
rect 22606 39200 22922 39201
rect 22606 39136 22612 39200
rect 22676 39136 22692 39200
rect 22756 39136 22772 39200
rect 22836 39136 22852 39200
rect 22916 39136 22922 39200
rect 22606 39135 22922 39136
rect 27606 39200 27922 39201
rect 27606 39136 27612 39200
rect 27676 39136 27692 39200
rect 27756 39136 27772 39200
rect 27836 39136 27852 39200
rect 27916 39136 27922 39200
rect 27606 39135 27922 39136
rect 32606 39200 32922 39201
rect 32606 39136 32612 39200
rect 32676 39136 32692 39200
rect 32756 39136 32772 39200
rect 32836 39136 32852 39200
rect 32916 39136 32922 39200
rect 32606 39135 32922 39136
rect 37606 39200 37922 39201
rect 37606 39136 37612 39200
rect 37676 39136 37692 39200
rect 37756 39136 37772 39200
rect 37836 39136 37852 39200
rect 37916 39136 37922 39200
rect 37606 39135 37922 39136
rect 20161 38994 20227 38997
rect 24577 38994 24643 38997
rect 20161 38992 24643 38994
rect 20161 38936 20166 38992
rect 20222 38936 24582 38992
rect 24638 38936 24643 38992
rect 20161 38934 24643 38936
rect 20161 38931 20227 38934
rect 24577 38931 24643 38934
rect 29085 38994 29151 38997
rect 29361 38994 29427 38997
rect 29085 38992 29427 38994
rect 29085 38936 29090 38992
rect 29146 38936 29366 38992
rect 29422 38936 29427 38992
rect 29085 38934 29427 38936
rect 29085 38931 29151 38934
rect 29361 38931 29427 38934
rect 20345 38858 20411 38861
rect 24301 38858 24367 38861
rect 20345 38856 24367 38858
rect 20345 38800 20350 38856
rect 20406 38800 24306 38856
rect 24362 38800 24367 38856
rect 20345 38798 24367 38800
rect 20345 38795 20411 38798
rect 24301 38795 24367 38798
rect 23238 38660 23244 38724
rect 23308 38722 23314 38724
rect 23381 38722 23447 38725
rect 23308 38720 23447 38722
rect 23308 38664 23386 38720
rect 23442 38664 23447 38720
rect 23308 38662 23447 38664
rect 23308 38660 23314 38662
rect 23381 38659 23447 38662
rect 28993 38722 29059 38725
rect 29545 38722 29611 38725
rect 28993 38720 29611 38722
rect 28993 38664 28998 38720
rect 29054 38664 29550 38720
rect 29606 38664 29611 38720
rect 28993 38662 29611 38664
rect 28993 38659 29059 38662
rect 29545 38659 29611 38662
rect 1946 38656 2262 38657
rect 1946 38592 1952 38656
rect 2016 38592 2032 38656
rect 2096 38592 2112 38656
rect 2176 38592 2192 38656
rect 2256 38592 2262 38656
rect 1946 38591 2262 38592
rect 6946 38656 7262 38657
rect 6946 38592 6952 38656
rect 7016 38592 7032 38656
rect 7096 38592 7112 38656
rect 7176 38592 7192 38656
rect 7256 38592 7262 38656
rect 6946 38591 7262 38592
rect 11946 38656 12262 38657
rect 11946 38592 11952 38656
rect 12016 38592 12032 38656
rect 12096 38592 12112 38656
rect 12176 38592 12192 38656
rect 12256 38592 12262 38656
rect 11946 38591 12262 38592
rect 16946 38656 17262 38657
rect 16946 38592 16952 38656
rect 17016 38592 17032 38656
rect 17096 38592 17112 38656
rect 17176 38592 17192 38656
rect 17256 38592 17262 38656
rect 16946 38591 17262 38592
rect 21946 38656 22262 38657
rect 21946 38592 21952 38656
rect 22016 38592 22032 38656
rect 22096 38592 22112 38656
rect 22176 38592 22192 38656
rect 22256 38592 22262 38656
rect 21946 38591 22262 38592
rect 26946 38656 27262 38657
rect 26946 38592 26952 38656
rect 27016 38592 27032 38656
rect 27096 38592 27112 38656
rect 27176 38592 27192 38656
rect 27256 38592 27262 38656
rect 26946 38591 27262 38592
rect 31946 38656 32262 38657
rect 31946 38592 31952 38656
rect 32016 38592 32032 38656
rect 32096 38592 32112 38656
rect 32176 38592 32192 38656
rect 32256 38592 32262 38656
rect 31946 38591 32262 38592
rect 36946 38656 37262 38657
rect 36946 38592 36952 38656
rect 37016 38592 37032 38656
rect 37096 38592 37112 38656
rect 37176 38592 37192 38656
rect 37256 38592 37262 38656
rect 36946 38591 37262 38592
rect 24761 38452 24827 38453
rect 24710 38450 24716 38452
rect 24670 38390 24716 38450
rect 24780 38448 24827 38452
rect 24822 38392 24827 38448
rect 24710 38388 24716 38390
rect 24780 38388 24827 38392
rect 24761 38387 24827 38388
rect 2606 38112 2922 38113
rect 2606 38048 2612 38112
rect 2676 38048 2692 38112
rect 2756 38048 2772 38112
rect 2836 38048 2852 38112
rect 2916 38048 2922 38112
rect 2606 38047 2922 38048
rect 7606 38112 7922 38113
rect 7606 38048 7612 38112
rect 7676 38048 7692 38112
rect 7756 38048 7772 38112
rect 7836 38048 7852 38112
rect 7916 38048 7922 38112
rect 7606 38047 7922 38048
rect 12606 38112 12922 38113
rect 12606 38048 12612 38112
rect 12676 38048 12692 38112
rect 12756 38048 12772 38112
rect 12836 38048 12852 38112
rect 12916 38048 12922 38112
rect 12606 38047 12922 38048
rect 17606 38112 17922 38113
rect 17606 38048 17612 38112
rect 17676 38048 17692 38112
rect 17756 38048 17772 38112
rect 17836 38048 17852 38112
rect 17916 38048 17922 38112
rect 17606 38047 17922 38048
rect 22606 38112 22922 38113
rect 22606 38048 22612 38112
rect 22676 38048 22692 38112
rect 22756 38048 22772 38112
rect 22836 38048 22852 38112
rect 22916 38048 22922 38112
rect 22606 38047 22922 38048
rect 27606 38112 27922 38113
rect 27606 38048 27612 38112
rect 27676 38048 27692 38112
rect 27756 38048 27772 38112
rect 27836 38048 27852 38112
rect 27916 38048 27922 38112
rect 27606 38047 27922 38048
rect 32606 38112 32922 38113
rect 32606 38048 32612 38112
rect 32676 38048 32692 38112
rect 32756 38048 32772 38112
rect 32836 38048 32852 38112
rect 32916 38048 32922 38112
rect 32606 38047 32922 38048
rect 37606 38112 37922 38113
rect 37606 38048 37612 38112
rect 37676 38048 37692 38112
rect 37756 38048 37772 38112
rect 37836 38048 37852 38112
rect 37916 38048 37922 38112
rect 37606 38047 37922 38048
rect 25221 38044 25287 38045
rect 25221 38042 25268 38044
rect 25176 38040 25268 38042
rect 25176 37984 25226 38040
rect 25176 37982 25268 37984
rect 25221 37980 25268 37982
rect 25332 37980 25338 38044
rect 25221 37979 25287 37980
rect 1946 37568 2262 37569
rect 1946 37504 1952 37568
rect 2016 37504 2032 37568
rect 2096 37504 2112 37568
rect 2176 37504 2192 37568
rect 2256 37504 2262 37568
rect 1946 37503 2262 37504
rect 6946 37568 7262 37569
rect 6946 37504 6952 37568
rect 7016 37504 7032 37568
rect 7096 37504 7112 37568
rect 7176 37504 7192 37568
rect 7256 37504 7262 37568
rect 6946 37503 7262 37504
rect 11946 37568 12262 37569
rect 11946 37504 11952 37568
rect 12016 37504 12032 37568
rect 12096 37504 12112 37568
rect 12176 37504 12192 37568
rect 12256 37504 12262 37568
rect 11946 37503 12262 37504
rect 16946 37568 17262 37569
rect 16946 37504 16952 37568
rect 17016 37504 17032 37568
rect 17096 37504 17112 37568
rect 17176 37504 17192 37568
rect 17256 37504 17262 37568
rect 16946 37503 17262 37504
rect 21946 37568 22262 37569
rect 21946 37504 21952 37568
rect 22016 37504 22032 37568
rect 22096 37504 22112 37568
rect 22176 37504 22192 37568
rect 22256 37504 22262 37568
rect 21946 37503 22262 37504
rect 26946 37568 27262 37569
rect 26946 37504 26952 37568
rect 27016 37504 27032 37568
rect 27096 37504 27112 37568
rect 27176 37504 27192 37568
rect 27256 37504 27262 37568
rect 26946 37503 27262 37504
rect 31946 37568 32262 37569
rect 31946 37504 31952 37568
rect 32016 37504 32032 37568
rect 32096 37504 32112 37568
rect 32176 37504 32192 37568
rect 32256 37504 32262 37568
rect 31946 37503 32262 37504
rect 36946 37568 37262 37569
rect 36946 37504 36952 37568
rect 37016 37504 37032 37568
rect 37096 37504 37112 37568
rect 37176 37504 37192 37568
rect 37256 37504 37262 37568
rect 36946 37503 37262 37504
rect 2606 37024 2922 37025
rect 2606 36960 2612 37024
rect 2676 36960 2692 37024
rect 2756 36960 2772 37024
rect 2836 36960 2852 37024
rect 2916 36960 2922 37024
rect 2606 36959 2922 36960
rect 7606 37024 7922 37025
rect 7606 36960 7612 37024
rect 7676 36960 7692 37024
rect 7756 36960 7772 37024
rect 7836 36960 7852 37024
rect 7916 36960 7922 37024
rect 7606 36959 7922 36960
rect 12606 37024 12922 37025
rect 12606 36960 12612 37024
rect 12676 36960 12692 37024
rect 12756 36960 12772 37024
rect 12836 36960 12852 37024
rect 12916 36960 12922 37024
rect 12606 36959 12922 36960
rect 17606 37024 17922 37025
rect 17606 36960 17612 37024
rect 17676 36960 17692 37024
rect 17756 36960 17772 37024
rect 17836 36960 17852 37024
rect 17916 36960 17922 37024
rect 17606 36959 17922 36960
rect 22606 37024 22922 37025
rect 22606 36960 22612 37024
rect 22676 36960 22692 37024
rect 22756 36960 22772 37024
rect 22836 36960 22852 37024
rect 22916 36960 22922 37024
rect 22606 36959 22922 36960
rect 27606 37024 27922 37025
rect 27606 36960 27612 37024
rect 27676 36960 27692 37024
rect 27756 36960 27772 37024
rect 27836 36960 27852 37024
rect 27916 36960 27922 37024
rect 27606 36959 27922 36960
rect 32606 37024 32922 37025
rect 32606 36960 32612 37024
rect 32676 36960 32692 37024
rect 32756 36960 32772 37024
rect 32836 36960 32852 37024
rect 32916 36960 32922 37024
rect 32606 36959 32922 36960
rect 37606 37024 37922 37025
rect 37606 36960 37612 37024
rect 37676 36960 37692 37024
rect 37756 36960 37772 37024
rect 37836 36960 37852 37024
rect 37916 36960 37922 37024
rect 37606 36959 37922 36960
rect 4153 36682 4219 36685
rect 23749 36682 23815 36685
rect 4153 36680 23815 36682
rect 4153 36624 4158 36680
rect 4214 36624 23754 36680
rect 23810 36624 23815 36680
rect 4153 36622 23815 36624
rect 4153 36619 4219 36622
rect 23749 36619 23815 36622
rect 1946 36480 2262 36481
rect 1946 36416 1952 36480
rect 2016 36416 2032 36480
rect 2096 36416 2112 36480
rect 2176 36416 2192 36480
rect 2256 36416 2262 36480
rect 1946 36415 2262 36416
rect 6946 36480 7262 36481
rect 6946 36416 6952 36480
rect 7016 36416 7032 36480
rect 7096 36416 7112 36480
rect 7176 36416 7192 36480
rect 7256 36416 7262 36480
rect 6946 36415 7262 36416
rect 11946 36480 12262 36481
rect 11946 36416 11952 36480
rect 12016 36416 12032 36480
rect 12096 36416 12112 36480
rect 12176 36416 12192 36480
rect 12256 36416 12262 36480
rect 11946 36415 12262 36416
rect 16946 36480 17262 36481
rect 16946 36416 16952 36480
rect 17016 36416 17032 36480
rect 17096 36416 17112 36480
rect 17176 36416 17192 36480
rect 17256 36416 17262 36480
rect 16946 36415 17262 36416
rect 21946 36480 22262 36481
rect 21946 36416 21952 36480
rect 22016 36416 22032 36480
rect 22096 36416 22112 36480
rect 22176 36416 22192 36480
rect 22256 36416 22262 36480
rect 21946 36415 22262 36416
rect 26946 36480 27262 36481
rect 26946 36416 26952 36480
rect 27016 36416 27032 36480
rect 27096 36416 27112 36480
rect 27176 36416 27192 36480
rect 27256 36416 27262 36480
rect 26946 36415 27262 36416
rect 31946 36480 32262 36481
rect 31946 36416 31952 36480
rect 32016 36416 32032 36480
rect 32096 36416 32112 36480
rect 32176 36416 32192 36480
rect 32256 36416 32262 36480
rect 31946 36415 32262 36416
rect 36946 36480 37262 36481
rect 36946 36416 36952 36480
rect 37016 36416 37032 36480
rect 37096 36416 37112 36480
rect 37176 36416 37192 36480
rect 37256 36416 37262 36480
rect 36946 36415 37262 36416
rect 2606 35936 2922 35937
rect 2606 35872 2612 35936
rect 2676 35872 2692 35936
rect 2756 35872 2772 35936
rect 2836 35872 2852 35936
rect 2916 35872 2922 35936
rect 2606 35871 2922 35872
rect 7606 35936 7922 35937
rect 7606 35872 7612 35936
rect 7676 35872 7692 35936
rect 7756 35872 7772 35936
rect 7836 35872 7852 35936
rect 7916 35872 7922 35936
rect 7606 35871 7922 35872
rect 12606 35936 12922 35937
rect 12606 35872 12612 35936
rect 12676 35872 12692 35936
rect 12756 35872 12772 35936
rect 12836 35872 12852 35936
rect 12916 35872 12922 35936
rect 12606 35871 12922 35872
rect 17606 35936 17922 35937
rect 17606 35872 17612 35936
rect 17676 35872 17692 35936
rect 17756 35872 17772 35936
rect 17836 35872 17852 35936
rect 17916 35872 17922 35936
rect 17606 35871 17922 35872
rect 22606 35936 22922 35937
rect 22606 35872 22612 35936
rect 22676 35872 22692 35936
rect 22756 35872 22772 35936
rect 22836 35872 22852 35936
rect 22916 35872 22922 35936
rect 22606 35871 22922 35872
rect 27606 35936 27922 35937
rect 27606 35872 27612 35936
rect 27676 35872 27692 35936
rect 27756 35872 27772 35936
rect 27836 35872 27852 35936
rect 27916 35872 27922 35936
rect 27606 35871 27922 35872
rect 32606 35936 32922 35937
rect 32606 35872 32612 35936
rect 32676 35872 32692 35936
rect 32756 35872 32772 35936
rect 32836 35872 32852 35936
rect 32916 35872 32922 35936
rect 32606 35871 32922 35872
rect 37606 35936 37922 35937
rect 37606 35872 37612 35936
rect 37676 35872 37692 35936
rect 37756 35872 37772 35936
rect 37836 35872 37852 35936
rect 37916 35872 37922 35936
rect 37606 35871 37922 35872
rect 1946 35392 2262 35393
rect 1946 35328 1952 35392
rect 2016 35328 2032 35392
rect 2096 35328 2112 35392
rect 2176 35328 2192 35392
rect 2256 35328 2262 35392
rect 1946 35327 2262 35328
rect 6946 35392 7262 35393
rect 6946 35328 6952 35392
rect 7016 35328 7032 35392
rect 7096 35328 7112 35392
rect 7176 35328 7192 35392
rect 7256 35328 7262 35392
rect 6946 35327 7262 35328
rect 11946 35392 12262 35393
rect 11946 35328 11952 35392
rect 12016 35328 12032 35392
rect 12096 35328 12112 35392
rect 12176 35328 12192 35392
rect 12256 35328 12262 35392
rect 11946 35327 12262 35328
rect 16946 35392 17262 35393
rect 16946 35328 16952 35392
rect 17016 35328 17032 35392
rect 17096 35328 17112 35392
rect 17176 35328 17192 35392
rect 17256 35328 17262 35392
rect 16946 35327 17262 35328
rect 21946 35392 22262 35393
rect 21946 35328 21952 35392
rect 22016 35328 22032 35392
rect 22096 35328 22112 35392
rect 22176 35328 22192 35392
rect 22256 35328 22262 35392
rect 21946 35327 22262 35328
rect 26946 35392 27262 35393
rect 26946 35328 26952 35392
rect 27016 35328 27032 35392
rect 27096 35328 27112 35392
rect 27176 35328 27192 35392
rect 27256 35328 27262 35392
rect 26946 35327 27262 35328
rect 31946 35392 32262 35393
rect 31946 35328 31952 35392
rect 32016 35328 32032 35392
rect 32096 35328 32112 35392
rect 32176 35328 32192 35392
rect 32256 35328 32262 35392
rect 31946 35327 32262 35328
rect 36946 35392 37262 35393
rect 36946 35328 36952 35392
rect 37016 35328 37032 35392
rect 37096 35328 37112 35392
rect 37176 35328 37192 35392
rect 37256 35328 37262 35392
rect 36946 35327 37262 35328
rect 6729 35186 6795 35189
rect 15193 35186 15259 35189
rect 6729 35184 15259 35186
rect 6729 35128 6734 35184
rect 6790 35128 15198 35184
rect 15254 35128 15259 35184
rect 6729 35126 15259 35128
rect 6729 35123 6795 35126
rect 15193 35123 15259 35126
rect 8201 35050 8267 35053
rect 8158 35048 8267 35050
rect 8158 34992 8206 35048
rect 8262 34992 8267 35048
rect 8158 34987 8267 34992
rect 2606 34848 2922 34849
rect 2606 34784 2612 34848
rect 2676 34784 2692 34848
rect 2756 34784 2772 34848
rect 2836 34784 2852 34848
rect 2916 34784 2922 34848
rect 2606 34783 2922 34784
rect 7606 34848 7922 34849
rect 7606 34784 7612 34848
rect 7676 34784 7692 34848
rect 7756 34784 7772 34848
rect 7836 34784 7852 34848
rect 7916 34784 7922 34848
rect 7606 34783 7922 34784
rect 8158 34781 8218 34987
rect 12606 34848 12922 34849
rect 12606 34784 12612 34848
rect 12676 34784 12692 34848
rect 12756 34784 12772 34848
rect 12836 34784 12852 34848
rect 12916 34784 12922 34848
rect 12606 34783 12922 34784
rect 17606 34848 17922 34849
rect 17606 34784 17612 34848
rect 17676 34784 17692 34848
rect 17756 34784 17772 34848
rect 17836 34784 17852 34848
rect 17916 34784 17922 34848
rect 17606 34783 17922 34784
rect 22606 34848 22922 34849
rect 22606 34784 22612 34848
rect 22676 34784 22692 34848
rect 22756 34784 22772 34848
rect 22836 34784 22852 34848
rect 22916 34784 22922 34848
rect 22606 34783 22922 34784
rect 27606 34848 27922 34849
rect 27606 34784 27612 34848
rect 27676 34784 27692 34848
rect 27756 34784 27772 34848
rect 27836 34784 27852 34848
rect 27916 34784 27922 34848
rect 27606 34783 27922 34784
rect 32606 34848 32922 34849
rect 32606 34784 32612 34848
rect 32676 34784 32692 34848
rect 32756 34784 32772 34848
rect 32836 34784 32852 34848
rect 32916 34784 32922 34848
rect 32606 34783 32922 34784
rect 37606 34848 37922 34849
rect 37606 34784 37612 34848
rect 37676 34784 37692 34848
rect 37756 34784 37772 34848
rect 37836 34784 37852 34848
rect 37916 34784 37922 34848
rect 37606 34783 37922 34784
rect 7373 34778 7439 34781
rect 7373 34776 7482 34778
rect 7373 34720 7378 34776
rect 7434 34720 7482 34776
rect 7373 34715 7482 34720
rect 8158 34776 8267 34781
rect 8158 34720 8206 34776
rect 8262 34720 8267 34776
rect 8158 34718 8267 34720
rect 8201 34715 8267 34718
rect 7422 34509 7482 34715
rect 7422 34504 7531 34509
rect 7422 34448 7470 34504
rect 7526 34448 7531 34504
rect 7422 34446 7531 34448
rect 7465 34443 7531 34446
rect 1946 34304 2262 34305
rect 1946 34240 1952 34304
rect 2016 34240 2032 34304
rect 2096 34240 2112 34304
rect 2176 34240 2192 34304
rect 2256 34240 2262 34304
rect 1946 34239 2262 34240
rect 6946 34304 7262 34305
rect 6946 34240 6952 34304
rect 7016 34240 7032 34304
rect 7096 34240 7112 34304
rect 7176 34240 7192 34304
rect 7256 34240 7262 34304
rect 6946 34239 7262 34240
rect 11946 34304 12262 34305
rect 11946 34240 11952 34304
rect 12016 34240 12032 34304
rect 12096 34240 12112 34304
rect 12176 34240 12192 34304
rect 12256 34240 12262 34304
rect 11946 34239 12262 34240
rect 16946 34304 17262 34305
rect 16946 34240 16952 34304
rect 17016 34240 17032 34304
rect 17096 34240 17112 34304
rect 17176 34240 17192 34304
rect 17256 34240 17262 34304
rect 16946 34239 17262 34240
rect 21946 34304 22262 34305
rect 21946 34240 21952 34304
rect 22016 34240 22032 34304
rect 22096 34240 22112 34304
rect 22176 34240 22192 34304
rect 22256 34240 22262 34304
rect 21946 34239 22262 34240
rect 26946 34304 27262 34305
rect 26946 34240 26952 34304
rect 27016 34240 27032 34304
rect 27096 34240 27112 34304
rect 27176 34240 27192 34304
rect 27256 34240 27262 34304
rect 26946 34239 27262 34240
rect 31946 34304 32262 34305
rect 31946 34240 31952 34304
rect 32016 34240 32032 34304
rect 32096 34240 32112 34304
rect 32176 34240 32192 34304
rect 32256 34240 32262 34304
rect 31946 34239 32262 34240
rect 36946 34304 37262 34305
rect 36946 34240 36952 34304
rect 37016 34240 37032 34304
rect 37096 34240 37112 34304
rect 37176 34240 37192 34304
rect 37256 34240 37262 34304
rect 36946 34239 37262 34240
rect 2606 33760 2922 33761
rect 2606 33696 2612 33760
rect 2676 33696 2692 33760
rect 2756 33696 2772 33760
rect 2836 33696 2852 33760
rect 2916 33696 2922 33760
rect 2606 33695 2922 33696
rect 7606 33760 7922 33761
rect 7606 33696 7612 33760
rect 7676 33696 7692 33760
rect 7756 33696 7772 33760
rect 7836 33696 7852 33760
rect 7916 33696 7922 33760
rect 7606 33695 7922 33696
rect 12606 33760 12922 33761
rect 12606 33696 12612 33760
rect 12676 33696 12692 33760
rect 12756 33696 12772 33760
rect 12836 33696 12852 33760
rect 12916 33696 12922 33760
rect 12606 33695 12922 33696
rect 17606 33760 17922 33761
rect 17606 33696 17612 33760
rect 17676 33696 17692 33760
rect 17756 33696 17772 33760
rect 17836 33696 17852 33760
rect 17916 33696 17922 33760
rect 17606 33695 17922 33696
rect 22606 33760 22922 33761
rect 22606 33696 22612 33760
rect 22676 33696 22692 33760
rect 22756 33696 22772 33760
rect 22836 33696 22852 33760
rect 22916 33696 22922 33760
rect 22606 33695 22922 33696
rect 27606 33760 27922 33761
rect 27606 33696 27612 33760
rect 27676 33696 27692 33760
rect 27756 33696 27772 33760
rect 27836 33696 27852 33760
rect 27916 33696 27922 33760
rect 27606 33695 27922 33696
rect 32606 33760 32922 33761
rect 32606 33696 32612 33760
rect 32676 33696 32692 33760
rect 32756 33696 32772 33760
rect 32836 33696 32852 33760
rect 32916 33696 32922 33760
rect 32606 33695 32922 33696
rect 37606 33760 37922 33761
rect 37606 33696 37612 33760
rect 37676 33696 37692 33760
rect 37756 33696 37772 33760
rect 37836 33696 37852 33760
rect 37916 33696 37922 33760
rect 37606 33695 37922 33696
rect 1946 33216 2262 33217
rect 1946 33152 1952 33216
rect 2016 33152 2032 33216
rect 2096 33152 2112 33216
rect 2176 33152 2192 33216
rect 2256 33152 2262 33216
rect 1946 33151 2262 33152
rect 6946 33216 7262 33217
rect 6946 33152 6952 33216
rect 7016 33152 7032 33216
rect 7096 33152 7112 33216
rect 7176 33152 7192 33216
rect 7256 33152 7262 33216
rect 6946 33151 7262 33152
rect 11946 33216 12262 33217
rect 11946 33152 11952 33216
rect 12016 33152 12032 33216
rect 12096 33152 12112 33216
rect 12176 33152 12192 33216
rect 12256 33152 12262 33216
rect 11946 33151 12262 33152
rect 16946 33216 17262 33217
rect 16946 33152 16952 33216
rect 17016 33152 17032 33216
rect 17096 33152 17112 33216
rect 17176 33152 17192 33216
rect 17256 33152 17262 33216
rect 16946 33151 17262 33152
rect 21946 33216 22262 33217
rect 21946 33152 21952 33216
rect 22016 33152 22032 33216
rect 22096 33152 22112 33216
rect 22176 33152 22192 33216
rect 22256 33152 22262 33216
rect 21946 33151 22262 33152
rect 26946 33216 27262 33217
rect 26946 33152 26952 33216
rect 27016 33152 27032 33216
rect 27096 33152 27112 33216
rect 27176 33152 27192 33216
rect 27256 33152 27262 33216
rect 26946 33151 27262 33152
rect 31946 33216 32262 33217
rect 31946 33152 31952 33216
rect 32016 33152 32032 33216
rect 32096 33152 32112 33216
rect 32176 33152 32192 33216
rect 32256 33152 32262 33216
rect 31946 33151 32262 33152
rect 36946 33216 37262 33217
rect 36946 33152 36952 33216
rect 37016 33152 37032 33216
rect 37096 33152 37112 33216
rect 37176 33152 37192 33216
rect 37256 33152 37262 33216
rect 36946 33151 37262 33152
rect 2606 32672 2922 32673
rect 2606 32608 2612 32672
rect 2676 32608 2692 32672
rect 2756 32608 2772 32672
rect 2836 32608 2852 32672
rect 2916 32608 2922 32672
rect 2606 32607 2922 32608
rect 7606 32672 7922 32673
rect 7606 32608 7612 32672
rect 7676 32608 7692 32672
rect 7756 32608 7772 32672
rect 7836 32608 7852 32672
rect 7916 32608 7922 32672
rect 7606 32607 7922 32608
rect 12606 32672 12922 32673
rect 12606 32608 12612 32672
rect 12676 32608 12692 32672
rect 12756 32608 12772 32672
rect 12836 32608 12852 32672
rect 12916 32608 12922 32672
rect 12606 32607 12922 32608
rect 17606 32672 17922 32673
rect 17606 32608 17612 32672
rect 17676 32608 17692 32672
rect 17756 32608 17772 32672
rect 17836 32608 17852 32672
rect 17916 32608 17922 32672
rect 17606 32607 17922 32608
rect 22606 32672 22922 32673
rect 22606 32608 22612 32672
rect 22676 32608 22692 32672
rect 22756 32608 22772 32672
rect 22836 32608 22852 32672
rect 22916 32608 22922 32672
rect 22606 32607 22922 32608
rect 27606 32672 27922 32673
rect 27606 32608 27612 32672
rect 27676 32608 27692 32672
rect 27756 32608 27772 32672
rect 27836 32608 27852 32672
rect 27916 32608 27922 32672
rect 27606 32607 27922 32608
rect 32606 32672 32922 32673
rect 32606 32608 32612 32672
rect 32676 32608 32692 32672
rect 32756 32608 32772 32672
rect 32836 32608 32852 32672
rect 32916 32608 32922 32672
rect 32606 32607 32922 32608
rect 37606 32672 37922 32673
rect 37606 32608 37612 32672
rect 37676 32608 37692 32672
rect 37756 32608 37772 32672
rect 37836 32608 37852 32672
rect 37916 32608 37922 32672
rect 37606 32607 37922 32608
rect 1946 32128 2262 32129
rect 1946 32064 1952 32128
rect 2016 32064 2032 32128
rect 2096 32064 2112 32128
rect 2176 32064 2192 32128
rect 2256 32064 2262 32128
rect 1946 32063 2262 32064
rect 6946 32128 7262 32129
rect 6946 32064 6952 32128
rect 7016 32064 7032 32128
rect 7096 32064 7112 32128
rect 7176 32064 7192 32128
rect 7256 32064 7262 32128
rect 6946 32063 7262 32064
rect 11946 32128 12262 32129
rect 11946 32064 11952 32128
rect 12016 32064 12032 32128
rect 12096 32064 12112 32128
rect 12176 32064 12192 32128
rect 12256 32064 12262 32128
rect 11946 32063 12262 32064
rect 16946 32128 17262 32129
rect 16946 32064 16952 32128
rect 17016 32064 17032 32128
rect 17096 32064 17112 32128
rect 17176 32064 17192 32128
rect 17256 32064 17262 32128
rect 16946 32063 17262 32064
rect 21946 32128 22262 32129
rect 21946 32064 21952 32128
rect 22016 32064 22032 32128
rect 22096 32064 22112 32128
rect 22176 32064 22192 32128
rect 22256 32064 22262 32128
rect 21946 32063 22262 32064
rect 26946 32128 27262 32129
rect 26946 32064 26952 32128
rect 27016 32064 27032 32128
rect 27096 32064 27112 32128
rect 27176 32064 27192 32128
rect 27256 32064 27262 32128
rect 26946 32063 27262 32064
rect 31946 32128 32262 32129
rect 31946 32064 31952 32128
rect 32016 32064 32032 32128
rect 32096 32064 32112 32128
rect 32176 32064 32192 32128
rect 32256 32064 32262 32128
rect 31946 32063 32262 32064
rect 36946 32128 37262 32129
rect 36946 32064 36952 32128
rect 37016 32064 37032 32128
rect 37096 32064 37112 32128
rect 37176 32064 37192 32128
rect 37256 32064 37262 32128
rect 36946 32063 37262 32064
rect 2606 31584 2922 31585
rect 2606 31520 2612 31584
rect 2676 31520 2692 31584
rect 2756 31520 2772 31584
rect 2836 31520 2852 31584
rect 2916 31520 2922 31584
rect 2606 31519 2922 31520
rect 7606 31584 7922 31585
rect 7606 31520 7612 31584
rect 7676 31520 7692 31584
rect 7756 31520 7772 31584
rect 7836 31520 7852 31584
rect 7916 31520 7922 31584
rect 7606 31519 7922 31520
rect 12606 31584 12922 31585
rect 12606 31520 12612 31584
rect 12676 31520 12692 31584
rect 12756 31520 12772 31584
rect 12836 31520 12852 31584
rect 12916 31520 12922 31584
rect 12606 31519 12922 31520
rect 17606 31584 17922 31585
rect 17606 31520 17612 31584
rect 17676 31520 17692 31584
rect 17756 31520 17772 31584
rect 17836 31520 17852 31584
rect 17916 31520 17922 31584
rect 17606 31519 17922 31520
rect 22606 31584 22922 31585
rect 22606 31520 22612 31584
rect 22676 31520 22692 31584
rect 22756 31520 22772 31584
rect 22836 31520 22852 31584
rect 22916 31520 22922 31584
rect 22606 31519 22922 31520
rect 27606 31584 27922 31585
rect 27606 31520 27612 31584
rect 27676 31520 27692 31584
rect 27756 31520 27772 31584
rect 27836 31520 27852 31584
rect 27916 31520 27922 31584
rect 27606 31519 27922 31520
rect 32606 31584 32922 31585
rect 32606 31520 32612 31584
rect 32676 31520 32692 31584
rect 32756 31520 32772 31584
rect 32836 31520 32852 31584
rect 32916 31520 32922 31584
rect 32606 31519 32922 31520
rect 37606 31584 37922 31585
rect 37606 31520 37612 31584
rect 37676 31520 37692 31584
rect 37756 31520 37772 31584
rect 37836 31520 37852 31584
rect 37916 31520 37922 31584
rect 37606 31519 37922 31520
rect 0 31378 800 31408
rect 1393 31378 1459 31381
rect 0 31376 1459 31378
rect 0 31320 1398 31376
rect 1454 31320 1459 31376
rect 0 31318 1459 31320
rect 0 31288 800 31318
rect 1393 31315 1459 31318
rect 40493 31378 40559 31381
rect 41200 31378 42000 31408
rect 40493 31376 42000 31378
rect 40493 31320 40498 31376
rect 40554 31320 42000 31376
rect 40493 31318 42000 31320
rect 40493 31315 40559 31318
rect 41200 31288 42000 31318
rect 9489 31242 9555 31245
rect 30598 31242 30604 31244
rect 9489 31240 30604 31242
rect 9489 31184 9494 31240
rect 9550 31184 30604 31240
rect 9489 31182 30604 31184
rect 9489 31179 9555 31182
rect 30598 31180 30604 31182
rect 30668 31180 30674 31244
rect 23238 31044 23244 31108
rect 23308 31106 23314 31108
rect 23381 31106 23447 31109
rect 23308 31104 23447 31106
rect 23308 31048 23386 31104
rect 23442 31048 23447 31104
rect 23308 31046 23447 31048
rect 23308 31044 23314 31046
rect 23381 31043 23447 31046
rect 1946 31040 2262 31041
rect 1946 30976 1952 31040
rect 2016 30976 2032 31040
rect 2096 30976 2112 31040
rect 2176 30976 2192 31040
rect 2256 30976 2262 31040
rect 1946 30975 2262 30976
rect 6946 31040 7262 31041
rect 6946 30976 6952 31040
rect 7016 30976 7032 31040
rect 7096 30976 7112 31040
rect 7176 30976 7192 31040
rect 7256 30976 7262 31040
rect 6946 30975 7262 30976
rect 11946 31040 12262 31041
rect 11946 30976 11952 31040
rect 12016 30976 12032 31040
rect 12096 30976 12112 31040
rect 12176 30976 12192 31040
rect 12256 30976 12262 31040
rect 11946 30975 12262 30976
rect 16946 31040 17262 31041
rect 16946 30976 16952 31040
rect 17016 30976 17032 31040
rect 17096 30976 17112 31040
rect 17176 30976 17192 31040
rect 17256 30976 17262 31040
rect 16946 30975 17262 30976
rect 21946 31040 22262 31041
rect 21946 30976 21952 31040
rect 22016 30976 22032 31040
rect 22096 30976 22112 31040
rect 22176 30976 22192 31040
rect 22256 30976 22262 31040
rect 21946 30975 22262 30976
rect 26946 31040 27262 31041
rect 26946 30976 26952 31040
rect 27016 30976 27032 31040
rect 27096 30976 27112 31040
rect 27176 30976 27192 31040
rect 27256 30976 27262 31040
rect 26946 30975 27262 30976
rect 31946 31040 32262 31041
rect 31946 30976 31952 31040
rect 32016 30976 32032 31040
rect 32096 30976 32112 31040
rect 32176 30976 32192 31040
rect 32256 30976 32262 31040
rect 31946 30975 32262 30976
rect 36946 31040 37262 31041
rect 36946 30976 36952 31040
rect 37016 30976 37032 31040
rect 37096 30976 37112 31040
rect 37176 30976 37192 31040
rect 37256 30976 37262 31040
rect 36946 30975 37262 30976
rect 2606 30496 2922 30497
rect 2606 30432 2612 30496
rect 2676 30432 2692 30496
rect 2756 30432 2772 30496
rect 2836 30432 2852 30496
rect 2916 30432 2922 30496
rect 2606 30431 2922 30432
rect 7606 30496 7922 30497
rect 7606 30432 7612 30496
rect 7676 30432 7692 30496
rect 7756 30432 7772 30496
rect 7836 30432 7852 30496
rect 7916 30432 7922 30496
rect 7606 30431 7922 30432
rect 12606 30496 12922 30497
rect 12606 30432 12612 30496
rect 12676 30432 12692 30496
rect 12756 30432 12772 30496
rect 12836 30432 12852 30496
rect 12916 30432 12922 30496
rect 12606 30431 12922 30432
rect 17606 30496 17922 30497
rect 17606 30432 17612 30496
rect 17676 30432 17692 30496
rect 17756 30432 17772 30496
rect 17836 30432 17852 30496
rect 17916 30432 17922 30496
rect 17606 30431 17922 30432
rect 22606 30496 22922 30497
rect 22606 30432 22612 30496
rect 22676 30432 22692 30496
rect 22756 30432 22772 30496
rect 22836 30432 22852 30496
rect 22916 30432 22922 30496
rect 22606 30431 22922 30432
rect 27606 30496 27922 30497
rect 27606 30432 27612 30496
rect 27676 30432 27692 30496
rect 27756 30432 27772 30496
rect 27836 30432 27852 30496
rect 27916 30432 27922 30496
rect 27606 30431 27922 30432
rect 32606 30496 32922 30497
rect 32606 30432 32612 30496
rect 32676 30432 32692 30496
rect 32756 30432 32772 30496
rect 32836 30432 32852 30496
rect 32916 30432 32922 30496
rect 32606 30431 32922 30432
rect 37606 30496 37922 30497
rect 37606 30432 37612 30496
rect 37676 30432 37692 30496
rect 37756 30432 37772 30496
rect 37836 30432 37852 30496
rect 37916 30432 37922 30496
rect 37606 30431 37922 30432
rect 1946 29952 2262 29953
rect 1946 29888 1952 29952
rect 2016 29888 2032 29952
rect 2096 29888 2112 29952
rect 2176 29888 2192 29952
rect 2256 29888 2262 29952
rect 1946 29887 2262 29888
rect 6946 29952 7262 29953
rect 6946 29888 6952 29952
rect 7016 29888 7032 29952
rect 7096 29888 7112 29952
rect 7176 29888 7192 29952
rect 7256 29888 7262 29952
rect 6946 29887 7262 29888
rect 11946 29952 12262 29953
rect 11946 29888 11952 29952
rect 12016 29888 12032 29952
rect 12096 29888 12112 29952
rect 12176 29888 12192 29952
rect 12256 29888 12262 29952
rect 11946 29887 12262 29888
rect 16946 29952 17262 29953
rect 16946 29888 16952 29952
rect 17016 29888 17032 29952
rect 17096 29888 17112 29952
rect 17176 29888 17192 29952
rect 17256 29888 17262 29952
rect 16946 29887 17262 29888
rect 21946 29952 22262 29953
rect 21946 29888 21952 29952
rect 22016 29888 22032 29952
rect 22096 29888 22112 29952
rect 22176 29888 22192 29952
rect 22256 29888 22262 29952
rect 21946 29887 22262 29888
rect 26946 29952 27262 29953
rect 26946 29888 26952 29952
rect 27016 29888 27032 29952
rect 27096 29888 27112 29952
rect 27176 29888 27192 29952
rect 27256 29888 27262 29952
rect 26946 29887 27262 29888
rect 31946 29952 32262 29953
rect 31946 29888 31952 29952
rect 32016 29888 32032 29952
rect 32096 29888 32112 29952
rect 32176 29888 32192 29952
rect 32256 29888 32262 29952
rect 31946 29887 32262 29888
rect 36946 29952 37262 29953
rect 36946 29888 36952 29952
rect 37016 29888 37032 29952
rect 37096 29888 37112 29952
rect 37176 29888 37192 29952
rect 37256 29888 37262 29952
rect 36946 29887 37262 29888
rect 2606 29408 2922 29409
rect 2606 29344 2612 29408
rect 2676 29344 2692 29408
rect 2756 29344 2772 29408
rect 2836 29344 2852 29408
rect 2916 29344 2922 29408
rect 2606 29343 2922 29344
rect 7606 29408 7922 29409
rect 7606 29344 7612 29408
rect 7676 29344 7692 29408
rect 7756 29344 7772 29408
rect 7836 29344 7852 29408
rect 7916 29344 7922 29408
rect 7606 29343 7922 29344
rect 12606 29408 12922 29409
rect 12606 29344 12612 29408
rect 12676 29344 12692 29408
rect 12756 29344 12772 29408
rect 12836 29344 12852 29408
rect 12916 29344 12922 29408
rect 12606 29343 12922 29344
rect 17606 29408 17922 29409
rect 17606 29344 17612 29408
rect 17676 29344 17692 29408
rect 17756 29344 17772 29408
rect 17836 29344 17852 29408
rect 17916 29344 17922 29408
rect 17606 29343 17922 29344
rect 22606 29408 22922 29409
rect 22606 29344 22612 29408
rect 22676 29344 22692 29408
rect 22756 29344 22772 29408
rect 22836 29344 22852 29408
rect 22916 29344 22922 29408
rect 22606 29343 22922 29344
rect 27606 29408 27922 29409
rect 27606 29344 27612 29408
rect 27676 29344 27692 29408
rect 27756 29344 27772 29408
rect 27836 29344 27852 29408
rect 27916 29344 27922 29408
rect 27606 29343 27922 29344
rect 32606 29408 32922 29409
rect 32606 29344 32612 29408
rect 32676 29344 32692 29408
rect 32756 29344 32772 29408
rect 32836 29344 32852 29408
rect 32916 29344 32922 29408
rect 32606 29343 32922 29344
rect 37606 29408 37922 29409
rect 37606 29344 37612 29408
rect 37676 29344 37692 29408
rect 37756 29344 37772 29408
rect 37836 29344 37852 29408
rect 37916 29344 37922 29408
rect 37606 29343 37922 29344
rect 1946 28864 2262 28865
rect 1946 28800 1952 28864
rect 2016 28800 2032 28864
rect 2096 28800 2112 28864
rect 2176 28800 2192 28864
rect 2256 28800 2262 28864
rect 1946 28799 2262 28800
rect 6946 28864 7262 28865
rect 6946 28800 6952 28864
rect 7016 28800 7032 28864
rect 7096 28800 7112 28864
rect 7176 28800 7192 28864
rect 7256 28800 7262 28864
rect 6946 28799 7262 28800
rect 11946 28864 12262 28865
rect 11946 28800 11952 28864
rect 12016 28800 12032 28864
rect 12096 28800 12112 28864
rect 12176 28800 12192 28864
rect 12256 28800 12262 28864
rect 11946 28799 12262 28800
rect 16946 28864 17262 28865
rect 16946 28800 16952 28864
rect 17016 28800 17032 28864
rect 17096 28800 17112 28864
rect 17176 28800 17192 28864
rect 17256 28800 17262 28864
rect 16946 28799 17262 28800
rect 21946 28864 22262 28865
rect 21946 28800 21952 28864
rect 22016 28800 22032 28864
rect 22096 28800 22112 28864
rect 22176 28800 22192 28864
rect 22256 28800 22262 28864
rect 21946 28799 22262 28800
rect 26946 28864 27262 28865
rect 26946 28800 26952 28864
rect 27016 28800 27032 28864
rect 27096 28800 27112 28864
rect 27176 28800 27192 28864
rect 27256 28800 27262 28864
rect 26946 28799 27262 28800
rect 31946 28864 32262 28865
rect 31946 28800 31952 28864
rect 32016 28800 32032 28864
rect 32096 28800 32112 28864
rect 32176 28800 32192 28864
rect 32256 28800 32262 28864
rect 31946 28799 32262 28800
rect 36946 28864 37262 28865
rect 36946 28800 36952 28864
rect 37016 28800 37032 28864
rect 37096 28800 37112 28864
rect 37176 28800 37192 28864
rect 37256 28800 37262 28864
rect 36946 28799 37262 28800
rect 2606 28320 2922 28321
rect 2606 28256 2612 28320
rect 2676 28256 2692 28320
rect 2756 28256 2772 28320
rect 2836 28256 2852 28320
rect 2916 28256 2922 28320
rect 2606 28255 2922 28256
rect 7606 28320 7922 28321
rect 7606 28256 7612 28320
rect 7676 28256 7692 28320
rect 7756 28256 7772 28320
rect 7836 28256 7852 28320
rect 7916 28256 7922 28320
rect 7606 28255 7922 28256
rect 12606 28320 12922 28321
rect 12606 28256 12612 28320
rect 12676 28256 12692 28320
rect 12756 28256 12772 28320
rect 12836 28256 12852 28320
rect 12916 28256 12922 28320
rect 12606 28255 12922 28256
rect 17606 28320 17922 28321
rect 17606 28256 17612 28320
rect 17676 28256 17692 28320
rect 17756 28256 17772 28320
rect 17836 28256 17852 28320
rect 17916 28256 17922 28320
rect 17606 28255 17922 28256
rect 22606 28320 22922 28321
rect 22606 28256 22612 28320
rect 22676 28256 22692 28320
rect 22756 28256 22772 28320
rect 22836 28256 22852 28320
rect 22916 28256 22922 28320
rect 22606 28255 22922 28256
rect 27606 28320 27922 28321
rect 27606 28256 27612 28320
rect 27676 28256 27692 28320
rect 27756 28256 27772 28320
rect 27836 28256 27852 28320
rect 27916 28256 27922 28320
rect 27606 28255 27922 28256
rect 32606 28320 32922 28321
rect 32606 28256 32612 28320
rect 32676 28256 32692 28320
rect 32756 28256 32772 28320
rect 32836 28256 32852 28320
rect 32916 28256 32922 28320
rect 32606 28255 32922 28256
rect 37606 28320 37922 28321
rect 37606 28256 37612 28320
rect 37676 28256 37692 28320
rect 37756 28256 37772 28320
rect 37836 28256 37852 28320
rect 37916 28256 37922 28320
rect 37606 28255 37922 28256
rect 1946 27776 2262 27777
rect 1946 27712 1952 27776
rect 2016 27712 2032 27776
rect 2096 27712 2112 27776
rect 2176 27712 2192 27776
rect 2256 27712 2262 27776
rect 1946 27711 2262 27712
rect 6946 27776 7262 27777
rect 6946 27712 6952 27776
rect 7016 27712 7032 27776
rect 7096 27712 7112 27776
rect 7176 27712 7192 27776
rect 7256 27712 7262 27776
rect 6946 27711 7262 27712
rect 11946 27776 12262 27777
rect 11946 27712 11952 27776
rect 12016 27712 12032 27776
rect 12096 27712 12112 27776
rect 12176 27712 12192 27776
rect 12256 27712 12262 27776
rect 11946 27711 12262 27712
rect 16946 27776 17262 27777
rect 16946 27712 16952 27776
rect 17016 27712 17032 27776
rect 17096 27712 17112 27776
rect 17176 27712 17192 27776
rect 17256 27712 17262 27776
rect 16946 27711 17262 27712
rect 21946 27776 22262 27777
rect 21946 27712 21952 27776
rect 22016 27712 22032 27776
rect 22096 27712 22112 27776
rect 22176 27712 22192 27776
rect 22256 27712 22262 27776
rect 21946 27711 22262 27712
rect 26946 27776 27262 27777
rect 26946 27712 26952 27776
rect 27016 27712 27032 27776
rect 27096 27712 27112 27776
rect 27176 27712 27192 27776
rect 27256 27712 27262 27776
rect 26946 27711 27262 27712
rect 31946 27776 32262 27777
rect 31946 27712 31952 27776
rect 32016 27712 32032 27776
rect 32096 27712 32112 27776
rect 32176 27712 32192 27776
rect 32256 27712 32262 27776
rect 31946 27711 32262 27712
rect 36946 27776 37262 27777
rect 36946 27712 36952 27776
rect 37016 27712 37032 27776
rect 37096 27712 37112 27776
rect 37176 27712 37192 27776
rect 37256 27712 37262 27776
rect 36946 27711 37262 27712
rect 2606 27232 2922 27233
rect 2606 27168 2612 27232
rect 2676 27168 2692 27232
rect 2756 27168 2772 27232
rect 2836 27168 2852 27232
rect 2916 27168 2922 27232
rect 2606 27167 2922 27168
rect 7606 27232 7922 27233
rect 7606 27168 7612 27232
rect 7676 27168 7692 27232
rect 7756 27168 7772 27232
rect 7836 27168 7852 27232
rect 7916 27168 7922 27232
rect 7606 27167 7922 27168
rect 12606 27232 12922 27233
rect 12606 27168 12612 27232
rect 12676 27168 12692 27232
rect 12756 27168 12772 27232
rect 12836 27168 12852 27232
rect 12916 27168 12922 27232
rect 12606 27167 12922 27168
rect 17606 27232 17922 27233
rect 17606 27168 17612 27232
rect 17676 27168 17692 27232
rect 17756 27168 17772 27232
rect 17836 27168 17852 27232
rect 17916 27168 17922 27232
rect 17606 27167 17922 27168
rect 22606 27232 22922 27233
rect 22606 27168 22612 27232
rect 22676 27168 22692 27232
rect 22756 27168 22772 27232
rect 22836 27168 22852 27232
rect 22916 27168 22922 27232
rect 22606 27167 22922 27168
rect 27606 27232 27922 27233
rect 27606 27168 27612 27232
rect 27676 27168 27692 27232
rect 27756 27168 27772 27232
rect 27836 27168 27852 27232
rect 27916 27168 27922 27232
rect 27606 27167 27922 27168
rect 32606 27232 32922 27233
rect 32606 27168 32612 27232
rect 32676 27168 32692 27232
rect 32756 27168 32772 27232
rect 32836 27168 32852 27232
rect 32916 27168 32922 27232
rect 32606 27167 32922 27168
rect 37606 27232 37922 27233
rect 37606 27168 37612 27232
rect 37676 27168 37692 27232
rect 37756 27168 37772 27232
rect 37836 27168 37852 27232
rect 37916 27168 37922 27232
rect 37606 27167 37922 27168
rect 17309 27026 17375 27029
rect 17174 27024 17375 27026
rect 17174 26968 17314 27024
rect 17370 26968 17375 27024
rect 17174 26966 17375 26968
rect 16573 26890 16639 26893
rect 17174 26890 17234 26966
rect 17309 26963 17375 26966
rect 16573 26888 17234 26890
rect 16573 26832 16578 26888
rect 16634 26832 17234 26888
rect 16573 26830 17234 26832
rect 16573 26827 16639 26830
rect 1946 26688 2262 26689
rect 1946 26624 1952 26688
rect 2016 26624 2032 26688
rect 2096 26624 2112 26688
rect 2176 26624 2192 26688
rect 2256 26624 2262 26688
rect 1946 26623 2262 26624
rect 6946 26688 7262 26689
rect 6946 26624 6952 26688
rect 7016 26624 7032 26688
rect 7096 26624 7112 26688
rect 7176 26624 7192 26688
rect 7256 26624 7262 26688
rect 6946 26623 7262 26624
rect 11946 26688 12262 26689
rect 11946 26624 11952 26688
rect 12016 26624 12032 26688
rect 12096 26624 12112 26688
rect 12176 26624 12192 26688
rect 12256 26624 12262 26688
rect 11946 26623 12262 26624
rect 16946 26688 17262 26689
rect 16946 26624 16952 26688
rect 17016 26624 17032 26688
rect 17096 26624 17112 26688
rect 17176 26624 17192 26688
rect 17256 26624 17262 26688
rect 16946 26623 17262 26624
rect 21946 26688 22262 26689
rect 21946 26624 21952 26688
rect 22016 26624 22032 26688
rect 22096 26624 22112 26688
rect 22176 26624 22192 26688
rect 22256 26624 22262 26688
rect 21946 26623 22262 26624
rect 26946 26688 27262 26689
rect 26946 26624 26952 26688
rect 27016 26624 27032 26688
rect 27096 26624 27112 26688
rect 27176 26624 27192 26688
rect 27256 26624 27262 26688
rect 26946 26623 27262 26624
rect 31946 26688 32262 26689
rect 31946 26624 31952 26688
rect 32016 26624 32032 26688
rect 32096 26624 32112 26688
rect 32176 26624 32192 26688
rect 32256 26624 32262 26688
rect 31946 26623 32262 26624
rect 36946 26688 37262 26689
rect 36946 26624 36952 26688
rect 37016 26624 37032 26688
rect 37096 26624 37112 26688
rect 37176 26624 37192 26688
rect 37256 26624 37262 26688
rect 36946 26623 37262 26624
rect 18454 26284 18460 26348
rect 18524 26346 18530 26348
rect 24945 26346 25011 26349
rect 18524 26344 25011 26346
rect 18524 26288 24950 26344
rect 25006 26288 25011 26344
rect 18524 26286 25011 26288
rect 18524 26284 18530 26286
rect 24945 26283 25011 26286
rect 2606 26144 2922 26145
rect 2606 26080 2612 26144
rect 2676 26080 2692 26144
rect 2756 26080 2772 26144
rect 2836 26080 2852 26144
rect 2916 26080 2922 26144
rect 2606 26079 2922 26080
rect 7606 26144 7922 26145
rect 7606 26080 7612 26144
rect 7676 26080 7692 26144
rect 7756 26080 7772 26144
rect 7836 26080 7852 26144
rect 7916 26080 7922 26144
rect 7606 26079 7922 26080
rect 12606 26144 12922 26145
rect 12606 26080 12612 26144
rect 12676 26080 12692 26144
rect 12756 26080 12772 26144
rect 12836 26080 12852 26144
rect 12916 26080 12922 26144
rect 12606 26079 12922 26080
rect 17606 26144 17922 26145
rect 17606 26080 17612 26144
rect 17676 26080 17692 26144
rect 17756 26080 17772 26144
rect 17836 26080 17852 26144
rect 17916 26080 17922 26144
rect 17606 26079 17922 26080
rect 22606 26144 22922 26145
rect 22606 26080 22612 26144
rect 22676 26080 22692 26144
rect 22756 26080 22772 26144
rect 22836 26080 22852 26144
rect 22916 26080 22922 26144
rect 22606 26079 22922 26080
rect 27606 26144 27922 26145
rect 27606 26080 27612 26144
rect 27676 26080 27692 26144
rect 27756 26080 27772 26144
rect 27836 26080 27852 26144
rect 27916 26080 27922 26144
rect 27606 26079 27922 26080
rect 32606 26144 32922 26145
rect 32606 26080 32612 26144
rect 32676 26080 32692 26144
rect 32756 26080 32772 26144
rect 32836 26080 32852 26144
rect 32916 26080 32922 26144
rect 32606 26079 32922 26080
rect 37606 26144 37922 26145
rect 37606 26080 37612 26144
rect 37676 26080 37692 26144
rect 37756 26080 37772 26144
rect 37836 26080 37852 26144
rect 37916 26080 37922 26144
rect 37606 26079 37922 26080
rect 1946 25600 2262 25601
rect 1946 25536 1952 25600
rect 2016 25536 2032 25600
rect 2096 25536 2112 25600
rect 2176 25536 2192 25600
rect 2256 25536 2262 25600
rect 1946 25535 2262 25536
rect 6946 25600 7262 25601
rect 6946 25536 6952 25600
rect 7016 25536 7032 25600
rect 7096 25536 7112 25600
rect 7176 25536 7192 25600
rect 7256 25536 7262 25600
rect 6946 25535 7262 25536
rect 11946 25600 12262 25601
rect 11946 25536 11952 25600
rect 12016 25536 12032 25600
rect 12096 25536 12112 25600
rect 12176 25536 12192 25600
rect 12256 25536 12262 25600
rect 11946 25535 12262 25536
rect 16946 25600 17262 25601
rect 16946 25536 16952 25600
rect 17016 25536 17032 25600
rect 17096 25536 17112 25600
rect 17176 25536 17192 25600
rect 17256 25536 17262 25600
rect 16946 25535 17262 25536
rect 21946 25600 22262 25601
rect 21946 25536 21952 25600
rect 22016 25536 22032 25600
rect 22096 25536 22112 25600
rect 22176 25536 22192 25600
rect 22256 25536 22262 25600
rect 21946 25535 22262 25536
rect 26946 25600 27262 25601
rect 26946 25536 26952 25600
rect 27016 25536 27032 25600
rect 27096 25536 27112 25600
rect 27176 25536 27192 25600
rect 27256 25536 27262 25600
rect 26946 25535 27262 25536
rect 31946 25600 32262 25601
rect 31946 25536 31952 25600
rect 32016 25536 32032 25600
rect 32096 25536 32112 25600
rect 32176 25536 32192 25600
rect 32256 25536 32262 25600
rect 31946 25535 32262 25536
rect 36946 25600 37262 25601
rect 36946 25536 36952 25600
rect 37016 25536 37032 25600
rect 37096 25536 37112 25600
rect 37176 25536 37192 25600
rect 37256 25536 37262 25600
rect 36946 25535 37262 25536
rect 2606 25056 2922 25057
rect 2606 24992 2612 25056
rect 2676 24992 2692 25056
rect 2756 24992 2772 25056
rect 2836 24992 2852 25056
rect 2916 24992 2922 25056
rect 2606 24991 2922 24992
rect 7606 25056 7922 25057
rect 7606 24992 7612 25056
rect 7676 24992 7692 25056
rect 7756 24992 7772 25056
rect 7836 24992 7852 25056
rect 7916 24992 7922 25056
rect 7606 24991 7922 24992
rect 12606 25056 12922 25057
rect 12606 24992 12612 25056
rect 12676 24992 12692 25056
rect 12756 24992 12772 25056
rect 12836 24992 12852 25056
rect 12916 24992 12922 25056
rect 12606 24991 12922 24992
rect 17606 25056 17922 25057
rect 17606 24992 17612 25056
rect 17676 24992 17692 25056
rect 17756 24992 17772 25056
rect 17836 24992 17852 25056
rect 17916 24992 17922 25056
rect 17606 24991 17922 24992
rect 22606 25056 22922 25057
rect 22606 24992 22612 25056
rect 22676 24992 22692 25056
rect 22756 24992 22772 25056
rect 22836 24992 22852 25056
rect 22916 24992 22922 25056
rect 22606 24991 22922 24992
rect 27606 25056 27922 25057
rect 27606 24992 27612 25056
rect 27676 24992 27692 25056
rect 27756 24992 27772 25056
rect 27836 24992 27852 25056
rect 27916 24992 27922 25056
rect 27606 24991 27922 24992
rect 32606 25056 32922 25057
rect 32606 24992 32612 25056
rect 32676 24992 32692 25056
rect 32756 24992 32772 25056
rect 32836 24992 32852 25056
rect 32916 24992 32922 25056
rect 32606 24991 32922 24992
rect 37606 25056 37922 25057
rect 37606 24992 37612 25056
rect 37676 24992 37692 25056
rect 37756 24992 37772 25056
rect 37836 24992 37852 25056
rect 37916 24992 37922 25056
rect 37606 24991 37922 24992
rect 1946 24512 2262 24513
rect 1946 24448 1952 24512
rect 2016 24448 2032 24512
rect 2096 24448 2112 24512
rect 2176 24448 2192 24512
rect 2256 24448 2262 24512
rect 1946 24447 2262 24448
rect 6946 24512 7262 24513
rect 6946 24448 6952 24512
rect 7016 24448 7032 24512
rect 7096 24448 7112 24512
rect 7176 24448 7192 24512
rect 7256 24448 7262 24512
rect 6946 24447 7262 24448
rect 11946 24512 12262 24513
rect 11946 24448 11952 24512
rect 12016 24448 12032 24512
rect 12096 24448 12112 24512
rect 12176 24448 12192 24512
rect 12256 24448 12262 24512
rect 11946 24447 12262 24448
rect 16946 24512 17262 24513
rect 16946 24448 16952 24512
rect 17016 24448 17032 24512
rect 17096 24448 17112 24512
rect 17176 24448 17192 24512
rect 17256 24448 17262 24512
rect 16946 24447 17262 24448
rect 21946 24512 22262 24513
rect 21946 24448 21952 24512
rect 22016 24448 22032 24512
rect 22096 24448 22112 24512
rect 22176 24448 22192 24512
rect 22256 24448 22262 24512
rect 21946 24447 22262 24448
rect 26946 24512 27262 24513
rect 26946 24448 26952 24512
rect 27016 24448 27032 24512
rect 27096 24448 27112 24512
rect 27176 24448 27192 24512
rect 27256 24448 27262 24512
rect 26946 24447 27262 24448
rect 31946 24512 32262 24513
rect 31946 24448 31952 24512
rect 32016 24448 32032 24512
rect 32096 24448 32112 24512
rect 32176 24448 32192 24512
rect 32256 24448 32262 24512
rect 31946 24447 32262 24448
rect 36946 24512 37262 24513
rect 36946 24448 36952 24512
rect 37016 24448 37032 24512
rect 37096 24448 37112 24512
rect 37176 24448 37192 24512
rect 37256 24448 37262 24512
rect 36946 24447 37262 24448
rect 2606 23968 2922 23969
rect 2606 23904 2612 23968
rect 2676 23904 2692 23968
rect 2756 23904 2772 23968
rect 2836 23904 2852 23968
rect 2916 23904 2922 23968
rect 2606 23903 2922 23904
rect 7606 23968 7922 23969
rect 7606 23904 7612 23968
rect 7676 23904 7692 23968
rect 7756 23904 7772 23968
rect 7836 23904 7852 23968
rect 7916 23904 7922 23968
rect 7606 23903 7922 23904
rect 12606 23968 12922 23969
rect 12606 23904 12612 23968
rect 12676 23904 12692 23968
rect 12756 23904 12772 23968
rect 12836 23904 12852 23968
rect 12916 23904 12922 23968
rect 12606 23903 12922 23904
rect 17606 23968 17922 23969
rect 17606 23904 17612 23968
rect 17676 23904 17692 23968
rect 17756 23904 17772 23968
rect 17836 23904 17852 23968
rect 17916 23904 17922 23968
rect 17606 23903 17922 23904
rect 22606 23968 22922 23969
rect 22606 23904 22612 23968
rect 22676 23904 22692 23968
rect 22756 23904 22772 23968
rect 22836 23904 22852 23968
rect 22916 23904 22922 23968
rect 22606 23903 22922 23904
rect 27606 23968 27922 23969
rect 27606 23904 27612 23968
rect 27676 23904 27692 23968
rect 27756 23904 27772 23968
rect 27836 23904 27852 23968
rect 27916 23904 27922 23968
rect 27606 23903 27922 23904
rect 32606 23968 32922 23969
rect 32606 23904 32612 23968
rect 32676 23904 32692 23968
rect 32756 23904 32772 23968
rect 32836 23904 32852 23968
rect 32916 23904 32922 23968
rect 32606 23903 32922 23904
rect 37606 23968 37922 23969
rect 37606 23904 37612 23968
rect 37676 23904 37692 23968
rect 37756 23904 37772 23968
rect 37836 23904 37852 23968
rect 37916 23904 37922 23968
rect 37606 23903 37922 23904
rect 1946 23424 2262 23425
rect 1946 23360 1952 23424
rect 2016 23360 2032 23424
rect 2096 23360 2112 23424
rect 2176 23360 2192 23424
rect 2256 23360 2262 23424
rect 1946 23359 2262 23360
rect 6946 23424 7262 23425
rect 6946 23360 6952 23424
rect 7016 23360 7032 23424
rect 7096 23360 7112 23424
rect 7176 23360 7192 23424
rect 7256 23360 7262 23424
rect 6946 23359 7262 23360
rect 11946 23424 12262 23425
rect 11946 23360 11952 23424
rect 12016 23360 12032 23424
rect 12096 23360 12112 23424
rect 12176 23360 12192 23424
rect 12256 23360 12262 23424
rect 11946 23359 12262 23360
rect 16946 23424 17262 23425
rect 16946 23360 16952 23424
rect 17016 23360 17032 23424
rect 17096 23360 17112 23424
rect 17176 23360 17192 23424
rect 17256 23360 17262 23424
rect 16946 23359 17262 23360
rect 21946 23424 22262 23425
rect 21946 23360 21952 23424
rect 22016 23360 22032 23424
rect 22096 23360 22112 23424
rect 22176 23360 22192 23424
rect 22256 23360 22262 23424
rect 21946 23359 22262 23360
rect 26946 23424 27262 23425
rect 26946 23360 26952 23424
rect 27016 23360 27032 23424
rect 27096 23360 27112 23424
rect 27176 23360 27192 23424
rect 27256 23360 27262 23424
rect 26946 23359 27262 23360
rect 31946 23424 32262 23425
rect 31946 23360 31952 23424
rect 32016 23360 32032 23424
rect 32096 23360 32112 23424
rect 32176 23360 32192 23424
rect 32256 23360 32262 23424
rect 31946 23359 32262 23360
rect 36946 23424 37262 23425
rect 36946 23360 36952 23424
rect 37016 23360 37032 23424
rect 37096 23360 37112 23424
rect 37176 23360 37192 23424
rect 37256 23360 37262 23424
rect 36946 23359 37262 23360
rect 2606 22880 2922 22881
rect 2606 22816 2612 22880
rect 2676 22816 2692 22880
rect 2756 22816 2772 22880
rect 2836 22816 2852 22880
rect 2916 22816 2922 22880
rect 2606 22815 2922 22816
rect 7606 22880 7922 22881
rect 7606 22816 7612 22880
rect 7676 22816 7692 22880
rect 7756 22816 7772 22880
rect 7836 22816 7852 22880
rect 7916 22816 7922 22880
rect 7606 22815 7922 22816
rect 12606 22880 12922 22881
rect 12606 22816 12612 22880
rect 12676 22816 12692 22880
rect 12756 22816 12772 22880
rect 12836 22816 12852 22880
rect 12916 22816 12922 22880
rect 12606 22815 12922 22816
rect 17606 22880 17922 22881
rect 17606 22816 17612 22880
rect 17676 22816 17692 22880
rect 17756 22816 17772 22880
rect 17836 22816 17852 22880
rect 17916 22816 17922 22880
rect 17606 22815 17922 22816
rect 22606 22880 22922 22881
rect 22606 22816 22612 22880
rect 22676 22816 22692 22880
rect 22756 22816 22772 22880
rect 22836 22816 22852 22880
rect 22916 22816 22922 22880
rect 22606 22815 22922 22816
rect 27606 22880 27922 22881
rect 27606 22816 27612 22880
rect 27676 22816 27692 22880
rect 27756 22816 27772 22880
rect 27836 22816 27852 22880
rect 27916 22816 27922 22880
rect 27606 22815 27922 22816
rect 32606 22880 32922 22881
rect 32606 22816 32612 22880
rect 32676 22816 32692 22880
rect 32756 22816 32772 22880
rect 32836 22816 32852 22880
rect 32916 22816 32922 22880
rect 32606 22815 32922 22816
rect 37606 22880 37922 22881
rect 37606 22816 37612 22880
rect 37676 22816 37692 22880
rect 37756 22816 37772 22880
rect 37836 22816 37852 22880
rect 37916 22816 37922 22880
rect 37606 22815 37922 22816
rect 14917 22812 14983 22813
rect 14917 22810 14964 22812
rect 14872 22808 14964 22810
rect 14872 22752 14922 22808
rect 14872 22750 14964 22752
rect 14917 22748 14964 22750
rect 15028 22748 15034 22812
rect 14917 22747 14983 22748
rect 841 22538 907 22541
rect 798 22536 907 22538
rect 798 22480 846 22536
rect 902 22480 907 22536
rect 798 22475 907 22480
rect 798 22432 858 22475
rect 0 22342 858 22432
rect 40493 22402 40559 22405
rect 41200 22402 42000 22432
rect 40493 22400 42000 22402
rect 40493 22344 40498 22400
rect 40554 22344 42000 22400
rect 40493 22342 42000 22344
rect 0 22312 800 22342
rect 40493 22339 40559 22342
rect 1946 22336 2262 22337
rect 1946 22272 1952 22336
rect 2016 22272 2032 22336
rect 2096 22272 2112 22336
rect 2176 22272 2192 22336
rect 2256 22272 2262 22336
rect 1946 22271 2262 22272
rect 6946 22336 7262 22337
rect 6946 22272 6952 22336
rect 7016 22272 7032 22336
rect 7096 22272 7112 22336
rect 7176 22272 7192 22336
rect 7256 22272 7262 22336
rect 6946 22271 7262 22272
rect 11946 22336 12262 22337
rect 11946 22272 11952 22336
rect 12016 22272 12032 22336
rect 12096 22272 12112 22336
rect 12176 22272 12192 22336
rect 12256 22272 12262 22336
rect 11946 22271 12262 22272
rect 16946 22336 17262 22337
rect 16946 22272 16952 22336
rect 17016 22272 17032 22336
rect 17096 22272 17112 22336
rect 17176 22272 17192 22336
rect 17256 22272 17262 22336
rect 16946 22271 17262 22272
rect 21946 22336 22262 22337
rect 21946 22272 21952 22336
rect 22016 22272 22032 22336
rect 22096 22272 22112 22336
rect 22176 22272 22192 22336
rect 22256 22272 22262 22336
rect 21946 22271 22262 22272
rect 26946 22336 27262 22337
rect 26946 22272 26952 22336
rect 27016 22272 27032 22336
rect 27096 22272 27112 22336
rect 27176 22272 27192 22336
rect 27256 22272 27262 22336
rect 26946 22271 27262 22272
rect 31946 22336 32262 22337
rect 31946 22272 31952 22336
rect 32016 22272 32032 22336
rect 32096 22272 32112 22336
rect 32176 22272 32192 22336
rect 32256 22272 32262 22336
rect 31946 22271 32262 22272
rect 36946 22336 37262 22337
rect 36946 22272 36952 22336
rect 37016 22272 37032 22336
rect 37096 22272 37112 22336
rect 37176 22272 37192 22336
rect 37256 22272 37262 22336
rect 41200 22312 42000 22342
rect 36946 22271 37262 22272
rect 2606 21792 2922 21793
rect 2606 21728 2612 21792
rect 2676 21728 2692 21792
rect 2756 21728 2772 21792
rect 2836 21728 2852 21792
rect 2916 21728 2922 21792
rect 2606 21727 2922 21728
rect 7606 21792 7922 21793
rect 7606 21728 7612 21792
rect 7676 21728 7692 21792
rect 7756 21728 7772 21792
rect 7836 21728 7852 21792
rect 7916 21728 7922 21792
rect 7606 21727 7922 21728
rect 12606 21792 12922 21793
rect 12606 21728 12612 21792
rect 12676 21728 12692 21792
rect 12756 21728 12772 21792
rect 12836 21728 12852 21792
rect 12916 21728 12922 21792
rect 12606 21727 12922 21728
rect 17606 21792 17922 21793
rect 17606 21728 17612 21792
rect 17676 21728 17692 21792
rect 17756 21728 17772 21792
rect 17836 21728 17852 21792
rect 17916 21728 17922 21792
rect 17606 21727 17922 21728
rect 22606 21792 22922 21793
rect 22606 21728 22612 21792
rect 22676 21728 22692 21792
rect 22756 21728 22772 21792
rect 22836 21728 22852 21792
rect 22916 21728 22922 21792
rect 22606 21727 22922 21728
rect 27606 21792 27922 21793
rect 27606 21728 27612 21792
rect 27676 21728 27692 21792
rect 27756 21728 27772 21792
rect 27836 21728 27852 21792
rect 27916 21728 27922 21792
rect 27606 21727 27922 21728
rect 32606 21792 32922 21793
rect 32606 21728 32612 21792
rect 32676 21728 32692 21792
rect 32756 21728 32772 21792
rect 32836 21728 32852 21792
rect 32916 21728 32922 21792
rect 32606 21727 32922 21728
rect 37606 21792 37922 21793
rect 37606 21728 37612 21792
rect 37676 21728 37692 21792
rect 37756 21728 37772 21792
rect 37836 21728 37852 21792
rect 37916 21728 37922 21792
rect 37606 21727 37922 21728
rect 1946 21248 2262 21249
rect 1946 21184 1952 21248
rect 2016 21184 2032 21248
rect 2096 21184 2112 21248
rect 2176 21184 2192 21248
rect 2256 21184 2262 21248
rect 1946 21183 2262 21184
rect 6946 21248 7262 21249
rect 6946 21184 6952 21248
rect 7016 21184 7032 21248
rect 7096 21184 7112 21248
rect 7176 21184 7192 21248
rect 7256 21184 7262 21248
rect 6946 21183 7262 21184
rect 11946 21248 12262 21249
rect 11946 21184 11952 21248
rect 12016 21184 12032 21248
rect 12096 21184 12112 21248
rect 12176 21184 12192 21248
rect 12256 21184 12262 21248
rect 11946 21183 12262 21184
rect 16946 21248 17262 21249
rect 16946 21184 16952 21248
rect 17016 21184 17032 21248
rect 17096 21184 17112 21248
rect 17176 21184 17192 21248
rect 17256 21184 17262 21248
rect 16946 21183 17262 21184
rect 21946 21248 22262 21249
rect 21946 21184 21952 21248
rect 22016 21184 22032 21248
rect 22096 21184 22112 21248
rect 22176 21184 22192 21248
rect 22256 21184 22262 21248
rect 21946 21183 22262 21184
rect 26946 21248 27262 21249
rect 26946 21184 26952 21248
rect 27016 21184 27032 21248
rect 27096 21184 27112 21248
rect 27176 21184 27192 21248
rect 27256 21184 27262 21248
rect 26946 21183 27262 21184
rect 31946 21248 32262 21249
rect 31946 21184 31952 21248
rect 32016 21184 32032 21248
rect 32096 21184 32112 21248
rect 32176 21184 32192 21248
rect 32256 21184 32262 21248
rect 31946 21183 32262 21184
rect 36946 21248 37262 21249
rect 36946 21184 36952 21248
rect 37016 21184 37032 21248
rect 37096 21184 37112 21248
rect 37176 21184 37192 21248
rect 37256 21184 37262 21248
rect 36946 21183 37262 21184
rect 2606 20704 2922 20705
rect 2606 20640 2612 20704
rect 2676 20640 2692 20704
rect 2756 20640 2772 20704
rect 2836 20640 2852 20704
rect 2916 20640 2922 20704
rect 2606 20639 2922 20640
rect 7606 20704 7922 20705
rect 7606 20640 7612 20704
rect 7676 20640 7692 20704
rect 7756 20640 7772 20704
rect 7836 20640 7852 20704
rect 7916 20640 7922 20704
rect 7606 20639 7922 20640
rect 12606 20704 12922 20705
rect 12606 20640 12612 20704
rect 12676 20640 12692 20704
rect 12756 20640 12772 20704
rect 12836 20640 12852 20704
rect 12916 20640 12922 20704
rect 12606 20639 12922 20640
rect 17606 20704 17922 20705
rect 17606 20640 17612 20704
rect 17676 20640 17692 20704
rect 17756 20640 17772 20704
rect 17836 20640 17852 20704
rect 17916 20640 17922 20704
rect 17606 20639 17922 20640
rect 22606 20704 22922 20705
rect 22606 20640 22612 20704
rect 22676 20640 22692 20704
rect 22756 20640 22772 20704
rect 22836 20640 22852 20704
rect 22916 20640 22922 20704
rect 22606 20639 22922 20640
rect 27606 20704 27922 20705
rect 27606 20640 27612 20704
rect 27676 20640 27692 20704
rect 27756 20640 27772 20704
rect 27836 20640 27852 20704
rect 27916 20640 27922 20704
rect 27606 20639 27922 20640
rect 32606 20704 32922 20705
rect 32606 20640 32612 20704
rect 32676 20640 32692 20704
rect 32756 20640 32772 20704
rect 32836 20640 32852 20704
rect 32916 20640 32922 20704
rect 32606 20639 32922 20640
rect 37606 20704 37922 20705
rect 37606 20640 37612 20704
rect 37676 20640 37692 20704
rect 37756 20640 37772 20704
rect 37836 20640 37852 20704
rect 37916 20640 37922 20704
rect 37606 20639 37922 20640
rect 1946 20160 2262 20161
rect 1946 20096 1952 20160
rect 2016 20096 2032 20160
rect 2096 20096 2112 20160
rect 2176 20096 2192 20160
rect 2256 20096 2262 20160
rect 1946 20095 2262 20096
rect 6946 20160 7262 20161
rect 6946 20096 6952 20160
rect 7016 20096 7032 20160
rect 7096 20096 7112 20160
rect 7176 20096 7192 20160
rect 7256 20096 7262 20160
rect 6946 20095 7262 20096
rect 11946 20160 12262 20161
rect 11946 20096 11952 20160
rect 12016 20096 12032 20160
rect 12096 20096 12112 20160
rect 12176 20096 12192 20160
rect 12256 20096 12262 20160
rect 11946 20095 12262 20096
rect 16946 20160 17262 20161
rect 16946 20096 16952 20160
rect 17016 20096 17032 20160
rect 17096 20096 17112 20160
rect 17176 20096 17192 20160
rect 17256 20096 17262 20160
rect 16946 20095 17262 20096
rect 21946 20160 22262 20161
rect 21946 20096 21952 20160
rect 22016 20096 22032 20160
rect 22096 20096 22112 20160
rect 22176 20096 22192 20160
rect 22256 20096 22262 20160
rect 21946 20095 22262 20096
rect 26946 20160 27262 20161
rect 26946 20096 26952 20160
rect 27016 20096 27032 20160
rect 27096 20096 27112 20160
rect 27176 20096 27192 20160
rect 27256 20096 27262 20160
rect 26946 20095 27262 20096
rect 31946 20160 32262 20161
rect 31946 20096 31952 20160
rect 32016 20096 32032 20160
rect 32096 20096 32112 20160
rect 32176 20096 32192 20160
rect 32256 20096 32262 20160
rect 31946 20095 32262 20096
rect 36946 20160 37262 20161
rect 36946 20096 36952 20160
rect 37016 20096 37032 20160
rect 37096 20096 37112 20160
rect 37176 20096 37192 20160
rect 37256 20096 37262 20160
rect 36946 20095 37262 20096
rect 2606 19616 2922 19617
rect 2606 19552 2612 19616
rect 2676 19552 2692 19616
rect 2756 19552 2772 19616
rect 2836 19552 2852 19616
rect 2916 19552 2922 19616
rect 2606 19551 2922 19552
rect 7606 19616 7922 19617
rect 7606 19552 7612 19616
rect 7676 19552 7692 19616
rect 7756 19552 7772 19616
rect 7836 19552 7852 19616
rect 7916 19552 7922 19616
rect 7606 19551 7922 19552
rect 12606 19616 12922 19617
rect 12606 19552 12612 19616
rect 12676 19552 12692 19616
rect 12756 19552 12772 19616
rect 12836 19552 12852 19616
rect 12916 19552 12922 19616
rect 12606 19551 12922 19552
rect 17606 19616 17922 19617
rect 17606 19552 17612 19616
rect 17676 19552 17692 19616
rect 17756 19552 17772 19616
rect 17836 19552 17852 19616
rect 17916 19552 17922 19616
rect 17606 19551 17922 19552
rect 22606 19616 22922 19617
rect 22606 19552 22612 19616
rect 22676 19552 22692 19616
rect 22756 19552 22772 19616
rect 22836 19552 22852 19616
rect 22916 19552 22922 19616
rect 22606 19551 22922 19552
rect 27606 19616 27922 19617
rect 27606 19552 27612 19616
rect 27676 19552 27692 19616
rect 27756 19552 27772 19616
rect 27836 19552 27852 19616
rect 27916 19552 27922 19616
rect 27606 19551 27922 19552
rect 32606 19616 32922 19617
rect 32606 19552 32612 19616
rect 32676 19552 32692 19616
rect 32756 19552 32772 19616
rect 32836 19552 32852 19616
rect 32916 19552 32922 19616
rect 32606 19551 32922 19552
rect 37606 19616 37922 19617
rect 37606 19552 37612 19616
rect 37676 19552 37692 19616
rect 37756 19552 37772 19616
rect 37836 19552 37852 19616
rect 37916 19552 37922 19616
rect 37606 19551 37922 19552
rect 1946 19072 2262 19073
rect 1946 19008 1952 19072
rect 2016 19008 2032 19072
rect 2096 19008 2112 19072
rect 2176 19008 2192 19072
rect 2256 19008 2262 19072
rect 1946 19007 2262 19008
rect 6946 19072 7262 19073
rect 6946 19008 6952 19072
rect 7016 19008 7032 19072
rect 7096 19008 7112 19072
rect 7176 19008 7192 19072
rect 7256 19008 7262 19072
rect 6946 19007 7262 19008
rect 11946 19072 12262 19073
rect 11946 19008 11952 19072
rect 12016 19008 12032 19072
rect 12096 19008 12112 19072
rect 12176 19008 12192 19072
rect 12256 19008 12262 19072
rect 11946 19007 12262 19008
rect 16946 19072 17262 19073
rect 16946 19008 16952 19072
rect 17016 19008 17032 19072
rect 17096 19008 17112 19072
rect 17176 19008 17192 19072
rect 17256 19008 17262 19072
rect 16946 19007 17262 19008
rect 21946 19072 22262 19073
rect 21946 19008 21952 19072
rect 22016 19008 22032 19072
rect 22096 19008 22112 19072
rect 22176 19008 22192 19072
rect 22256 19008 22262 19072
rect 21946 19007 22262 19008
rect 26946 19072 27262 19073
rect 26946 19008 26952 19072
rect 27016 19008 27032 19072
rect 27096 19008 27112 19072
rect 27176 19008 27192 19072
rect 27256 19008 27262 19072
rect 26946 19007 27262 19008
rect 31946 19072 32262 19073
rect 31946 19008 31952 19072
rect 32016 19008 32032 19072
rect 32096 19008 32112 19072
rect 32176 19008 32192 19072
rect 32256 19008 32262 19072
rect 31946 19007 32262 19008
rect 36946 19072 37262 19073
rect 36946 19008 36952 19072
rect 37016 19008 37032 19072
rect 37096 19008 37112 19072
rect 37176 19008 37192 19072
rect 37256 19008 37262 19072
rect 36946 19007 37262 19008
rect 2606 18528 2922 18529
rect 2606 18464 2612 18528
rect 2676 18464 2692 18528
rect 2756 18464 2772 18528
rect 2836 18464 2852 18528
rect 2916 18464 2922 18528
rect 2606 18463 2922 18464
rect 7606 18528 7922 18529
rect 7606 18464 7612 18528
rect 7676 18464 7692 18528
rect 7756 18464 7772 18528
rect 7836 18464 7852 18528
rect 7916 18464 7922 18528
rect 7606 18463 7922 18464
rect 12606 18528 12922 18529
rect 12606 18464 12612 18528
rect 12676 18464 12692 18528
rect 12756 18464 12772 18528
rect 12836 18464 12852 18528
rect 12916 18464 12922 18528
rect 12606 18463 12922 18464
rect 17606 18528 17922 18529
rect 17606 18464 17612 18528
rect 17676 18464 17692 18528
rect 17756 18464 17772 18528
rect 17836 18464 17852 18528
rect 17916 18464 17922 18528
rect 17606 18463 17922 18464
rect 22606 18528 22922 18529
rect 22606 18464 22612 18528
rect 22676 18464 22692 18528
rect 22756 18464 22772 18528
rect 22836 18464 22852 18528
rect 22916 18464 22922 18528
rect 22606 18463 22922 18464
rect 27606 18528 27922 18529
rect 27606 18464 27612 18528
rect 27676 18464 27692 18528
rect 27756 18464 27772 18528
rect 27836 18464 27852 18528
rect 27916 18464 27922 18528
rect 27606 18463 27922 18464
rect 32606 18528 32922 18529
rect 32606 18464 32612 18528
rect 32676 18464 32692 18528
rect 32756 18464 32772 18528
rect 32836 18464 32852 18528
rect 32916 18464 32922 18528
rect 32606 18463 32922 18464
rect 37606 18528 37922 18529
rect 37606 18464 37612 18528
rect 37676 18464 37692 18528
rect 37756 18464 37772 18528
rect 37836 18464 37852 18528
rect 37916 18464 37922 18528
rect 37606 18463 37922 18464
rect 1946 17984 2262 17985
rect 1946 17920 1952 17984
rect 2016 17920 2032 17984
rect 2096 17920 2112 17984
rect 2176 17920 2192 17984
rect 2256 17920 2262 17984
rect 1946 17919 2262 17920
rect 6946 17984 7262 17985
rect 6946 17920 6952 17984
rect 7016 17920 7032 17984
rect 7096 17920 7112 17984
rect 7176 17920 7192 17984
rect 7256 17920 7262 17984
rect 6946 17919 7262 17920
rect 11946 17984 12262 17985
rect 11946 17920 11952 17984
rect 12016 17920 12032 17984
rect 12096 17920 12112 17984
rect 12176 17920 12192 17984
rect 12256 17920 12262 17984
rect 11946 17919 12262 17920
rect 16946 17984 17262 17985
rect 16946 17920 16952 17984
rect 17016 17920 17032 17984
rect 17096 17920 17112 17984
rect 17176 17920 17192 17984
rect 17256 17920 17262 17984
rect 16946 17919 17262 17920
rect 21946 17984 22262 17985
rect 21946 17920 21952 17984
rect 22016 17920 22032 17984
rect 22096 17920 22112 17984
rect 22176 17920 22192 17984
rect 22256 17920 22262 17984
rect 21946 17919 22262 17920
rect 26946 17984 27262 17985
rect 26946 17920 26952 17984
rect 27016 17920 27032 17984
rect 27096 17920 27112 17984
rect 27176 17920 27192 17984
rect 27256 17920 27262 17984
rect 26946 17919 27262 17920
rect 31946 17984 32262 17985
rect 31946 17920 31952 17984
rect 32016 17920 32032 17984
rect 32096 17920 32112 17984
rect 32176 17920 32192 17984
rect 32256 17920 32262 17984
rect 31946 17919 32262 17920
rect 36946 17984 37262 17985
rect 36946 17920 36952 17984
rect 37016 17920 37032 17984
rect 37096 17920 37112 17984
rect 37176 17920 37192 17984
rect 37256 17920 37262 17984
rect 36946 17919 37262 17920
rect 2606 17440 2922 17441
rect 2606 17376 2612 17440
rect 2676 17376 2692 17440
rect 2756 17376 2772 17440
rect 2836 17376 2852 17440
rect 2916 17376 2922 17440
rect 2606 17375 2922 17376
rect 7606 17440 7922 17441
rect 7606 17376 7612 17440
rect 7676 17376 7692 17440
rect 7756 17376 7772 17440
rect 7836 17376 7852 17440
rect 7916 17376 7922 17440
rect 7606 17375 7922 17376
rect 12606 17440 12922 17441
rect 12606 17376 12612 17440
rect 12676 17376 12692 17440
rect 12756 17376 12772 17440
rect 12836 17376 12852 17440
rect 12916 17376 12922 17440
rect 12606 17375 12922 17376
rect 17606 17440 17922 17441
rect 17606 17376 17612 17440
rect 17676 17376 17692 17440
rect 17756 17376 17772 17440
rect 17836 17376 17852 17440
rect 17916 17376 17922 17440
rect 17606 17375 17922 17376
rect 22606 17440 22922 17441
rect 22606 17376 22612 17440
rect 22676 17376 22692 17440
rect 22756 17376 22772 17440
rect 22836 17376 22852 17440
rect 22916 17376 22922 17440
rect 22606 17375 22922 17376
rect 27606 17440 27922 17441
rect 27606 17376 27612 17440
rect 27676 17376 27692 17440
rect 27756 17376 27772 17440
rect 27836 17376 27852 17440
rect 27916 17376 27922 17440
rect 27606 17375 27922 17376
rect 32606 17440 32922 17441
rect 32606 17376 32612 17440
rect 32676 17376 32692 17440
rect 32756 17376 32772 17440
rect 32836 17376 32852 17440
rect 32916 17376 32922 17440
rect 32606 17375 32922 17376
rect 37606 17440 37922 17441
rect 37606 17376 37612 17440
rect 37676 17376 37692 17440
rect 37756 17376 37772 17440
rect 37836 17376 37852 17440
rect 37916 17376 37922 17440
rect 37606 17375 37922 17376
rect 1946 16896 2262 16897
rect 1946 16832 1952 16896
rect 2016 16832 2032 16896
rect 2096 16832 2112 16896
rect 2176 16832 2192 16896
rect 2256 16832 2262 16896
rect 1946 16831 2262 16832
rect 6946 16896 7262 16897
rect 6946 16832 6952 16896
rect 7016 16832 7032 16896
rect 7096 16832 7112 16896
rect 7176 16832 7192 16896
rect 7256 16832 7262 16896
rect 6946 16831 7262 16832
rect 11946 16896 12262 16897
rect 11946 16832 11952 16896
rect 12016 16832 12032 16896
rect 12096 16832 12112 16896
rect 12176 16832 12192 16896
rect 12256 16832 12262 16896
rect 11946 16831 12262 16832
rect 16946 16896 17262 16897
rect 16946 16832 16952 16896
rect 17016 16832 17032 16896
rect 17096 16832 17112 16896
rect 17176 16832 17192 16896
rect 17256 16832 17262 16896
rect 16946 16831 17262 16832
rect 21946 16896 22262 16897
rect 21946 16832 21952 16896
rect 22016 16832 22032 16896
rect 22096 16832 22112 16896
rect 22176 16832 22192 16896
rect 22256 16832 22262 16896
rect 21946 16831 22262 16832
rect 26946 16896 27262 16897
rect 26946 16832 26952 16896
rect 27016 16832 27032 16896
rect 27096 16832 27112 16896
rect 27176 16832 27192 16896
rect 27256 16832 27262 16896
rect 26946 16831 27262 16832
rect 31946 16896 32262 16897
rect 31946 16832 31952 16896
rect 32016 16832 32032 16896
rect 32096 16832 32112 16896
rect 32176 16832 32192 16896
rect 32256 16832 32262 16896
rect 31946 16831 32262 16832
rect 36946 16896 37262 16897
rect 36946 16832 36952 16896
rect 37016 16832 37032 16896
rect 37096 16832 37112 16896
rect 37176 16832 37192 16896
rect 37256 16832 37262 16896
rect 36946 16831 37262 16832
rect 2606 16352 2922 16353
rect 2606 16288 2612 16352
rect 2676 16288 2692 16352
rect 2756 16288 2772 16352
rect 2836 16288 2852 16352
rect 2916 16288 2922 16352
rect 2606 16287 2922 16288
rect 7606 16352 7922 16353
rect 7606 16288 7612 16352
rect 7676 16288 7692 16352
rect 7756 16288 7772 16352
rect 7836 16288 7852 16352
rect 7916 16288 7922 16352
rect 7606 16287 7922 16288
rect 12606 16352 12922 16353
rect 12606 16288 12612 16352
rect 12676 16288 12692 16352
rect 12756 16288 12772 16352
rect 12836 16288 12852 16352
rect 12916 16288 12922 16352
rect 12606 16287 12922 16288
rect 17606 16352 17922 16353
rect 17606 16288 17612 16352
rect 17676 16288 17692 16352
rect 17756 16288 17772 16352
rect 17836 16288 17852 16352
rect 17916 16288 17922 16352
rect 17606 16287 17922 16288
rect 22606 16352 22922 16353
rect 22606 16288 22612 16352
rect 22676 16288 22692 16352
rect 22756 16288 22772 16352
rect 22836 16288 22852 16352
rect 22916 16288 22922 16352
rect 22606 16287 22922 16288
rect 27606 16352 27922 16353
rect 27606 16288 27612 16352
rect 27676 16288 27692 16352
rect 27756 16288 27772 16352
rect 27836 16288 27852 16352
rect 27916 16288 27922 16352
rect 27606 16287 27922 16288
rect 32606 16352 32922 16353
rect 32606 16288 32612 16352
rect 32676 16288 32692 16352
rect 32756 16288 32772 16352
rect 32836 16288 32852 16352
rect 32916 16288 32922 16352
rect 32606 16287 32922 16288
rect 37606 16352 37922 16353
rect 37606 16288 37612 16352
rect 37676 16288 37692 16352
rect 37756 16288 37772 16352
rect 37836 16288 37852 16352
rect 37916 16288 37922 16352
rect 37606 16287 37922 16288
rect 1946 15808 2262 15809
rect 1946 15744 1952 15808
rect 2016 15744 2032 15808
rect 2096 15744 2112 15808
rect 2176 15744 2192 15808
rect 2256 15744 2262 15808
rect 1946 15743 2262 15744
rect 6946 15808 7262 15809
rect 6946 15744 6952 15808
rect 7016 15744 7032 15808
rect 7096 15744 7112 15808
rect 7176 15744 7192 15808
rect 7256 15744 7262 15808
rect 6946 15743 7262 15744
rect 11946 15808 12262 15809
rect 11946 15744 11952 15808
rect 12016 15744 12032 15808
rect 12096 15744 12112 15808
rect 12176 15744 12192 15808
rect 12256 15744 12262 15808
rect 11946 15743 12262 15744
rect 16946 15808 17262 15809
rect 16946 15744 16952 15808
rect 17016 15744 17032 15808
rect 17096 15744 17112 15808
rect 17176 15744 17192 15808
rect 17256 15744 17262 15808
rect 16946 15743 17262 15744
rect 21946 15808 22262 15809
rect 21946 15744 21952 15808
rect 22016 15744 22032 15808
rect 22096 15744 22112 15808
rect 22176 15744 22192 15808
rect 22256 15744 22262 15808
rect 21946 15743 22262 15744
rect 26946 15808 27262 15809
rect 26946 15744 26952 15808
rect 27016 15744 27032 15808
rect 27096 15744 27112 15808
rect 27176 15744 27192 15808
rect 27256 15744 27262 15808
rect 26946 15743 27262 15744
rect 31946 15808 32262 15809
rect 31946 15744 31952 15808
rect 32016 15744 32032 15808
rect 32096 15744 32112 15808
rect 32176 15744 32192 15808
rect 32256 15744 32262 15808
rect 31946 15743 32262 15744
rect 36946 15808 37262 15809
rect 36946 15744 36952 15808
rect 37016 15744 37032 15808
rect 37096 15744 37112 15808
rect 37176 15744 37192 15808
rect 37256 15744 37262 15808
rect 36946 15743 37262 15744
rect 2606 15264 2922 15265
rect 2606 15200 2612 15264
rect 2676 15200 2692 15264
rect 2756 15200 2772 15264
rect 2836 15200 2852 15264
rect 2916 15200 2922 15264
rect 2606 15199 2922 15200
rect 7606 15264 7922 15265
rect 7606 15200 7612 15264
rect 7676 15200 7692 15264
rect 7756 15200 7772 15264
rect 7836 15200 7852 15264
rect 7916 15200 7922 15264
rect 7606 15199 7922 15200
rect 12606 15264 12922 15265
rect 12606 15200 12612 15264
rect 12676 15200 12692 15264
rect 12756 15200 12772 15264
rect 12836 15200 12852 15264
rect 12916 15200 12922 15264
rect 12606 15199 12922 15200
rect 17606 15264 17922 15265
rect 17606 15200 17612 15264
rect 17676 15200 17692 15264
rect 17756 15200 17772 15264
rect 17836 15200 17852 15264
rect 17916 15200 17922 15264
rect 17606 15199 17922 15200
rect 22606 15264 22922 15265
rect 22606 15200 22612 15264
rect 22676 15200 22692 15264
rect 22756 15200 22772 15264
rect 22836 15200 22852 15264
rect 22916 15200 22922 15264
rect 22606 15199 22922 15200
rect 27606 15264 27922 15265
rect 27606 15200 27612 15264
rect 27676 15200 27692 15264
rect 27756 15200 27772 15264
rect 27836 15200 27852 15264
rect 27916 15200 27922 15264
rect 27606 15199 27922 15200
rect 32606 15264 32922 15265
rect 32606 15200 32612 15264
rect 32676 15200 32692 15264
rect 32756 15200 32772 15264
rect 32836 15200 32852 15264
rect 32916 15200 32922 15264
rect 32606 15199 32922 15200
rect 37606 15264 37922 15265
rect 37606 15200 37612 15264
rect 37676 15200 37692 15264
rect 37756 15200 37772 15264
rect 37836 15200 37852 15264
rect 37916 15200 37922 15264
rect 37606 15199 37922 15200
rect 22369 15058 22435 15061
rect 24894 15058 24900 15060
rect 22369 15056 24900 15058
rect 22369 15000 22374 15056
rect 22430 15000 24900 15056
rect 22369 14998 24900 15000
rect 22369 14995 22435 14998
rect 24894 14996 24900 14998
rect 24964 15058 24970 15060
rect 35341 15058 35407 15061
rect 24964 15056 35407 15058
rect 24964 15000 35346 15056
rect 35402 15000 35407 15056
rect 24964 14998 35407 15000
rect 24964 14996 24970 14998
rect 35341 14995 35407 14998
rect 1946 14720 2262 14721
rect 1946 14656 1952 14720
rect 2016 14656 2032 14720
rect 2096 14656 2112 14720
rect 2176 14656 2192 14720
rect 2256 14656 2262 14720
rect 1946 14655 2262 14656
rect 6946 14720 7262 14721
rect 6946 14656 6952 14720
rect 7016 14656 7032 14720
rect 7096 14656 7112 14720
rect 7176 14656 7192 14720
rect 7256 14656 7262 14720
rect 6946 14655 7262 14656
rect 11946 14720 12262 14721
rect 11946 14656 11952 14720
rect 12016 14656 12032 14720
rect 12096 14656 12112 14720
rect 12176 14656 12192 14720
rect 12256 14656 12262 14720
rect 11946 14655 12262 14656
rect 16946 14720 17262 14721
rect 16946 14656 16952 14720
rect 17016 14656 17032 14720
rect 17096 14656 17112 14720
rect 17176 14656 17192 14720
rect 17256 14656 17262 14720
rect 16946 14655 17262 14656
rect 21946 14720 22262 14721
rect 21946 14656 21952 14720
rect 22016 14656 22032 14720
rect 22096 14656 22112 14720
rect 22176 14656 22192 14720
rect 22256 14656 22262 14720
rect 21946 14655 22262 14656
rect 26946 14720 27262 14721
rect 26946 14656 26952 14720
rect 27016 14656 27032 14720
rect 27096 14656 27112 14720
rect 27176 14656 27192 14720
rect 27256 14656 27262 14720
rect 26946 14655 27262 14656
rect 31946 14720 32262 14721
rect 31946 14656 31952 14720
rect 32016 14656 32032 14720
rect 32096 14656 32112 14720
rect 32176 14656 32192 14720
rect 32256 14656 32262 14720
rect 31946 14655 32262 14656
rect 36946 14720 37262 14721
rect 36946 14656 36952 14720
rect 37016 14656 37032 14720
rect 37096 14656 37112 14720
rect 37176 14656 37192 14720
rect 37256 14656 37262 14720
rect 36946 14655 37262 14656
rect 2606 14176 2922 14177
rect 2606 14112 2612 14176
rect 2676 14112 2692 14176
rect 2756 14112 2772 14176
rect 2836 14112 2852 14176
rect 2916 14112 2922 14176
rect 2606 14111 2922 14112
rect 7606 14176 7922 14177
rect 7606 14112 7612 14176
rect 7676 14112 7692 14176
rect 7756 14112 7772 14176
rect 7836 14112 7852 14176
rect 7916 14112 7922 14176
rect 7606 14111 7922 14112
rect 12606 14176 12922 14177
rect 12606 14112 12612 14176
rect 12676 14112 12692 14176
rect 12756 14112 12772 14176
rect 12836 14112 12852 14176
rect 12916 14112 12922 14176
rect 12606 14111 12922 14112
rect 17606 14176 17922 14177
rect 17606 14112 17612 14176
rect 17676 14112 17692 14176
rect 17756 14112 17772 14176
rect 17836 14112 17852 14176
rect 17916 14112 17922 14176
rect 17606 14111 17922 14112
rect 22606 14176 22922 14177
rect 22606 14112 22612 14176
rect 22676 14112 22692 14176
rect 22756 14112 22772 14176
rect 22836 14112 22852 14176
rect 22916 14112 22922 14176
rect 22606 14111 22922 14112
rect 27606 14176 27922 14177
rect 27606 14112 27612 14176
rect 27676 14112 27692 14176
rect 27756 14112 27772 14176
rect 27836 14112 27852 14176
rect 27916 14112 27922 14176
rect 27606 14111 27922 14112
rect 32606 14176 32922 14177
rect 32606 14112 32612 14176
rect 32676 14112 32692 14176
rect 32756 14112 32772 14176
rect 32836 14112 32852 14176
rect 32916 14112 32922 14176
rect 32606 14111 32922 14112
rect 37606 14176 37922 14177
rect 37606 14112 37612 14176
rect 37676 14112 37692 14176
rect 37756 14112 37772 14176
rect 37836 14112 37852 14176
rect 37916 14112 37922 14176
rect 37606 14111 37922 14112
rect 1946 13632 2262 13633
rect 1946 13568 1952 13632
rect 2016 13568 2032 13632
rect 2096 13568 2112 13632
rect 2176 13568 2192 13632
rect 2256 13568 2262 13632
rect 1946 13567 2262 13568
rect 6946 13632 7262 13633
rect 6946 13568 6952 13632
rect 7016 13568 7032 13632
rect 7096 13568 7112 13632
rect 7176 13568 7192 13632
rect 7256 13568 7262 13632
rect 6946 13567 7262 13568
rect 11946 13632 12262 13633
rect 11946 13568 11952 13632
rect 12016 13568 12032 13632
rect 12096 13568 12112 13632
rect 12176 13568 12192 13632
rect 12256 13568 12262 13632
rect 11946 13567 12262 13568
rect 16946 13632 17262 13633
rect 16946 13568 16952 13632
rect 17016 13568 17032 13632
rect 17096 13568 17112 13632
rect 17176 13568 17192 13632
rect 17256 13568 17262 13632
rect 16946 13567 17262 13568
rect 21946 13632 22262 13633
rect 21946 13568 21952 13632
rect 22016 13568 22032 13632
rect 22096 13568 22112 13632
rect 22176 13568 22192 13632
rect 22256 13568 22262 13632
rect 21946 13567 22262 13568
rect 26946 13632 27262 13633
rect 26946 13568 26952 13632
rect 27016 13568 27032 13632
rect 27096 13568 27112 13632
rect 27176 13568 27192 13632
rect 27256 13568 27262 13632
rect 26946 13567 27262 13568
rect 31946 13632 32262 13633
rect 31946 13568 31952 13632
rect 32016 13568 32032 13632
rect 32096 13568 32112 13632
rect 32176 13568 32192 13632
rect 32256 13568 32262 13632
rect 31946 13567 32262 13568
rect 36946 13632 37262 13633
rect 36946 13568 36952 13632
rect 37016 13568 37032 13632
rect 37096 13568 37112 13632
rect 37176 13568 37192 13632
rect 37256 13568 37262 13632
rect 36946 13567 37262 13568
rect 0 13426 800 13456
rect 1393 13426 1459 13429
rect 0 13424 1459 13426
rect 0 13368 1398 13424
rect 1454 13368 1459 13424
rect 0 13366 1459 13368
rect 0 13336 800 13366
rect 1393 13363 1459 13366
rect 16573 13426 16639 13429
rect 21582 13426 21588 13428
rect 16573 13424 21588 13426
rect 16573 13368 16578 13424
rect 16634 13368 21588 13424
rect 16573 13366 21588 13368
rect 16573 13363 16639 13366
rect 21582 13364 21588 13366
rect 21652 13364 21658 13428
rect 39941 13426 40007 13429
rect 41200 13426 42000 13456
rect 39941 13424 42000 13426
rect 39941 13368 39946 13424
rect 40002 13368 42000 13424
rect 39941 13366 42000 13368
rect 39941 13363 40007 13366
rect 41200 13336 42000 13366
rect 2606 13088 2922 13089
rect 2606 13024 2612 13088
rect 2676 13024 2692 13088
rect 2756 13024 2772 13088
rect 2836 13024 2852 13088
rect 2916 13024 2922 13088
rect 2606 13023 2922 13024
rect 7606 13088 7922 13089
rect 7606 13024 7612 13088
rect 7676 13024 7692 13088
rect 7756 13024 7772 13088
rect 7836 13024 7852 13088
rect 7916 13024 7922 13088
rect 7606 13023 7922 13024
rect 12606 13088 12922 13089
rect 12606 13024 12612 13088
rect 12676 13024 12692 13088
rect 12756 13024 12772 13088
rect 12836 13024 12852 13088
rect 12916 13024 12922 13088
rect 12606 13023 12922 13024
rect 17606 13088 17922 13089
rect 17606 13024 17612 13088
rect 17676 13024 17692 13088
rect 17756 13024 17772 13088
rect 17836 13024 17852 13088
rect 17916 13024 17922 13088
rect 17606 13023 17922 13024
rect 22606 13088 22922 13089
rect 22606 13024 22612 13088
rect 22676 13024 22692 13088
rect 22756 13024 22772 13088
rect 22836 13024 22852 13088
rect 22916 13024 22922 13088
rect 22606 13023 22922 13024
rect 27606 13088 27922 13089
rect 27606 13024 27612 13088
rect 27676 13024 27692 13088
rect 27756 13024 27772 13088
rect 27836 13024 27852 13088
rect 27916 13024 27922 13088
rect 27606 13023 27922 13024
rect 32606 13088 32922 13089
rect 32606 13024 32612 13088
rect 32676 13024 32692 13088
rect 32756 13024 32772 13088
rect 32836 13024 32852 13088
rect 32916 13024 32922 13088
rect 32606 13023 32922 13024
rect 37606 13088 37922 13089
rect 37606 13024 37612 13088
rect 37676 13024 37692 13088
rect 37756 13024 37772 13088
rect 37836 13024 37852 13088
rect 37916 13024 37922 13088
rect 37606 13023 37922 13024
rect 1946 12544 2262 12545
rect 1946 12480 1952 12544
rect 2016 12480 2032 12544
rect 2096 12480 2112 12544
rect 2176 12480 2192 12544
rect 2256 12480 2262 12544
rect 1946 12479 2262 12480
rect 6946 12544 7262 12545
rect 6946 12480 6952 12544
rect 7016 12480 7032 12544
rect 7096 12480 7112 12544
rect 7176 12480 7192 12544
rect 7256 12480 7262 12544
rect 6946 12479 7262 12480
rect 11946 12544 12262 12545
rect 11946 12480 11952 12544
rect 12016 12480 12032 12544
rect 12096 12480 12112 12544
rect 12176 12480 12192 12544
rect 12256 12480 12262 12544
rect 11946 12479 12262 12480
rect 16946 12544 17262 12545
rect 16946 12480 16952 12544
rect 17016 12480 17032 12544
rect 17096 12480 17112 12544
rect 17176 12480 17192 12544
rect 17256 12480 17262 12544
rect 16946 12479 17262 12480
rect 21946 12544 22262 12545
rect 21946 12480 21952 12544
rect 22016 12480 22032 12544
rect 22096 12480 22112 12544
rect 22176 12480 22192 12544
rect 22256 12480 22262 12544
rect 21946 12479 22262 12480
rect 26946 12544 27262 12545
rect 26946 12480 26952 12544
rect 27016 12480 27032 12544
rect 27096 12480 27112 12544
rect 27176 12480 27192 12544
rect 27256 12480 27262 12544
rect 26946 12479 27262 12480
rect 31946 12544 32262 12545
rect 31946 12480 31952 12544
rect 32016 12480 32032 12544
rect 32096 12480 32112 12544
rect 32176 12480 32192 12544
rect 32256 12480 32262 12544
rect 31946 12479 32262 12480
rect 36946 12544 37262 12545
rect 36946 12480 36952 12544
rect 37016 12480 37032 12544
rect 37096 12480 37112 12544
rect 37176 12480 37192 12544
rect 37256 12480 37262 12544
rect 36946 12479 37262 12480
rect 20478 12140 20484 12204
rect 20548 12202 20554 12204
rect 24853 12202 24919 12205
rect 20548 12200 24919 12202
rect 20548 12144 24858 12200
rect 24914 12144 24919 12200
rect 20548 12142 24919 12144
rect 20548 12140 20554 12142
rect 24853 12139 24919 12142
rect 2606 12000 2922 12001
rect 2606 11936 2612 12000
rect 2676 11936 2692 12000
rect 2756 11936 2772 12000
rect 2836 11936 2852 12000
rect 2916 11936 2922 12000
rect 2606 11935 2922 11936
rect 7606 12000 7922 12001
rect 7606 11936 7612 12000
rect 7676 11936 7692 12000
rect 7756 11936 7772 12000
rect 7836 11936 7852 12000
rect 7916 11936 7922 12000
rect 7606 11935 7922 11936
rect 12606 12000 12922 12001
rect 12606 11936 12612 12000
rect 12676 11936 12692 12000
rect 12756 11936 12772 12000
rect 12836 11936 12852 12000
rect 12916 11936 12922 12000
rect 12606 11935 12922 11936
rect 17606 12000 17922 12001
rect 17606 11936 17612 12000
rect 17676 11936 17692 12000
rect 17756 11936 17772 12000
rect 17836 11936 17852 12000
rect 17916 11936 17922 12000
rect 17606 11935 17922 11936
rect 22606 12000 22922 12001
rect 22606 11936 22612 12000
rect 22676 11936 22692 12000
rect 22756 11936 22772 12000
rect 22836 11936 22852 12000
rect 22916 11936 22922 12000
rect 22606 11935 22922 11936
rect 27606 12000 27922 12001
rect 27606 11936 27612 12000
rect 27676 11936 27692 12000
rect 27756 11936 27772 12000
rect 27836 11936 27852 12000
rect 27916 11936 27922 12000
rect 27606 11935 27922 11936
rect 32606 12000 32922 12001
rect 32606 11936 32612 12000
rect 32676 11936 32692 12000
rect 32756 11936 32772 12000
rect 32836 11936 32852 12000
rect 32916 11936 32922 12000
rect 32606 11935 32922 11936
rect 37606 12000 37922 12001
rect 37606 11936 37612 12000
rect 37676 11936 37692 12000
rect 37756 11936 37772 12000
rect 37836 11936 37852 12000
rect 37916 11936 37922 12000
rect 37606 11935 37922 11936
rect 3785 11658 3851 11661
rect 34830 11658 34836 11660
rect 3785 11656 34836 11658
rect 3785 11600 3790 11656
rect 3846 11600 34836 11656
rect 3785 11598 34836 11600
rect 3785 11595 3851 11598
rect 34830 11596 34836 11598
rect 34900 11596 34906 11660
rect 1946 11456 2262 11457
rect 1946 11392 1952 11456
rect 2016 11392 2032 11456
rect 2096 11392 2112 11456
rect 2176 11392 2192 11456
rect 2256 11392 2262 11456
rect 1946 11391 2262 11392
rect 6946 11456 7262 11457
rect 6946 11392 6952 11456
rect 7016 11392 7032 11456
rect 7096 11392 7112 11456
rect 7176 11392 7192 11456
rect 7256 11392 7262 11456
rect 6946 11391 7262 11392
rect 11946 11456 12262 11457
rect 11946 11392 11952 11456
rect 12016 11392 12032 11456
rect 12096 11392 12112 11456
rect 12176 11392 12192 11456
rect 12256 11392 12262 11456
rect 11946 11391 12262 11392
rect 16946 11456 17262 11457
rect 16946 11392 16952 11456
rect 17016 11392 17032 11456
rect 17096 11392 17112 11456
rect 17176 11392 17192 11456
rect 17256 11392 17262 11456
rect 16946 11391 17262 11392
rect 21946 11456 22262 11457
rect 21946 11392 21952 11456
rect 22016 11392 22032 11456
rect 22096 11392 22112 11456
rect 22176 11392 22192 11456
rect 22256 11392 22262 11456
rect 21946 11391 22262 11392
rect 26946 11456 27262 11457
rect 26946 11392 26952 11456
rect 27016 11392 27032 11456
rect 27096 11392 27112 11456
rect 27176 11392 27192 11456
rect 27256 11392 27262 11456
rect 26946 11391 27262 11392
rect 31946 11456 32262 11457
rect 31946 11392 31952 11456
rect 32016 11392 32032 11456
rect 32096 11392 32112 11456
rect 32176 11392 32192 11456
rect 32256 11392 32262 11456
rect 31946 11391 32262 11392
rect 36946 11456 37262 11457
rect 36946 11392 36952 11456
rect 37016 11392 37032 11456
rect 37096 11392 37112 11456
rect 37176 11392 37192 11456
rect 37256 11392 37262 11456
rect 36946 11391 37262 11392
rect 1853 11114 1919 11117
rect 3366 11114 3372 11116
rect 1853 11112 3372 11114
rect 1853 11056 1858 11112
rect 1914 11056 3372 11112
rect 1853 11054 3372 11056
rect 1853 11051 1919 11054
rect 3366 11052 3372 11054
rect 3436 11052 3442 11116
rect 2606 10912 2922 10913
rect 2606 10848 2612 10912
rect 2676 10848 2692 10912
rect 2756 10848 2772 10912
rect 2836 10848 2852 10912
rect 2916 10848 2922 10912
rect 2606 10847 2922 10848
rect 7606 10912 7922 10913
rect 7606 10848 7612 10912
rect 7676 10848 7692 10912
rect 7756 10848 7772 10912
rect 7836 10848 7852 10912
rect 7916 10848 7922 10912
rect 7606 10847 7922 10848
rect 12606 10912 12922 10913
rect 12606 10848 12612 10912
rect 12676 10848 12692 10912
rect 12756 10848 12772 10912
rect 12836 10848 12852 10912
rect 12916 10848 12922 10912
rect 12606 10847 12922 10848
rect 17606 10912 17922 10913
rect 17606 10848 17612 10912
rect 17676 10848 17692 10912
rect 17756 10848 17772 10912
rect 17836 10848 17852 10912
rect 17916 10848 17922 10912
rect 17606 10847 17922 10848
rect 22606 10912 22922 10913
rect 22606 10848 22612 10912
rect 22676 10848 22692 10912
rect 22756 10848 22772 10912
rect 22836 10848 22852 10912
rect 22916 10848 22922 10912
rect 22606 10847 22922 10848
rect 27606 10912 27922 10913
rect 27606 10848 27612 10912
rect 27676 10848 27692 10912
rect 27756 10848 27772 10912
rect 27836 10848 27852 10912
rect 27916 10848 27922 10912
rect 27606 10847 27922 10848
rect 32606 10912 32922 10913
rect 32606 10848 32612 10912
rect 32676 10848 32692 10912
rect 32756 10848 32772 10912
rect 32836 10848 32852 10912
rect 32916 10848 32922 10912
rect 32606 10847 32922 10848
rect 37606 10912 37922 10913
rect 37606 10848 37612 10912
rect 37676 10848 37692 10912
rect 37756 10848 37772 10912
rect 37836 10848 37852 10912
rect 37916 10848 37922 10912
rect 37606 10847 37922 10848
rect 1946 10368 2262 10369
rect 1946 10304 1952 10368
rect 2016 10304 2032 10368
rect 2096 10304 2112 10368
rect 2176 10304 2192 10368
rect 2256 10304 2262 10368
rect 1946 10303 2262 10304
rect 6946 10368 7262 10369
rect 6946 10304 6952 10368
rect 7016 10304 7032 10368
rect 7096 10304 7112 10368
rect 7176 10304 7192 10368
rect 7256 10304 7262 10368
rect 6946 10303 7262 10304
rect 11946 10368 12262 10369
rect 11946 10304 11952 10368
rect 12016 10304 12032 10368
rect 12096 10304 12112 10368
rect 12176 10304 12192 10368
rect 12256 10304 12262 10368
rect 11946 10303 12262 10304
rect 16946 10368 17262 10369
rect 16946 10304 16952 10368
rect 17016 10304 17032 10368
rect 17096 10304 17112 10368
rect 17176 10304 17192 10368
rect 17256 10304 17262 10368
rect 16946 10303 17262 10304
rect 21946 10368 22262 10369
rect 21946 10304 21952 10368
rect 22016 10304 22032 10368
rect 22096 10304 22112 10368
rect 22176 10304 22192 10368
rect 22256 10304 22262 10368
rect 21946 10303 22262 10304
rect 26946 10368 27262 10369
rect 26946 10304 26952 10368
rect 27016 10304 27032 10368
rect 27096 10304 27112 10368
rect 27176 10304 27192 10368
rect 27256 10304 27262 10368
rect 26946 10303 27262 10304
rect 31946 10368 32262 10369
rect 31946 10304 31952 10368
rect 32016 10304 32032 10368
rect 32096 10304 32112 10368
rect 32176 10304 32192 10368
rect 32256 10304 32262 10368
rect 31946 10303 32262 10304
rect 36946 10368 37262 10369
rect 36946 10304 36952 10368
rect 37016 10304 37032 10368
rect 37096 10304 37112 10368
rect 37176 10304 37192 10368
rect 37256 10304 37262 10368
rect 36946 10303 37262 10304
rect 2606 9824 2922 9825
rect 2606 9760 2612 9824
rect 2676 9760 2692 9824
rect 2756 9760 2772 9824
rect 2836 9760 2852 9824
rect 2916 9760 2922 9824
rect 2606 9759 2922 9760
rect 7606 9824 7922 9825
rect 7606 9760 7612 9824
rect 7676 9760 7692 9824
rect 7756 9760 7772 9824
rect 7836 9760 7852 9824
rect 7916 9760 7922 9824
rect 7606 9759 7922 9760
rect 12606 9824 12922 9825
rect 12606 9760 12612 9824
rect 12676 9760 12692 9824
rect 12756 9760 12772 9824
rect 12836 9760 12852 9824
rect 12916 9760 12922 9824
rect 12606 9759 12922 9760
rect 17606 9824 17922 9825
rect 17606 9760 17612 9824
rect 17676 9760 17692 9824
rect 17756 9760 17772 9824
rect 17836 9760 17852 9824
rect 17916 9760 17922 9824
rect 17606 9759 17922 9760
rect 22606 9824 22922 9825
rect 22606 9760 22612 9824
rect 22676 9760 22692 9824
rect 22756 9760 22772 9824
rect 22836 9760 22852 9824
rect 22916 9760 22922 9824
rect 22606 9759 22922 9760
rect 27606 9824 27922 9825
rect 27606 9760 27612 9824
rect 27676 9760 27692 9824
rect 27756 9760 27772 9824
rect 27836 9760 27852 9824
rect 27916 9760 27922 9824
rect 27606 9759 27922 9760
rect 32606 9824 32922 9825
rect 32606 9760 32612 9824
rect 32676 9760 32692 9824
rect 32756 9760 32772 9824
rect 32836 9760 32852 9824
rect 32916 9760 32922 9824
rect 32606 9759 32922 9760
rect 37606 9824 37922 9825
rect 37606 9760 37612 9824
rect 37676 9760 37692 9824
rect 37756 9760 37772 9824
rect 37836 9760 37852 9824
rect 37916 9760 37922 9824
rect 37606 9759 37922 9760
rect 1946 9280 2262 9281
rect 1946 9216 1952 9280
rect 2016 9216 2032 9280
rect 2096 9216 2112 9280
rect 2176 9216 2192 9280
rect 2256 9216 2262 9280
rect 1946 9215 2262 9216
rect 6946 9280 7262 9281
rect 6946 9216 6952 9280
rect 7016 9216 7032 9280
rect 7096 9216 7112 9280
rect 7176 9216 7192 9280
rect 7256 9216 7262 9280
rect 6946 9215 7262 9216
rect 11946 9280 12262 9281
rect 11946 9216 11952 9280
rect 12016 9216 12032 9280
rect 12096 9216 12112 9280
rect 12176 9216 12192 9280
rect 12256 9216 12262 9280
rect 11946 9215 12262 9216
rect 16946 9280 17262 9281
rect 16946 9216 16952 9280
rect 17016 9216 17032 9280
rect 17096 9216 17112 9280
rect 17176 9216 17192 9280
rect 17256 9216 17262 9280
rect 16946 9215 17262 9216
rect 21946 9280 22262 9281
rect 21946 9216 21952 9280
rect 22016 9216 22032 9280
rect 22096 9216 22112 9280
rect 22176 9216 22192 9280
rect 22256 9216 22262 9280
rect 21946 9215 22262 9216
rect 26946 9280 27262 9281
rect 26946 9216 26952 9280
rect 27016 9216 27032 9280
rect 27096 9216 27112 9280
rect 27176 9216 27192 9280
rect 27256 9216 27262 9280
rect 26946 9215 27262 9216
rect 31946 9280 32262 9281
rect 31946 9216 31952 9280
rect 32016 9216 32032 9280
rect 32096 9216 32112 9280
rect 32176 9216 32192 9280
rect 32256 9216 32262 9280
rect 31946 9215 32262 9216
rect 36946 9280 37262 9281
rect 36946 9216 36952 9280
rect 37016 9216 37032 9280
rect 37096 9216 37112 9280
rect 37176 9216 37192 9280
rect 37256 9216 37262 9280
rect 36946 9215 37262 9216
rect 2606 8736 2922 8737
rect 2606 8672 2612 8736
rect 2676 8672 2692 8736
rect 2756 8672 2772 8736
rect 2836 8672 2852 8736
rect 2916 8672 2922 8736
rect 2606 8671 2922 8672
rect 7606 8736 7922 8737
rect 7606 8672 7612 8736
rect 7676 8672 7692 8736
rect 7756 8672 7772 8736
rect 7836 8672 7852 8736
rect 7916 8672 7922 8736
rect 7606 8671 7922 8672
rect 12606 8736 12922 8737
rect 12606 8672 12612 8736
rect 12676 8672 12692 8736
rect 12756 8672 12772 8736
rect 12836 8672 12852 8736
rect 12916 8672 12922 8736
rect 12606 8671 12922 8672
rect 17606 8736 17922 8737
rect 17606 8672 17612 8736
rect 17676 8672 17692 8736
rect 17756 8672 17772 8736
rect 17836 8672 17852 8736
rect 17916 8672 17922 8736
rect 17606 8671 17922 8672
rect 22606 8736 22922 8737
rect 22606 8672 22612 8736
rect 22676 8672 22692 8736
rect 22756 8672 22772 8736
rect 22836 8672 22852 8736
rect 22916 8672 22922 8736
rect 22606 8671 22922 8672
rect 27606 8736 27922 8737
rect 27606 8672 27612 8736
rect 27676 8672 27692 8736
rect 27756 8672 27772 8736
rect 27836 8672 27852 8736
rect 27916 8672 27922 8736
rect 27606 8671 27922 8672
rect 32606 8736 32922 8737
rect 32606 8672 32612 8736
rect 32676 8672 32692 8736
rect 32756 8672 32772 8736
rect 32836 8672 32852 8736
rect 32916 8672 32922 8736
rect 32606 8671 32922 8672
rect 37606 8736 37922 8737
rect 37606 8672 37612 8736
rect 37676 8672 37692 8736
rect 37756 8672 37772 8736
rect 37836 8672 37852 8736
rect 37916 8672 37922 8736
rect 37606 8671 37922 8672
rect 1946 8192 2262 8193
rect 1946 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2262 8192
rect 1946 8127 2262 8128
rect 6946 8192 7262 8193
rect 6946 8128 6952 8192
rect 7016 8128 7032 8192
rect 7096 8128 7112 8192
rect 7176 8128 7192 8192
rect 7256 8128 7262 8192
rect 6946 8127 7262 8128
rect 11946 8192 12262 8193
rect 11946 8128 11952 8192
rect 12016 8128 12032 8192
rect 12096 8128 12112 8192
rect 12176 8128 12192 8192
rect 12256 8128 12262 8192
rect 11946 8127 12262 8128
rect 16946 8192 17262 8193
rect 16946 8128 16952 8192
rect 17016 8128 17032 8192
rect 17096 8128 17112 8192
rect 17176 8128 17192 8192
rect 17256 8128 17262 8192
rect 16946 8127 17262 8128
rect 21946 8192 22262 8193
rect 21946 8128 21952 8192
rect 22016 8128 22032 8192
rect 22096 8128 22112 8192
rect 22176 8128 22192 8192
rect 22256 8128 22262 8192
rect 21946 8127 22262 8128
rect 26946 8192 27262 8193
rect 26946 8128 26952 8192
rect 27016 8128 27032 8192
rect 27096 8128 27112 8192
rect 27176 8128 27192 8192
rect 27256 8128 27262 8192
rect 26946 8127 27262 8128
rect 31946 8192 32262 8193
rect 31946 8128 31952 8192
rect 32016 8128 32032 8192
rect 32096 8128 32112 8192
rect 32176 8128 32192 8192
rect 32256 8128 32262 8192
rect 31946 8127 32262 8128
rect 36946 8192 37262 8193
rect 36946 8128 36952 8192
rect 37016 8128 37032 8192
rect 37096 8128 37112 8192
rect 37176 8128 37192 8192
rect 37256 8128 37262 8192
rect 36946 8127 37262 8128
rect 2606 7648 2922 7649
rect 2606 7584 2612 7648
rect 2676 7584 2692 7648
rect 2756 7584 2772 7648
rect 2836 7584 2852 7648
rect 2916 7584 2922 7648
rect 2606 7583 2922 7584
rect 7606 7648 7922 7649
rect 7606 7584 7612 7648
rect 7676 7584 7692 7648
rect 7756 7584 7772 7648
rect 7836 7584 7852 7648
rect 7916 7584 7922 7648
rect 7606 7583 7922 7584
rect 12606 7648 12922 7649
rect 12606 7584 12612 7648
rect 12676 7584 12692 7648
rect 12756 7584 12772 7648
rect 12836 7584 12852 7648
rect 12916 7584 12922 7648
rect 12606 7583 12922 7584
rect 17606 7648 17922 7649
rect 17606 7584 17612 7648
rect 17676 7584 17692 7648
rect 17756 7584 17772 7648
rect 17836 7584 17852 7648
rect 17916 7584 17922 7648
rect 17606 7583 17922 7584
rect 22606 7648 22922 7649
rect 22606 7584 22612 7648
rect 22676 7584 22692 7648
rect 22756 7584 22772 7648
rect 22836 7584 22852 7648
rect 22916 7584 22922 7648
rect 22606 7583 22922 7584
rect 27606 7648 27922 7649
rect 27606 7584 27612 7648
rect 27676 7584 27692 7648
rect 27756 7584 27772 7648
rect 27836 7584 27852 7648
rect 27916 7584 27922 7648
rect 27606 7583 27922 7584
rect 32606 7648 32922 7649
rect 32606 7584 32612 7648
rect 32676 7584 32692 7648
rect 32756 7584 32772 7648
rect 32836 7584 32852 7648
rect 32916 7584 32922 7648
rect 32606 7583 32922 7584
rect 37606 7648 37922 7649
rect 37606 7584 37612 7648
rect 37676 7584 37692 7648
rect 37756 7584 37772 7648
rect 37836 7584 37852 7648
rect 37916 7584 37922 7648
rect 37606 7583 37922 7584
rect 1946 7104 2262 7105
rect 1946 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2262 7104
rect 1946 7039 2262 7040
rect 6946 7104 7262 7105
rect 6946 7040 6952 7104
rect 7016 7040 7032 7104
rect 7096 7040 7112 7104
rect 7176 7040 7192 7104
rect 7256 7040 7262 7104
rect 6946 7039 7262 7040
rect 11946 7104 12262 7105
rect 11946 7040 11952 7104
rect 12016 7040 12032 7104
rect 12096 7040 12112 7104
rect 12176 7040 12192 7104
rect 12256 7040 12262 7104
rect 11946 7039 12262 7040
rect 16946 7104 17262 7105
rect 16946 7040 16952 7104
rect 17016 7040 17032 7104
rect 17096 7040 17112 7104
rect 17176 7040 17192 7104
rect 17256 7040 17262 7104
rect 16946 7039 17262 7040
rect 21946 7104 22262 7105
rect 21946 7040 21952 7104
rect 22016 7040 22032 7104
rect 22096 7040 22112 7104
rect 22176 7040 22192 7104
rect 22256 7040 22262 7104
rect 21946 7039 22262 7040
rect 26946 7104 27262 7105
rect 26946 7040 26952 7104
rect 27016 7040 27032 7104
rect 27096 7040 27112 7104
rect 27176 7040 27192 7104
rect 27256 7040 27262 7104
rect 26946 7039 27262 7040
rect 31946 7104 32262 7105
rect 31946 7040 31952 7104
rect 32016 7040 32032 7104
rect 32096 7040 32112 7104
rect 32176 7040 32192 7104
rect 32256 7040 32262 7104
rect 31946 7039 32262 7040
rect 36946 7104 37262 7105
rect 36946 7040 36952 7104
rect 37016 7040 37032 7104
rect 37096 7040 37112 7104
rect 37176 7040 37192 7104
rect 37256 7040 37262 7104
rect 36946 7039 37262 7040
rect 2606 6560 2922 6561
rect 2606 6496 2612 6560
rect 2676 6496 2692 6560
rect 2756 6496 2772 6560
rect 2836 6496 2852 6560
rect 2916 6496 2922 6560
rect 2606 6495 2922 6496
rect 7606 6560 7922 6561
rect 7606 6496 7612 6560
rect 7676 6496 7692 6560
rect 7756 6496 7772 6560
rect 7836 6496 7852 6560
rect 7916 6496 7922 6560
rect 7606 6495 7922 6496
rect 12606 6560 12922 6561
rect 12606 6496 12612 6560
rect 12676 6496 12692 6560
rect 12756 6496 12772 6560
rect 12836 6496 12852 6560
rect 12916 6496 12922 6560
rect 12606 6495 12922 6496
rect 17606 6560 17922 6561
rect 17606 6496 17612 6560
rect 17676 6496 17692 6560
rect 17756 6496 17772 6560
rect 17836 6496 17852 6560
rect 17916 6496 17922 6560
rect 17606 6495 17922 6496
rect 22606 6560 22922 6561
rect 22606 6496 22612 6560
rect 22676 6496 22692 6560
rect 22756 6496 22772 6560
rect 22836 6496 22852 6560
rect 22916 6496 22922 6560
rect 22606 6495 22922 6496
rect 27606 6560 27922 6561
rect 27606 6496 27612 6560
rect 27676 6496 27692 6560
rect 27756 6496 27772 6560
rect 27836 6496 27852 6560
rect 27916 6496 27922 6560
rect 27606 6495 27922 6496
rect 32606 6560 32922 6561
rect 32606 6496 32612 6560
rect 32676 6496 32692 6560
rect 32756 6496 32772 6560
rect 32836 6496 32852 6560
rect 32916 6496 32922 6560
rect 32606 6495 32922 6496
rect 37606 6560 37922 6561
rect 37606 6496 37612 6560
rect 37676 6496 37692 6560
rect 37756 6496 37772 6560
rect 37836 6496 37852 6560
rect 37916 6496 37922 6560
rect 37606 6495 37922 6496
rect 1946 6016 2262 6017
rect 1946 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2262 6016
rect 1946 5951 2262 5952
rect 6946 6016 7262 6017
rect 6946 5952 6952 6016
rect 7016 5952 7032 6016
rect 7096 5952 7112 6016
rect 7176 5952 7192 6016
rect 7256 5952 7262 6016
rect 6946 5951 7262 5952
rect 11946 6016 12262 6017
rect 11946 5952 11952 6016
rect 12016 5952 12032 6016
rect 12096 5952 12112 6016
rect 12176 5952 12192 6016
rect 12256 5952 12262 6016
rect 11946 5951 12262 5952
rect 16946 6016 17262 6017
rect 16946 5952 16952 6016
rect 17016 5952 17032 6016
rect 17096 5952 17112 6016
rect 17176 5952 17192 6016
rect 17256 5952 17262 6016
rect 16946 5951 17262 5952
rect 21946 6016 22262 6017
rect 21946 5952 21952 6016
rect 22016 5952 22032 6016
rect 22096 5952 22112 6016
rect 22176 5952 22192 6016
rect 22256 5952 22262 6016
rect 21946 5951 22262 5952
rect 26946 6016 27262 6017
rect 26946 5952 26952 6016
rect 27016 5952 27032 6016
rect 27096 5952 27112 6016
rect 27176 5952 27192 6016
rect 27256 5952 27262 6016
rect 26946 5951 27262 5952
rect 31946 6016 32262 6017
rect 31946 5952 31952 6016
rect 32016 5952 32032 6016
rect 32096 5952 32112 6016
rect 32176 5952 32192 6016
rect 32256 5952 32262 6016
rect 31946 5951 32262 5952
rect 36946 6016 37262 6017
rect 36946 5952 36952 6016
rect 37016 5952 37032 6016
rect 37096 5952 37112 6016
rect 37176 5952 37192 6016
rect 37256 5952 37262 6016
rect 36946 5951 37262 5952
rect 2606 5472 2922 5473
rect 2606 5408 2612 5472
rect 2676 5408 2692 5472
rect 2756 5408 2772 5472
rect 2836 5408 2852 5472
rect 2916 5408 2922 5472
rect 2606 5407 2922 5408
rect 7606 5472 7922 5473
rect 7606 5408 7612 5472
rect 7676 5408 7692 5472
rect 7756 5408 7772 5472
rect 7836 5408 7852 5472
rect 7916 5408 7922 5472
rect 7606 5407 7922 5408
rect 12606 5472 12922 5473
rect 12606 5408 12612 5472
rect 12676 5408 12692 5472
rect 12756 5408 12772 5472
rect 12836 5408 12852 5472
rect 12916 5408 12922 5472
rect 12606 5407 12922 5408
rect 17606 5472 17922 5473
rect 17606 5408 17612 5472
rect 17676 5408 17692 5472
rect 17756 5408 17772 5472
rect 17836 5408 17852 5472
rect 17916 5408 17922 5472
rect 17606 5407 17922 5408
rect 22606 5472 22922 5473
rect 22606 5408 22612 5472
rect 22676 5408 22692 5472
rect 22756 5408 22772 5472
rect 22836 5408 22852 5472
rect 22916 5408 22922 5472
rect 22606 5407 22922 5408
rect 27606 5472 27922 5473
rect 27606 5408 27612 5472
rect 27676 5408 27692 5472
rect 27756 5408 27772 5472
rect 27836 5408 27852 5472
rect 27916 5408 27922 5472
rect 27606 5407 27922 5408
rect 32606 5472 32922 5473
rect 32606 5408 32612 5472
rect 32676 5408 32692 5472
rect 32756 5408 32772 5472
rect 32836 5408 32852 5472
rect 32916 5408 32922 5472
rect 32606 5407 32922 5408
rect 37606 5472 37922 5473
rect 37606 5408 37612 5472
rect 37676 5408 37692 5472
rect 37756 5408 37772 5472
rect 37836 5408 37852 5472
rect 37916 5408 37922 5472
rect 37606 5407 37922 5408
rect 1946 4928 2262 4929
rect 1946 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2262 4928
rect 1946 4863 2262 4864
rect 6946 4928 7262 4929
rect 6946 4864 6952 4928
rect 7016 4864 7032 4928
rect 7096 4864 7112 4928
rect 7176 4864 7192 4928
rect 7256 4864 7262 4928
rect 6946 4863 7262 4864
rect 11946 4928 12262 4929
rect 11946 4864 11952 4928
rect 12016 4864 12032 4928
rect 12096 4864 12112 4928
rect 12176 4864 12192 4928
rect 12256 4864 12262 4928
rect 11946 4863 12262 4864
rect 16946 4928 17262 4929
rect 16946 4864 16952 4928
rect 17016 4864 17032 4928
rect 17096 4864 17112 4928
rect 17176 4864 17192 4928
rect 17256 4864 17262 4928
rect 16946 4863 17262 4864
rect 21946 4928 22262 4929
rect 21946 4864 21952 4928
rect 22016 4864 22032 4928
rect 22096 4864 22112 4928
rect 22176 4864 22192 4928
rect 22256 4864 22262 4928
rect 21946 4863 22262 4864
rect 26946 4928 27262 4929
rect 26946 4864 26952 4928
rect 27016 4864 27032 4928
rect 27096 4864 27112 4928
rect 27176 4864 27192 4928
rect 27256 4864 27262 4928
rect 26946 4863 27262 4864
rect 31946 4928 32262 4929
rect 31946 4864 31952 4928
rect 32016 4864 32032 4928
rect 32096 4864 32112 4928
rect 32176 4864 32192 4928
rect 32256 4864 32262 4928
rect 31946 4863 32262 4864
rect 36946 4928 37262 4929
rect 36946 4864 36952 4928
rect 37016 4864 37032 4928
rect 37096 4864 37112 4928
rect 37176 4864 37192 4928
rect 37256 4864 37262 4928
rect 36946 4863 37262 4864
rect 841 4586 907 4589
rect 798 4584 907 4586
rect 798 4528 846 4584
rect 902 4528 907 4584
rect 798 4523 907 4528
rect 798 4480 858 4523
rect 0 4390 858 4480
rect 40493 4450 40559 4453
rect 41200 4450 42000 4480
rect 40493 4448 42000 4450
rect 40493 4392 40498 4448
rect 40554 4392 42000 4448
rect 40493 4390 42000 4392
rect 0 4360 800 4390
rect 40493 4387 40559 4390
rect 2606 4384 2922 4385
rect 2606 4320 2612 4384
rect 2676 4320 2692 4384
rect 2756 4320 2772 4384
rect 2836 4320 2852 4384
rect 2916 4320 2922 4384
rect 2606 4319 2922 4320
rect 7606 4384 7922 4385
rect 7606 4320 7612 4384
rect 7676 4320 7692 4384
rect 7756 4320 7772 4384
rect 7836 4320 7852 4384
rect 7916 4320 7922 4384
rect 7606 4319 7922 4320
rect 12606 4384 12922 4385
rect 12606 4320 12612 4384
rect 12676 4320 12692 4384
rect 12756 4320 12772 4384
rect 12836 4320 12852 4384
rect 12916 4320 12922 4384
rect 12606 4319 12922 4320
rect 17606 4384 17922 4385
rect 17606 4320 17612 4384
rect 17676 4320 17692 4384
rect 17756 4320 17772 4384
rect 17836 4320 17852 4384
rect 17916 4320 17922 4384
rect 17606 4319 17922 4320
rect 22606 4384 22922 4385
rect 22606 4320 22612 4384
rect 22676 4320 22692 4384
rect 22756 4320 22772 4384
rect 22836 4320 22852 4384
rect 22916 4320 22922 4384
rect 22606 4319 22922 4320
rect 27606 4384 27922 4385
rect 27606 4320 27612 4384
rect 27676 4320 27692 4384
rect 27756 4320 27772 4384
rect 27836 4320 27852 4384
rect 27916 4320 27922 4384
rect 27606 4319 27922 4320
rect 32606 4384 32922 4385
rect 32606 4320 32612 4384
rect 32676 4320 32692 4384
rect 32756 4320 32772 4384
rect 32836 4320 32852 4384
rect 32916 4320 32922 4384
rect 32606 4319 32922 4320
rect 37606 4384 37922 4385
rect 37606 4320 37612 4384
rect 37676 4320 37692 4384
rect 37756 4320 37772 4384
rect 37836 4320 37852 4384
rect 37916 4320 37922 4384
rect 41200 4360 42000 4390
rect 37606 4319 37922 4320
rect 1946 3840 2262 3841
rect 1946 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2262 3840
rect 1946 3775 2262 3776
rect 6946 3840 7262 3841
rect 6946 3776 6952 3840
rect 7016 3776 7032 3840
rect 7096 3776 7112 3840
rect 7176 3776 7192 3840
rect 7256 3776 7262 3840
rect 6946 3775 7262 3776
rect 11946 3840 12262 3841
rect 11946 3776 11952 3840
rect 12016 3776 12032 3840
rect 12096 3776 12112 3840
rect 12176 3776 12192 3840
rect 12256 3776 12262 3840
rect 11946 3775 12262 3776
rect 16946 3840 17262 3841
rect 16946 3776 16952 3840
rect 17016 3776 17032 3840
rect 17096 3776 17112 3840
rect 17176 3776 17192 3840
rect 17256 3776 17262 3840
rect 16946 3775 17262 3776
rect 21946 3840 22262 3841
rect 21946 3776 21952 3840
rect 22016 3776 22032 3840
rect 22096 3776 22112 3840
rect 22176 3776 22192 3840
rect 22256 3776 22262 3840
rect 21946 3775 22262 3776
rect 26946 3840 27262 3841
rect 26946 3776 26952 3840
rect 27016 3776 27032 3840
rect 27096 3776 27112 3840
rect 27176 3776 27192 3840
rect 27256 3776 27262 3840
rect 26946 3775 27262 3776
rect 31946 3840 32262 3841
rect 31946 3776 31952 3840
rect 32016 3776 32032 3840
rect 32096 3776 32112 3840
rect 32176 3776 32192 3840
rect 32256 3776 32262 3840
rect 31946 3775 32262 3776
rect 36946 3840 37262 3841
rect 36946 3776 36952 3840
rect 37016 3776 37032 3840
rect 37096 3776 37112 3840
rect 37176 3776 37192 3840
rect 37256 3776 37262 3840
rect 36946 3775 37262 3776
rect 2606 3296 2922 3297
rect 2606 3232 2612 3296
rect 2676 3232 2692 3296
rect 2756 3232 2772 3296
rect 2836 3232 2852 3296
rect 2916 3232 2922 3296
rect 2606 3231 2922 3232
rect 7606 3296 7922 3297
rect 7606 3232 7612 3296
rect 7676 3232 7692 3296
rect 7756 3232 7772 3296
rect 7836 3232 7852 3296
rect 7916 3232 7922 3296
rect 7606 3231 7922 3232
rect 12606 3296 12922 3297
rect 12606 3232 12612 3296
rect 12676 3232 12692 3296
rect 12756 3232 12772 3296
rect 12836 3232 12852 3296
rect 12916 3232 12922 3296
rect 12606 3231 12922 3232
rect 17606 3296 17922 3297
rect 17606 3232 17612 3296
rect 17676 3232 17692 3296
rect 17756 3232 17772 3296
rect 17836 3232 17852 3296
rect 17916 3232 17922 3296
rect 17606 3231 17922 3232
rect 22606 3296 22922 3297
rect 22606 3232 22612 3296
rect 22676 3232 22692 3296
rect 22756 3232 22772 3296
rect 22836 3232 22852 3296
rect 22916 3232 22922 3296
rect 22606 3231 22922 3232
rect 27606 3296 27922 3297
rect 27606 3232 27612 3296
rect 27676 3232 27692 3296
rect 27756 3232 27772 3296
rect 27836 3232 27852 3296
rect 27916 3232 27922 3296
rect 27606 3231 27922 3232
rect 32606 3296 32922 3297
rect 32606 3232 32612 3296
rect 32676 3232 32692 3296
rect 32756 3232 32772 3296
rect 32836 3232 32852 3296
rect 32916 3232 32922 3296
rect 32606 3231 32922 3232
rect 37606 3296 37922 3297
rect 37606 3232 37612 3296
rect 37676 3232 37692 3296
rect 37756 3232 37772 3296
rect 37836 3232 37852 3296
rect 37916 3232 37922 3296
rect 37606 3231 37922 3232
rect 1946 2752 2262 2753
rect 1946 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2262 2752
rect 1946 2687 2262 2688
rect 6946 2752 7262 2753
rect 6946 2688 6952 2752
rect 7016 2688 7032 2752
rect 7096 2688 7112 2752
rect 7176 2688 7192 2752
rect 7256 2688 7262 2752
rect 6946 2687 7262 2688
rect 11946 2752 12262 2753
rect 11946 2688 11952 2752
rect 12016 2688 12032 2752
rect 12096 2688 12112 2752
rect 12176 2688 12192 2752
rect 12256 2688 12262 2752
rect 11946 2687 12262 2688
rect 16946 2752 17262 2753
rect 16946 2688 16952 2752
rect 17016 2688 17032 2752
rect 17096 2688 17112 2752
rect 17176 2688 17192 2752
rect 17256 2688 17262 2752
rect 16946 2687 17262 2688
rect 21946 2752 22262 2753
rect 21946 2688 21952 2752
rect 22016 2688 22032 2752
rect 22096 2688 22112 2752
rect 22176 2688 22192 2752
rect 22256 2688 22262 2752
rect 21946 2687 22262 2688
rect 26946 2752 27262 2753
rect 26946 2688 26952 2752
rect 27016 2688 27032 2752
rect 27096 2688 27112 2752
rect 27176 2688 27192 2752
rect 27256 2688 27262 2752
rect 26946 2687 27262 2688
rect 31946 2752 32262 2753
rect 31946 2688 31952 2752
rect 32016 2688 32032 2752
rect 32096 2688 32112 2752
rect 32176 2688 32192 2752
rect 32256 2688 32262 2752
rect 31946 2687 32262 2688
rect 36946 2752 37262 2753
rect 36946 2688 36952 2752
rect 37016 2688 37032 2752
rect 37096 2688 37112 2752
rect 37176 2688 37192 2752
rect 37256 2688 37262 2752
rect 36946 2687 37262 2688
rect 16430 2348 16436 2412
rect 16500 2410 16506 2412
rect 28625 2410 28691 2413
rect 16500 2408 28691 2410
rect 16500 2352 28630 2408
rect 28686 2352 28691 2408
rect 16500 2350 28691 2352
rect 16500 2348 16506 2350
rect 28625 2347 28691 2350
rect 2606 2208 2922 2209
rect 2606 2144 2612 2208
rect 2676 2144 2692 2208
rect 2756 2144 2772 2208
rect 2836 2144 2852 2208
rect 2916 2144 2922 2208
rect 2606 2143 2922 2144
rect 7606 2208 7922 2209
rect 7606 2144 7612 2208
rect 7676 2144 7692 2208
rect 7756 2144 7772 2208
rect 7836 2144 7852 2208
rect 7916 2144 7922 2208
rect 7606 2143 7922 2144
rect 12606 2208 12922 2209
rect 12606 2144 12612 2208
rect 12676 2144 12692 2208
rect 12756 2144 12772 2208
rect 12836 2144 12852 2208
rect 12916 2144 12922 2208
rect 12606 2143 12922 2144
rect 17606 2208 17922 2209
rect 17606 2144 17612 2208
rect 17676 2144 17692 2208
rect 17756 2144 17772 2208
rect 17836 2144 17852 2208
rect 17916 2144 17922 2208
rect 17606 2143 17922 2144
rect 22606 2208 22922 2209
rect 22606 2144 22612 2208
rect 22676 2144 22692 2208
rect 22756 2144 22772 2208
rect 22836 2144 22852 2208
rect 22916 2144 22922 2208
rect 22606 2143 22922 2144
rect 27606 2208 27922 2209
rect 27606 2144 27612 2208
rect 27676 2144 27692 2208
rect 27756 2144 27772 2208
rect 27836 2144 27852 2208
rect 27916 2144 27922 2208
rect 27606 2143 27922 2144
rect 32606 2208 32922 2209
rect 32606 2144 32612 2208
rect 32676 2144 32692 2208
rect 32756 2144 32772 2208
rect 32836 2144 32852 2208
rect 32916 2144 32922 2208
rect 32606 2143 32922 2144
rect 37606 2208 37922 2209
rect 37606 2144 37612 2208
rect 37676 2144 37692 2208
rect 37756 2144 37772 2208
rect 37836 2144 37852 2208
rect 37916 2144 37922 2208
rect 37606 2143 37922 2144
<< via3 >>
rect 2612 69660 2676 69664
rect 2612 69604 2616 69660
rect 2616 69604 2672 69660
rect 2672 69604 2676 69660
rect 2612 69600 2676 69604
rect 2692 69660 2756 69664
rect 2692 69604 2696 69660
rect 2696 69604 2752 69660
rect 2752 69604 2756 69660
rect 2692 69600 2756 69604
rect 2772 69660 2836 69664
rect 2772 69604 2776 69660
rect 2776 69604 2832 69660
rect 2832 69604 2836 69660
rect 2772 69600 2836 69604
rect 2852 69660 2916 69664
rect 2852 69604 2856 69660
rect 2856 69604 2912 69660
rect 2912 69604 2916 69660
rect 2852 69600 2916 69604
rect 7612 69660 7676 69664
rect 7612 69604 7616 69660
rect 7616 69604 7672 69660
rect 7672 69604 7676 69660
rect 7612 69600 7676 69604
rect 7692 69660 7756 69664
rect 7692 69604 7696 69660
rect 7696 69604 7752 69660
rect 7752 69604 7756 69660
rect 7692 69600 7756 69604
rect 7772 69660 7836 69664
rect 7772 69604 7776 69660
rect 7776 69604 7832 69660
rect 7832 69604 7836 69660
rect 7772 69600 7836 69604
rect 7852 69660 7916 69664
rect 7852 69604 7856 69660
rect 7856 69604 7912 69660
rect 7912 69604 7916 69660
rect 7852 69600 7916 69604
rect 12612 69660 12676 69664
rect 12612 69604 12616 69660
rect 12616 69604 12672 69660
rect 12672 69604 12676 69660
rect 12612 69600 12676 69604
rect 12692 69660 12756 69664
rect 12692 69604 12696 69660
rect 12696 69604 12752 69660
rect 12752 69604 12756 69660
rect 12692 69600 12756 69604
rect 12772 69660 12836 69664
rect 12772 69604 12776 69660
rect 12776 69604 12832 69660
rect 12832 69604 12836 69660
rect 12772 69600 12836 69604
rect 12852 69660 12916 69664
rect 12852 69604 12856 69660
rect 12856 69604 12912 69660
rect 12912 69604 12916 69660
rect 12852 69600 12916 69604
rect 17612 69660 17676 69664
rect 17612 69604 17616 69660
rect 17616 69604 17672 69660
rect 17672 69604 17676 69660
rect 17612 69600 17676 69604
rect 17692 69660 17756 69664
rect 17692 69604 17696 69660
rect 17696 69604 17752 69660
rect 17752 69604 17756 69660
rect 17692 69600 17756 69604
rect 17772 69660 17836 69664
rect 17772 69604 17776 69660
rect 17776 69604 17832 69660
rect 17832 69604 17836 69660
rect 17772 69600 17836 69604
rect 17852 69660 17916 69664
rect 17852 69604 17856 69660
rect 17856 69604 17912 69660
rect 17912 69604 17916 69660
rect 17852 69600 17916 69604
rect 22612 69660 22676 69664
rect 22612 69604 22616 69660
rect 22616 69604 22672 69660
rect 22672 69604 22676 69660
rect 22612 69600 22676 69604
rect 22692 69660 22756 69664
rect 22692 69604 22696 69660
rect 22696 69604 22752 69660
rect 22752 69604 22756 69660
rect 22692 69600 22756 69604
rect 22772 69660 22836 69664
rect 22772 69604 22776 69660
rect 22776 69604 22832 69660
rect 22832 69604 22836 69660
rect 22772 69600 22836 69604
rect 22852 69660 22916 69664
rect 22852 69604 22856 69660
rect 22856 69604 22912 69660
rect 22912 69604 22916 69660
rect 22852 69600 22916 69604
rect 27612 69660 27676 69664
rect 27612 69604 27616 69660
rect 27616 69604 27672 69660
rect 27672 69604 27676 69660
rect 27612 69600 27676 69604
rect 27692 69660 27756 69664
rect 27692 69604 27696 69660
rect 27696 69604 27752 69660
rect 27752 69604 27756 69660
rect 27692 69600 27756 69604
rect 27772 69660 27836 69664
rect 27772 69604 27776 69660
rect 27776 69604 27832 69660
rect 27832 69604 27836 69660
rect 27772 69600 27836 69604
rect 27852 69660 27916 69664
rect 27852 69604 27856 69660
rect 27856 69604 27912 69660
rect 27912 69604 27916 69660
rect 27852 69600 27916 69604
rect 32612 69660 32676 69664
rect 32612 69604 32616 69660
rect 32616 69604 32672 69660
rect 32672 69604 32676 69660
rect 32612 69600 32676 69604
rect 32692 69660 32756 69664
rect 32692 69604 32696 69660
rect 32696 69604 32752 69660
rect 32752 69604 32756 69660
rect 32692 69600 32756 69604
rect 32772 69660 32836 69664
rect 32772 69604 32776 69660
rect 32776 69604 32832 69660
rect 32832 69604 32836 69660
rect 32772 69600 32836 69604
rect 32852 69660 32916 69664
rect 32852 69604 32856 69660
rect 32856 69604 32912 69660
rect 32912 69604 32916 69660
rect 32852 69600 32916 69604
rect 37612 69660 37676 69664
rect 37612 69604 37616 69660
rect 37616 69604 37672 69660
rect 37672 69604 37676 69660
rect 37612 69600 37676 69604
rect 37692 69660 37756 69664
rect 37692 69604 37696 69660
rect 37696 69604 37752 69660
rect 37752 69604 37756 69660
rect 37692 69600 37756 69604
rect 37772 69660 37836 69664
rect 37772 69604 37776 69660
rect 37776 69604 37832 69660
rect 37832 69604 37836 69660
rect 37772 69600 37836 69604
rect 37852 69660 37916 69664
rect 37852 69604 37856 69660
rect 37856 69604 37912 69660
rect 37912 69604 37916 69660
rect 37852 69600 37916 69604
rect 1952 69116 2016 69120
rect 1952 69060 1956 69116
rect 1956 69060 2012 69116
rect 2012 69060 2016 69116
rect 1952 69056 2016 69060
rect 2032 69116 2096 69120
rect 2032 69060 2036 69116
rect 2036 69060 2092 69116
rect 2092 69060 2096 69116
rect 2032 69056 2096 69060
rect 2112 69116 2176 69120
rect 2112 69060 2116 69116
rect 2116 69060 2172 69116
rect 2172 69060 2176 69116
rect 2112 69056 2176 69060
rect 2192 69116 2256 69120
rect 2192 69060 2196 69116
rect 2196 69060 2252 69116
rect 2252 69060 2256 69116
rect 2192 69056 2256 69060
rect 6952 69116 7016 69120
rect 6952 69060 6956 69116
rect 6956 69060 7012 69116
rect 7012 69060 7016 69116
rect 6952 69056 7016 69060
rect 7032 69116 7096 69120
rect 7032 69060 7036 69116
rect 7036 69060 7092 69116
rect 7092 69060 7096 69116
rect 7032 69056 7096 69060
rect 7112 69116 7176 69120
rect 7112 69060 7116 69116
rect 7116 69060 7172 69116
rect 7172 69060 7176 69116
rect 7112 69056 7176 69060
rect 7192 69116 7256 69120
rect 7192 69060 7196 69116
rect 7196 69060 7252 69116
rect 7252 69060 7256 69116
rect 7192 69056 7256 69060
rect 11952 69116 12016 69120
rect 11952 69060 11956 69116
rect 11956 69060 12012 69116
rect 12012 69060 12016 69116
rect 11952 69056 12016 69060
rect 12032 69116 12096 69120
rect 12032 69060 12036 69116
rect 12036 69060 12092 69116
rect 12092 69060 12096 69116
rect 12032 69056 12096 69060
rect 12112 69116 12176 69120
rect 12112 69060 12116 69116
rect 12116 69060 12172 69116
rect 12172 69060 12176 69116
rect 12112 69056 12176 69060
rect 12192 69116 12256 69120
rect 12192 69060 12196 69116
rect 12196 69060 12252 69116
rect 12252 69060 12256 69116
rect 12192 69056 12256 69060
rect 16952 69116 17016 69120
rect 16952 69060 16956 69116
rect 16956 69060 17012 69116
rect 17012 69060 17016 69116
rect 16952 69056 17016 69060
rect 17032 69116 17096 69120
rect 17032 69060 17036 69116
rect 17036 69060 17092 69116
rect 17092 69060 17096 69116
rect 17032 69056 17096 69060
rect 17112 69116 17176 69120
rect 17112 69060 17116 69116
rect 17116 69060 17172 69116
rect 17172 69060 17176 69116
rect 17112 69056 17176 69060
rect 17192 69116 17256 69120
rect 17192 69060 17196 69116
rect 17196 69060 17252 69116
rect 17252 69060 17256 69116
rect 17192 69056 17256 69060
rect 21952 69116 22016 69120
rect 21952 69060 21956 69116
rect 21956 69060 22012 69116
rect 22012 69060 22016 69116
rect 21952 69056 22016 69060
rect 22032 69116 22096 69120
rect 22032 69060 22036 69116
rect 22036 69060 22092 69116
rect 22092 69060 22096 69116
rect 22032 69056 22096 69060
rect 22112 69116 22176 69120
rect 22112 69060 22116 69116
rect 22116 69060 22172 69116
rect 22172 69060 22176 69116
rect 22112 69056 22176 69060
rect 22192 69116 22256 69120
rect 22192 69060 22196 69116
rect 22196 69060 22252 69116
rect 22252 69060 22256 69116
rect 22192 69056 22256 69060
rect 26952 69116 27016 69120
rect 26952 69060 26956 69116
rect 26956 69060 27012 69116
rect 27012 69060 27016 69116
rect 26952 69056 27016 69060
rect 27032 69116 27096 69120
rect 27032 69060 27036 69116
rect 27036 69060 27092 69116
rect 27092 69060 27096 69116
rect 27032 69056 27096 69060
rect 27112 69116 27176 69120
rect 27112 69060 27116 69116
rect 27116 69060 27172 69116
rect 27172 69060 27176 69116
rect 27112 69056 27176 69060
rect 27192 69116 27256 69120
rect 27192 69060 27196 69116
rect 27196 69060 27252 69116
rect 27252 69060 27256 69116
rect 27192 69056 27256 69060
rect 31952 69116 32016 69120
rect 31952 69060 31956 69116
rect 31956 69060 32012 69116
rect 32012 69060 32016 69116
rect 31952 69056 32016 69060
rect 32032 69116 32096 69120
rect 32032 69060 32036 69116
rect 32036 69060 32092 69116
rect 32092 69060 32096 69116
rect 32032 69056 32096 69060
rect 32112 69116 32176 69120
rect 32112 69060 32116 69116
rect 32116 69060 32172 69116
rect 32172 69060 32176 69116
rect 32112 69056 32176 69060
rect 32192 69116 32256 69120
rect 32192 69060 32196 69116
rect 32196 69060 32252 69116
rect 32252 69060 32256 69116
rect 32192 69056 32256 69060
rect 36952 69116 37016 69120
rect 36952 69060 36956 69116
rect 36956 69060 37012 69116
rect 37012 69060 37016 69116
rect 36952 69056 37016 69060
rect 37032 69116 37096 69120
rect 37032 69060 37036 69116
rect 37036 69060 37092 69116
rect 37092 69060 37096 69116
rect 37032 69056 37096 69060
rect 37112 69116 37176 69120
rect 37112 69060 37116 69116
rect 37116 69060 37172 69116
rect 37172 69060 37176 69116
rect 37112 69056 37176 69060
rect 37192 69116 37256 69120
rect 37192 69060 37196 69116
rect 37196 69060 37252 69116
rect 37252 69060 37256 69116
rect 37192 69056 37256 69060
rect 2612 68572 2676 68576
rect 2612 68516 2616 68572
rect 2616 68516 2672 68572
rect 2672 68516 2676 68572
rect 2612 68512 2676 68516
rect 2692 68572 2756 68576
rect 2692 68516 2696 68572
rect 2696 68516 2752 68572
rect 2752 68516 2756 68572
rect 2692 68512 2756 68516
rect 2772 68572 2836 68576
rect 2772 68516 2776 68572
rect 2776 68516 2832 68572
rect 2832 68516 2836 68572
rect 2772 68512 2836 68516
rect 2852 68572 2916 68576
rect 2852 68516 2856 68572
rect 2856 68516 2912 68572
rect 2912 68516 2916 68572
rect 2852 68512 2916 68516
rect 7612 68572 7676 68576
rect 7612 68516 7616 68572
rect 7616 68516 7672 68572
rect 7672 68516 7676 68572
rect 7612 68512 7676 68516
rect 7692 68572 7756 68576
rect 7692 68516 7696 68572
rect 7696 68516 7752 68572
rect 7752 68516 7756 68572
rect 7692 68512 7756 68516
rect 7772 68572 7836 68576
rect 7772 68516 7776 68572
rect 7776 68516 7832 68572
rect 7832 68516 7836 68572
rect 7772 68512 7836 68516
rect 7852 68572 7916 68576
rect 7852 68516 7856 68572
rect 7856 68516 7912 68572
rect 7912 68516 7916 68572
rect 7852 68512 7916 68516
rect 12612 68572 12676 68576
rect 12612 68516 12616 68572
rect 12616 68516 12672 68572
rect 12672 68516 12676 68572
rect 12612 68512 12676 68516
rect 12692 68572 12756 68576
rect 12692 68516 12696 68572
rect 12696 68516 12752 68572
rect 12752 68516 12756 68572
rect 12692 68512 12756 68516
rect 12772 68572 12836 68576
rect 12772 68516 12776 68572
rect 12776 68516 12832 68572
rect 12832 68516 12836 68572
rect 12772 68512 12836 68516
rect 12852 68572 12916 68576
rect 12852 68516 12856 68572
rect 12856 68516 12912 68572
rect 12912 68516 12916 68572
rect 12852 68512 12916 68516
rect 17612 68572 17676 68576
rect 17612 68516 17616 68572
rect 17616 68516 17672 68572
rect 17672 68516 17676 68572
rect 17612 68512 17676 68516
rect 17692 68572 17756 68576
rect 17692 68516 17696 68572
rect 17696 68516 17752 68572
rect 17752 68516 17756 68572
rect 17692 68512 17756 68516
rect 17772 68572 17836 68576
rect 17772 68516 17776 68572
rect 17776 68516 17832 68572
rect 17832 68516 17836 68572
rect 17772 68512 17836 68516
rect 17852 68572 17916 68576
rect 17852 68516 17856 68572
rect 17856 68516 17912 68572
rect 17912 68516 17916 68572
rect 17852 68512 17916 68516
rect 22612 68572 22676 68576
rect 22612 68516 22616 68572
rect 22616 68516 22672 68572
rect 22672 68516 22676 68572
rect 22612 68512 22676 68516
rect 22692 68572 22756 68576
rect 22692 68516 22696 68572
rect 22696 68516 22752 68572
rect 22752 68516 22756 68572
rect 22692 68512 22756 68516
rect 22772 68572 22836 68576
rect 22772 68516 22776 68572
rect 22776 68516 22832 68572
rect 22832 68516 22836 68572
rect 22772 68512 22836 68516
rect 22852 68572 22916 68576
rect 22852 68516 22856 68572
rect 22856 68516 22912 68572
rect 22912 68516 22916 68572
rect 22852 68512 22916 68516
rect 27612 68572 27676 68576
rect 27612 68516 27616 68572
rect 27616 68516 27672 68572
rect 27672 68516 27676 68572
rect 27612 68512 27676 68516
rect 27692 68572 27756 68576
rect 27692 68516 27696 68572
rect 27696 68516 27752 68572
rect 27752 68516 27756 68572
rect 27692 68512 27756 68516
rect 27772 68572 27836 68576
rect 27772 68516 27776 68572
rect 27776 68516 27832 68572
rect 27832 68516 27836 68572
rect 27772 68512 27836 68516
rect 27852 68572 27916 68576
rect 27852 68516 27856 68572
rect 27856 68516 27912 68572
rect 27912 68516 27916 68572
rect 27852 68512 27916 68516
rect 32612 68572 32676 68576
rect 32612 68516 32616 68572
rect 32616 68516 32672 68572
rect 32672 68516 32676 68572
rect 32612 68512 32676 68516
rect 32692 68572 32756 68576
rect 32692 68516 32696 68572
rect 32696 68516 32752 68572
rect 32752 68516 32756 68572
rect 32692 68512 32756 68516
rect 32772 68572 32836 68576
rect 32772 68516 32776 68572
rect 32776 68516 32832 68572
rect 32832 68516 32836 68572
rect 32772 68512 32836 68516
rect 32852 68572 32916 68576
rect 32852 68516 32856 68572
rect 32856 68516 32912 68572
rect 32912 68516 32916 68572
rect 32852 68512 32916 68516
rect 37612 68572 37676 68576
rect 37612 68516 37616 68572
rect 37616 68516 37672 68572
rect 37672 68516 37676 68572
rect 37612 68512 37676 68516
rect 37692 68572 37756 68576
rect 37692 68516 37696 68572
rect 37696 68516 37752 68572
rect 37752 68516 37756 68572
rect 37692 68512 37756 68516
rect 37772 68572 37836 68576
rect 37772 68516 37776 68572
rect 37776 68516 37832 68572
rect 37832 68516 37836 68572
rect 37772 68512 37836 68516
rect 37852 68572 37916 68576
rect 37852 68516 37856 68572
rect 37856 68516 37912 68572
rect 37912 68516 37916 68572
rect 37852 68512 37916 68516
rect 1952 68028 2016 68032
rect 1952 67972 1956 68028
rect 1956 67972 2012 68028
rect 2012 67972 2016 68028
rect 1952 67968 2016 67972
rect 2032 68028 2096 68032
rect 2032 67972 2036 68028
rect 2036 67972 2092 68028
rect 2092 67972 2096 68028
rect 2032 67968 2096 67972
rect 2112 68028 2176 68032
rect 2112 67972 2116 68028
rect 2116 67972 2172 68028
rect 2172 67972 2176 68028
rect 2112 67968 2176 67972
rect 2192 68028 2256 68032
rect 2192 67972 2196 68028
rect 2196 67972 2252 68028
rect 2252 67972 2256 68028
rect 2192 67968 2256 67972
rect 6952 68028 7016 68032
rect 6952 67972 6956 68028
rect 6956 67972 7012 68028
rect 7012 67972 7016 68028
rect 6952 67968 7016 67972
rect 7032 68028 7096 68032
rect 7032 67972 7036 68028
rect 7036 67972 7092 68028
rect 7092 67972 7096 68028
rect 7032 67968 7096 67972
rect 7112 68028 7176 68032
rect 7112 67972 7116 68028
rect 7116 67972 7172 68028
rect 7172 67972 7176 68028
rect 7112 67968 7176 67972
rect 7192 68028 7256 68032
rect 7192 67972 7196 68028
rect 7196 67972 7252 68028
rect 7252 67972 7256 68028
rect 7192 67968 7256 67972
rect 11952 68028 12016 68032
rect 11952 67972 11956 68028
rect 11956 67972 12012 68028
rect 12012 67972 12016 68028
rect 11952 67968 12016 67972
rect 12032 68028 12096 68032
rect 12032 67972 12036 68028
rect 12036 67972 12092 68028
rect 12092 67972 12096 68028
rect 12032 67968 12096 67972
rect 12112 68028 12176 68032
rect 12112 67972 12116 68028
rect 12116 67972 12172 68028
rect 12172 67972 12176 68028
rect 12112 67968 12176 67972
rect 12192 68028 12256 68032
rect 12192 67972 12196 68028
rect 12196 67972 12252 68028
rect 12252 67972 12256 68028
rect 12192 67968 12256 67972
rect 16952 68028 17016 68032
rect 16952 67972 16956 68028
rect 16956 67972 17012 68028
rect 17012 67972 17016 68028
rect 16952 67968 17016 67972
rect 17032 68028 17096 68032
rect 17032 67972 17036 68028
rect 17036 67972 17092 68028
rect 17092 67972 17096 68028
rect 17032 67968 17096 67972
rect 17112 68028 17176 68032
rect 17112 67972 17116 68028
rect 17116 67972 17172 68028
rect 17172 67972 17176 68028
rect 17112 67968 17176 67972
rect 17192 68028 17256 68032
rect 17192 67972 17196 68028
rect 17196 67972 17252 68028
rect 17252 67972 17256 68028
rect 17192 67968 17256 67972
rect 21952 68028 22016 68032
rect 21952 67972 21956 68028
rect 21956 67972 22012 68028
rect 22012 67972 22016 68028
rect 21952 67968 22016 67972
rect 22032 68028 22096 68032
rect 22032 67972 22036 68028
rect 22036 67972 22092 68028
rect 22092 67972 22096 68028
rect 22032 67968 22096 67972
rect 22112 68028 22176 68032
rect 22112 67972 22116 68028
rect 22116 67972 22172 68028
rect 22172 67972 22176 68028
rect 22112 67968 22176 67972
rect 22192 68028 22256 68032
rect 22192 67972 22196 68028
rect 22196 67972 22252 68028
rect 22252 67972 22256 68028
rect 22192 67968 22256 67972
rect 26952 68028 27016 68032
rect 26952 67972 26956 68028
rect 26956 67972 27012 68028
rect 27012 67972 27016 68028
rect 26952 67968 27016 67972
rect 27032 68028 27096 68032
rect 27032 67972 27036 68028
rect 27036 67972 27092 68028
rect 27092 67972 27096 68028
rect 27032 67968 27096 67972
rect 27112 68028 27176 68032
rect 27112 67972 27116 68028
rect 27116 67972 27172 68028
rect 27172 67972 27176 68028
rect 27112 67968 27176 67972
rect 27192 68028 27256 68032
rect 27192 67972 27196 68028
rect 27196 67972 27252 68028
rect 27252 67972 27256 68028
rect 27192 67968 27256 67972
rect 31952 68028 32016 68032
rect 31952 67972 31956 68028
rect 31956 67972 32012 68028
rect 32012 67972 32016 68028
rect 31952 67968 32016 67972
rect 32032 68028 32096 68032
rect 32032 67972 32036 68028
rect 32036 67972 32092 68028
rect 32092 67972 32096 68028
rect 32032 67968 32096 67972
rect 32112 68028 32176 68032
rect 32112 67972 32116 68028
rect 32116 67972 32172 68028
rect 32172 67972 32176 68028
rect 32112 67968 32176 67972
rect 32192 68028 32256 68032
rect 32192 67972 32196 68028
rect 32196 67972 32252 68028
rect 32252 67972 32256 68028
rect 32192 67968 32256 67972
rect 36952 68028 37016 68032
rect 36952 67972 36956 68028
rect 36956 67972 37012 68028
rect 37012 67972 37016 68028
rect 36952 67968 37016 67972
rect 37032 68028 37096 68032
rect 37032 67972 37036 68028
rect 37036 67972 37092 68028
rect 37092 67972 37096 68028
rect 37032 67968 37096 67972
rect 37112 68028 37176 68032
rect 37112 67972 37116 68028
rect 37116 67972 37172 68028
rect 37172 67972 37176 68028
rect 37112 67968 37176 67972
rect 37192 68028 37256 68032
rect 37192 67972 37196 68028
rect 37196 67972 37252 68028
rect 37252 67972 37256 68028
rect 37192 67968 37256 67972
rect 14964 67764 15028 67828
rect 3372 67628 3436 67692
rect 2612 67484 2676 67488
rect 2612 67428 2616 67484
rect 2616 67428 2672 67484
rect 2672 67428 2676 67484
rect 2612 67424 2676 67428
rect 2692 67484 2756 67488
rect 2692 67428 2696 67484
rect 2696 67428 2752 67484
rect 2752 67428 2756 67484
rect 2692 67424 2756 67428
rect 2772 67484 2836 67488
rect 2772 67428 2776 67484
rect 2776 67428 2832 67484
rect 2832 67428 2836 67484
rect 2772 67424 2836 67428
rect 2852 67484 2916 67488
rect 2852 67428 2856 67484
rect 2856 67428 2912 67484
rect 2912 67428 2916 67484
rect 2852 67424 2916 67428
rect 7612 67484 7676 67488
rect 7612 67428 7616 67484
rect 7616 67428 7672 67484
rect 7672 67428 7676 67484
rect 7612 67424 7676 67428
rect 7692 67484 7756 67488
rect 7692 67428 7696 67484
rect 7696 67428 7752 67484
rect 7752 67428 7756 67484
rect 7692 67424 7756 67428
rect 7772 67484 7836 67488
rect 7772 67428 7776 67484
rect 7776 67428 7832 67484
rect 7832 67428 7836 67484
rect 7772 67424 7836 67428
rect 7852 67484 7916 67488
rect 7852 67428 7856 67484
rect 7856 67428 7912 67484
rect 7912 67428 7916 67484
rect 7852 67424 7916 67428
rect 12612 67484 12676 67488
rect 12612 67428 12616 67484
rect 12616 67428 12672 67484
rect 12672 67428 12676 67484
rect 12612 67424 12676 67428
rect 12692 67484 12756 67488
rect 12692 67428 12696 67484
rect 12696 67428 12752 67484
rect 12752 67428 12756 67484
rect 12692 67424 12756 67428
rect 12772 67484 12836 67488
rect 12772 67428 12776 67484
rect 12776 67428 12832 67484
rect 12832 67428 12836 67484
rect 12772 67424 12836 67428
rect 12852 67484 12916 67488
rect 12852 67428 12856 67484
rect 12856 67428 12912 67484
rect 12912 67428 12916 67484
rect 12852 67424 12916 67428
rect 17612 67484 17676 67488
rect 17612 67428 17616 67484
rect 17616 67428 17672 67484
rect 17672 67428 17676 67484
rect 17612 67424 17676 67428
rect 17692 67484 17756 67488
rect 17692 67428 17696 67484
rect 17696 67428 17752 67484
rect 17752 67428 17756 67484
rect 17692 67424 17756 67428
rect 17772 67484 17836 67488
rect 17772 67428 17776 67484
rect 17776 67428 17832 67484
rect 17832 67428 17836 67484
rect 17772 67424 17836 67428
rect 17852 67484 17916 67488
rect 17852 67428 17856 67484
rect 17856 67428 17912 67484
rect 17912 67428 17916 67484
rect 17852 67424 17916 67428
rect 22612 67484 22676 67488
rect 22612 67428 22616 67484
rect 22616 67428 22672 67484
rect 22672 67428 22676 67484
rect 22612 67424 22676 67428
rect 22692 67484 22756 67488
rect 22692 67428 22696 67484
rect 22696 67428 22752 67484
rect 22752 67428 22756 67484
rect 22692 67424 22756 67428
rect 22772 67484 22836 67488
rect 22772 67428 22776 67484
rect 22776 67428 22832 67484
rect 22832 67428 22836 67484
rect 22772 67424 22836 67428
rect 22852 67484 22916 67488
rect 22852 67428 22856 67484
rect 22856 67428 22912 67484
rect 22912 67428 22916 67484
rect 22852 67424 22916 67428
rect 27612 67484 27676 67488
rect 27612 67428 27616 67484
rect 27616 67428 27672 67484
rect 27672 67428 27676 67484
rect 27612 67424 27676 67428
rect 27692 67484 27756 67488
rect 27692 67428 27696 67484
rect 27696 67428 27752 67484
rect 27752 67428 27756 67484
rect 27692 67424 27756 67428
rect 27772 67484 27836 67488
rect 27772 67428 27776 67484
rect 27776 67428 27832 67484
rect 27832 67428 27836 67484
rect 27772 67424 27836 67428
rect 27852 67484 27916 67488
rect 27852 67428 27856 67484
rect 27856 67428 27912 67484
rect 27912 67428 27916 67484
rect 27852 67424 27916 67428
rect 32612 67484 32676 67488
rect 32612 67428 32616 67484
rect 32616 67428 32672 67484
rect 32672 67428 32676 67484
rect 32612 67424 32676 67428
rect 32692 67484 32756 67488
rect 32692 67428 32696 67484
rect 32696 67428 32752 67484
rect 32752 67428 32756 67484
rect 32692 67424 32756 67428
rect 32772 67484 32836 67488
rect 32772 67428 32776 67484
rect 32776 67428 32832 67484
rect 32832 67428 32836 67484
rect 32772 67424 32836 67428
rect 32852 67484 32916 67488
rect 32852 67428 32856 67484
rect 32856 67428 32912 67484
rect 32912 67428 32916 67484
rect 32852 67424 32916 67428
rect 37612 67484 37676 67488
rect 37612 67428 37616 67484
rect 37616 67428 37672 67484
rect 37672 67428 37676 67484
rect 37612 67424 37676 67428
rect 37692 67484 37756 67488
rect 37692 67428 37696 67484
rect 37696 67428 37752 67484
rect 37752 67428 37756 67484
rect 37692 67424 37756 67428
rect 37772 67484 37836 67488
rect 37772 67428 37776 67484
rect 37776 67428 37832 67484
rect 37832 67428 37836 67484
rect 37772 67424 37836 67428
rect 37852 67484 37916 67488
rect 37852 67428 37856 67484
rect 37856 67428 37912 67484
rect 37912 67428 37916 67484
rect 37852 67424 37916 67428
rect 1952 66940 2016 66944
rect 1952 66884 1956 66940
rect 1956 66884 2012 66940
rect 2012 66884 2016 66940
rect 1952 66880 2016 66884
rect 2032 66940 2096 66944
rect 2032 66884 2036 66940
rect 2036 66884 2092 66940
rect 2092 66884 2096 66940
rect 2032 66880 2096 66884
rect 2112 66940 2176 66944
rect 2112 66884 2116 66940
rect 2116 66884 2172 66940
rect 2172 66884 2176 66940
rect 2112 66880 2176 66884
rect 2192 66940 2256 66944
rect 2192 66884 2196 66940
rect 2196 66884 2252 66940
rect 2252 66884 2256 66940
rect 2192 66880 2256 66884
rect 6952 66940 7016 66944
rect 6952 66884 6956 66940
rect 6956 66884 7012 66940
rect 7012 66884 7016 66940
rect 6952 66880 7016 66884
rect 7032 66940 7096 66944
rect 7032 66884 7036 66940
rect 7036 66884 7092 66940
rect 7092 66884 7096 66940
rect 7032 66880 7096 66884
rect 7112 66940 7176 66944
rect 7112 66884 7116 66940
rect 7116 66884 7172 66940
rect 7172 66884 7176 66940
rect 7112 66880 7176 66884
rect 7192 66940 7256 66944
rect 7192 66884 7196 66940
rect 7196 66884 7252 66940
rect 7252 66884 7256 66940
rect 7192 66880 7256 66884
rect 11952 66940 12016 66944
rect 11952 66884 11956 66940
rect 11956 66884 12012 66940
rect 12012 66884 12016 66940
rect 11952 66880 12016 66884
rect 12032 66940 12096 66944
rect 12032 66884 12036 66940
rect 12036 66884 12092 66940
rect 12092 66884 12096 66940
rect 12032 66880 12096 66884
rect 12112 66940 12176 66944
rect 12112 66884 12116 66940
rect 12116 66884 12172 66940
rect 12172 66884 12176 66940
rect 12112 66880 12176 66884
rect 12192 66940 12256 66944
rect 12192 66884 12196 66940
rect 12196 66884 12252 66940
rect 12252 66884 12256 66940
rect 12192 66880 12256 66884
rect 16952 66940 17016 66944
rect 16952 66884 16956 66940
rect 16956 66884 17012 66940
rect 17012 66884 17016 66940
rect 16952 66880 17016 66884
rect 17032 66940 17096 66944
rect 17032 66884 17036 66940
rect 17036 66884 17092 66940
rect 17092 66884 17096 66940
rect 17032 66880 17096 66884
rect 17112 66940 17176 66944
rect 17112 66884 17116 66940
rect 17116 66884 17172 66940
rect 17172 66884 17176 66940
rect 17112 66880 17176 66884
rect 17192 66940 17256 66944
rect 17192 66884 17196 66940
rect 17196 66884 17252 66940
rect 17252 66884 17256 66940
rect 17192 66880 17256 66884
rect 21952 66940 22016 66944
rect 21952 66884 21956 66940
rect 21956 66884 22012 66940
rect 22012 66884 22016 66940
rect 21952 66880 22016 66884
rect 22032 66940 22096 66944
rect 22032 66884 22036 66940
rect 22036 66884 22092 66940
rect 22092 66884 22096 66940
rect 22032 66880 22096 66884
rect 22112 66940 22176 66944
rect 22112 66884 22116 66940
rect 22116 66884 22172 66940
rect 22172 66884 22176 66940
rect 22112 66880 22176 66884
rect 22192 66940 22256 66944
rect 22192 66884 22196 66940
rect 22196 66884 22252 66940
rect 22252 66884 22256 66940
rect 22192 66880 22256 66884
rect 26952 66940 27016 66944
rect 26952 66884 26956 66940
rect 26956 66884 27012 66940
rect 27012 66884 27016 66940
rect 26952 66880 27016 66884
rect 27032 66940 27096 66944
rect 27032 66884 27036 66940
rect 27036 66884 27092 66940
rect 27092 66884 27096 66940
rect 27032 66880 27096 66884
rect 27112 66940 27176 66944
rect 27112 66884 27116 66940
rect 27116 66884 27172 66940
rect 27172 66884 27176 66940
rect 27112 66880 27176 66884
rect 27192 66940 27256 66944
rect 27192 66884 27196 66940
rect 27196 66884 27252 66940
rect 27252 66884 27256 66940
rect 27192 66880 27256 66884
rect 31952 66940 32016 66944
rect 31952 66884 31956 66940
rect 31956 66884 32012 66940
rect 32012 66884 32016 66940
rect 31952 66880 32016 66884
rect 32032 66940 32096 66944
rect 32032 66884 32036 66940
rect 32036 66884 32092 66940
rect 32092 66884 32096 66940
rect 32032 66880 32096 66884
rect 32112 66940 32176 66944
rect 32112 66884 32116 66940
rect 32116 66884 32172 66940
rect 32172 66884 32176 66940
rect 32112 66880 32176 66884
rect 32192 66940 32256 66944
rect 32192 66884 32196 66940
rect 32196 66884 32252 66940
rect 32252 66884 32256 66940
rect 32192 66880 32256 66884
rect 36952 66940 37016 66944
rect 36952 66884 36956 66940
rect 36956 66884 37012 66940
rect 37012 66884 37016 66940
rect 36952 66880 37016 66884
rect 37032 66940 37096 66944
rect 37032 66884 37036 66940
rect 37036 66884 37092 66940
rect 37092 66884 37096 66940
rect 37032 66880 37096 66884
rect 37112 66940 37176 66944
rect 37112 66884 37116 66940
rect 37116 66884 37172 66940
rect 37172 66884 37176 66940
rect 37112 66880 37176 66884
rect 37192 66940 37256 66944
rect 37192 66884 37196 66940
rect 37196 66884 37252 66940
rect 37252 66884 37256 66940
rect 37192 66880 37256 66884
rect 2612 66396 2676 66400
rect 2612 66340 2616 66396
rect 2616 66340 2672 66396
rect 2672 66340 2676 66396
rect 2612 66336 2676 66340
rect 2692 66396 2756 66400
rect 2692 66340 2696 66396
rect 2696 66340 2752 66396
rect 2752 66340 2756 66396
rect 2692 66336 2756 66340
rect 2772 66396 2836 66400
rect 2772 66340 2776 66396
rect 2776 66340 2832 66396
rect 2832 66340 2836 66396
rect 2772 66336 2836 66340
rect 2852 66396 2916 66400
rect 2852 66340 2856 66396
rect 2856 66340 2912 66396
rect 2912 66340 2916 66396
rect 2852 66336 2916 66340
rect 7612 66396 7676 66400
rect 7612 66340 7616 66396
rect 7616 66340 7672 66396
rect 7672 66340 7676 66396
rect 7612 66336 7676 66340
rect 7692 66396 7756 66400
rect 7692 66340 7696 66396
rect 7696 66340 7752 66396
rect 7752 66340 7756 66396
rect 7692 66336 7756 66340
rect 7772 66396 7836 66400
rect 7772 66340 7776 66396
rect 7776 66340 7832 66396
rect 7832 66340 7836 66396
rect 7772 66336 7836 66340
rect 7852 66396 7916 66400
rect 7852 66340 7856 66396
rect 7856 66340 7912 66396
rect 7912 66340 7916 66396
rect 7852 66336 7916 66340
rect 12612 66396 12676 66400
rect 12612 66340 12616 66396
rect 12616 66340 12672 66396
rect 12672 66340 12676 66396
rect 12612 66336 12676 66340
rect 12692 66396 12756 66400
rect 12692 66340 12696 66396
rect 12696 66340 12752 66396
rect 12752 66340 12756 66396
rect 12692 66336 12756 66340
rect 12772 66396 12836 66400
rect 12772 66340 12776 66396
rect 12776 66340 12832 66396
rect 12832 66340 12836 66396
rect 12772 66336 12836 66340
rect 12852 66396 12916 66400
rect 12852 66340 12856 66396
rect 12856 66340 12912 66396
rect 12912 66340 12916 66396
rect 12852 66336 12916 66340
rect 17612 66396 17676 66400
rect 17612 66340 17616 66396
rect 17616 66340 17672 66396
rect 17672 66340 17676 66396
rect 17612 66336 17676 66340
rect 17692 66396 17756 66400
rect 17692 66340 17696 66396
rect 17696 66340 17752 66396
rect 17752 66340 17756 66396
rect 17692 66336 17756 66340
rect 17772 66396 17836 66400
rect 17772 66340 17776 66396
rect 17776 66340 17832 66396
rect 17832 66340 17836 66396
rect 17772 66336 17836 66340
rect 17852 66396 17916 66400
rect 17852 66340 17856 66396
rect 17856 66340 17912 66396
rect 17912 66340 17916 66396
rect 17852 66336 17916 66340
rect 22612 66396 22676 66400
rect 22612 66340 22616 66396
rect 22616 66340 22672 66396
rect 22672 66340 22676 66396
rect 22612 66336 22676 66340
rect 22692 66396 22756 66400
rect 22692 66340 22696 66396
rect 22696 66340 22752 66396
rect 22752 66340 22756 66396
rect 22692 66336 22756 66340
rect 22772 66396 22836 66400
rect 22772 66340 22776 66396
rect 22776 66340 22832 66396
rect 22832 66340 22836 66396
rect 22772 66336 22836 66340
rect 22852 66396 22916 66400
rect 22852 66340 22856 66396
rect 22856 66340 22912 66396
rect 22912 66340 22916 66396
rect 22852 66336 22916 66340
rect 27612 66396 27676 66400
rect 27612 66340 27616 66396
rect 27616 66340 27672 66396
rect 27672 66340 27676 66396
rect 27612 66336 27676 66340
rect 27692 66396 27756 66400
rect 27692 66340 27696 66396
rect 27696 66340 27752 66396
rect 27752 66340 27756 66396
rect 27692 66336 27756 66340
rect 27772 66396 27836 66400
rect 27772 66340 27776 66396
rect 27776 66340 27832 66396
rect 27832 66340 27836 66396
rect 27772 66336 27836 66340
rect 27852 66396 27916 66400
rect 27852 66340 27856 66396
rect 27856 66340 27912 66396
rect 27912 66340 27916 66396
rect 27852 66336 27916 66340
rect 32612 66396 32676 66400
rect 32612 66340 32616 66396
rect 32616 66340 32672 66396
rect 32672 66340 32676 66396
rect 32612 66336 32676 66340
rect 32692 66396 32756 66400
rect 32692 66340 32696 66396
rect 32696 66340 32752 66396
rect 32752 66340 32756 66396
rect 32692 66336 32756 66340
rect 32772 66396 32836 66400
rect 32772 66340 32776 66396
rect 32776 66340 32832 66396
rect 32832 66340 32836 66396
rect 32772 66336 32836 66340
rect 32852 66396 32916 66400
rect 32852 66340 32856 66396
rect 32856 66340 32912 66396
rect 32912 66340 32916 66396
rect 32852 66336 32916 66340
rect 37612 66396 37676 66400
rect 37612 66340 37616 66396
rect 37616 66340 37672 66396
rect 37672 66340 37676 66396
rect 37612 66336 37676 66340
rect 37692 66396 37756 66400
rect 37692 66340 37696 66396
rect 37696 66340 37752 66396
rect 37752 66340 37756 66396
rect 37692 66336 37756 66340
rect 37772 66396 37836 66400
rect 37772 66340 37776 66396
rect 37776 66340 37832 66396
rect 37832 66340 37836 66396
rect 37772 66336 37836 66340
rect 37852 66396 37916 66400
rect 37852 66340 37856 66396
rect 37856 66340 37912 66396
rect 37912 66340 37916 66396
rect 37852 66336 37916 66340
rect 1952 65852 2016 65856
rect 1952 65796 1956 65852
rect 1956 65796 2012 65852
rect 2012 65796 2016 65852
rect 1952 65792 2016 65796
rect 2032 65852 2096 65856
rect 2032 65796 2036 65852
rect 2036 65796 2092 65852
rect 2092 65796 2096 65852
rect 2032 65792 2096 65796
rect 2112 65852 2176 65856
rect 2112 65796 2116 65852
rect 2116 65796 2172 65852
rect 2172 65796 2176 65852
rect 2112 65792 2176 65796
rect 2192 65852 2256 65856
rect 2192 65796 2196 65852
rect 2196 65796 2252 65852
rect 2252 65796 2256 65852
rect 2192 65792 2256 65796
rect 6952 65852 7016 65856
rect 6952 65796 6956 65852
rect 6956 65796 7012 65852
rect 7012 65796 7016 65852
rect 6952 65792 7016 65796
rect 7032 65852 7096 65856
rect 7032 65796 7036 65852
rect 7036 65796 7092 65852
rect 7092 65796 7096 65852
rect 7032 65792 7096 65796
rect 7112 65852 7176 65856
rect 7112 65796 7116 65852
rect 7116 65796 7172 65852
rect 7172 65796 7176 65852
rect 7112 65792 7176 65796
rect 7192 65852 7256 65856
rect 7192 65796 7196 65852
rect 7196 65796 7252 65852
rect 7252 65796 7256 65852
rect 7192 65792 7256 65796
rect 11952 65852 12016 65856
rect 11952 65796 11956 65852
rect 11956 65796 12012 65852
rect 12012 65796 12016 65852
rect 11952 65792 12016 65796
rect 12032 65852 12096 65856
rect 12032 65796 12036 65852
rect 12036 65796 12092 65852
rect 12092 65796 12096 65852
rect 12032 65792 12096 65796
rect 12112 65852 12176 65856
rect 12112 65796 12116 65852
rect 12116 65796 12172 65852
rect 12172 65796 12176 65852
rect 12112 65792 12176 65796
rect 12192 65852 12256 65856
rect 12192 65796 12196 65852
rect 12196 65796 12252 65852
rect 12252 65796 12256 65852
rect 12192 65792 12256 65796
rect 16952 65852 17016 65856
rect 16952 65796 16956 65852
rect 16956 65796 17012 65852
rect 17012 65796 17016 65852
rect 16952 65792 17016 65796
rect 17032 65852 17096 65856
rect 17032 65796 17036 65852
rect 17036 65796 17092 65852
rect 17092 65796 17096 65852
rect 17032 65792 17096 65796
rect 17112 65852 17176 65856
rect 17112 65796 17116 65852
rect 17116 65796 17172 65852
rect 17172 65796 17176 65852
rect 17112 65792 17176 65796
rect 17192 65852 17256 65856
rect 17192 65796 17196 65852
rect 17196 65796 17252 65852
rect 17252 65796 17256 65852
rect 17192 65792 17256 65796
rect 21952 65852 22016 65856
rect 21952 65796 21956 65852
rect 21956 65796 22012 65852
rect 22012 65796 22016 65852
rect 21952 65792 22016 65796
rect 22032 65852 22096 65856
rect 22032 65796 22036 65852
rect 22036 65796 22092 65852
rect 22092 65796 22096 65852
rect 22032 65792 22096 65796
rect 22112 65852 22176 65856
rect 22112 65796 22116 65852
rect 22116 65796 22172 65852
rect 22172 65796 22176 65852
rect 22112 65792 22176 65796
rect 22192 65852 22256 65856
rect 22192 65796 22196 65852
rect 22196 65796 22252 65852
rect 22252 65796 22256 65852
rect 22192 65792 22256 65796
rect 26952 65852 27016 65856
rect 26952 65796 26956 65852
rect 26956 65796 27012 65852
rect 27012 65796 27016 65852
rect 26952 65792 27016 65796
rect 27032 65852 27096 65856
rect 27032 65796 27036 65852
rect 27036 65796 27092 65852
rect 27092 65796 27096 65852
rect 27032 65792 27096 65796
rect 27112 65852 27176 65856
rect 27112 65796 27116 65852
rect 27116 65796 27172 65852
rect 27172 65796 27176 65852
rect 27112 65792 27176 65796
rect 27192 65852 27256 65856
rect 27192 65796 27196 65852
rect 27196 65796 27252 65852
rect 27252 65796 27256 65852
rect 27192 65792 27256 65796
rect 31952 65852 32016 65856
rect 31952 65796 31956 65852
rect 31956 65796 32012 65852
rect 32012 65796 32016 65852
rect 31952 65792 32016 65796
rect 32032 65852 32096 65856
rect 32032 65796 32036 65852
rect 32036 65796 32092 65852
rect 32092 65796 32096 65852
rect 32032 65792 32096 65796
rect 32112 65852 32176 65856
rect 32112 65796 32116 65852
rect 32116 65796 32172 65852
rect 32172 65796 32176 65852
rect 32112 65792 32176 65796
rect 32192 65852 32256 65856
rect 32192 65796 32196 65852
rect 32196 65796 32252 65852
rect 32252 65796 32256 65852
rect 32192 65792 32256 65796
rect 36952 65852 37016 65856
rect 36952 65796 36956 65852
rect 36956 65796 37012 65852
rect 37012 65796 37016 65852
rect 36952 65792 37016 65796
rect 37032 65852 37096 65856
rect 37032 65796 37036 65852
rect 37036 65796 37092 65852
rect 37092 65796 37096 65852
rect 37032 65792 37096 65796
rect 37112 65852 37176 65856
rect 37112 65796 37116 65852
rect 37116 65796 37172 65852
rect 37172 65796 37176 65852
rect 37112 65792 37176 65796
rect 37192 65852 37256 65856
rect 37192 65796 37196 65852
rect 37196 65796 37252 65852
rect 37252 65796 37256 65852
rect 37192 65792 37256 65796
rect 23612 65452 23676 65516
rect 2612 65308 2676 65312
rect 2612 65252 2616 65308
rect 2616 65252 2672 65308
rect 2672 65252 2676 65308
rect 2612 65248 2676 65252
rect 2692 65308 2756 65312
rect 2692 65252 2696 65308
rect 2696 65252 2752 65308
rect 2752 65252 2756 65308
rect 2692 65248 2756 65252
rect 2772 65308 2836 65312
rect 2772 65252 2776 65308
rect 2776 65252 2832 65308
rect 2832 65252 2836 65308
rect 2772 65248 2836 65252
rect 2852 65308 2916 65312
rect 2852 65252 2856 65308
rect 2856 65252 2912 65308
rect 2912 65252 2916 65308
rect 2852 65248 2916 65252
rect 7612 65308 7676 65312
rect 7612 65252 7616 65308
rect 7616 65252 7672 65308
rect 7672 65252 7676 65308
rect 7612 65248 7676 65252
rect 7692 65308 7756 65312
rect 7692 65252 7696 65308
rect 7696 65252 7752 65308
rect 7752 65252 7756 65308
rect 7692 65248 7756 65252
rect 7772 65308 7836 65312
rect 7772 65252 7776 65308
rect 7776 65252 7832 65308
rect 7832 65252 7836 65308
rect 7772 65248 7836 65252
rect 7852 65308 7916 65312
rect 7852 65252 7856 65308
rect 7856 65252 7912 65308
rect 7912 65252 7916 65308
rect 7852 65248 7916 65252
rect 12612 65308 12676 65312
rect 12612 65252 12616 65308
rect 12616 65252 12672 65308
rect 12672 65252 12676 65308
rect 12612 65248 12676 65252
rect 12692 65308 12756 65312
rect 12692 65252 12696 65308
rect 12696 65252 12752 65308
rect 12752 65252 12756 65308
rect 12692 65248 12756 65252
rect 12772 65308 12836 65312
rect 12772 65252 12776 65308
rect 12776 65252 12832 65308
rect 12832 65252 12836 65308
rect 12772 65248 12836 65252
rect 12852 65308 12916 65312
rect 12852 65252 12856 65308
rect 12856 65252 12912 65308
rect 12912 65252 12916 65308
rect 12852 65248 12916 65252
rect 17612 65308 17676 65312
rect 17612 65252 17616 65308
rect 17616 65252 17672 65308
rect 17672 65252 17676 65308
rect 17612 65248 17676 65252
rect 17692 65308 17756 65312
rect 17692 65252 17696 65308
rect 17696 65252 17752 65308
rect 17752 65252 17756 65308
rect 17692 65248 17756 65252
rect 17772 65308 17836 65312
rect 17772 65252 17776 65308
rect 17776 65252 17832 65308
rect 17832 65252 17836 65308
rect 17772 65248 17836 65252
rect 17852 65308 17916 65312
rect 17852 65252 17856 65308
rect 17856 65252 17912 65308
rect 17912 65252 17916 65308
rect 17852 65248 17916 65252
rect 22612 65308 22676 65312
rect 22612 65252 22616 65308
rect 22616 65252 22672 65308
rect 22672 65252 22676 65308
rect 22612 65248 22676 65252
rect 22692 65308 22756 65312
rect 22692 65252 22696 65308
rect 22696 65252 22752 65308
rect 22752 65252 22756 65308
rect 22692 65248 22756 65252
rect 22772 65308 22836 65312
rect 22772 65252 22776 65308
rect 22776 65252 22832 65308
rect 22832 65252 22836 65308
rect 22772 65248 22836 65252
rect 22852 65308 22916 65312
rect 22852 65252 22856 65308
rect 22856 65252 22912 65308
rect 22912 65252 22916 65308
rect 22852 65248 22916 65252
rect 27612 65308 27676 65312
rect 27612 65252 27616 65308
rect 27616 65252 27672 65308
rect 27672 65252 27676 65308
rect 27612 65248 27676 65252
rect 27692 65308 27756 65312
rect 27692 65252 27696 65308
rect 27696 65252 27752 65308
rect 27752 65252 27756 65308
rect 27692 65248 27756 65252
rect 27772 65308 27836 65312
rect 27772 65252 27776 65308
rect 27776 65252 27832 65308
rect 27832 65252 27836 65308
rect 27772 65248 27836 65252
rect 27852 65308 27916 65312
rect 27852 65252 27856 65308
rect 27856 65252 27912 65308
rect 27912 65252 27916 65308
rect 27852 65248 27916 65252
rect 32612 65308 32676 65312
rect 32612 65252 32616 65308
rect 32616 65252 32672 65308
rect 32672 65252 32676 65308
rect 32612 65248 32676 65252
rect 32692 65308 32756 65312
rect 32692 65252 32696 65308
rect 32696 65252 32752 65308
rect 32752 65252 32756 65308
rect 32692 65248 32756 65252
rect 32772 65308 32836 65312
rect 32772 65252 32776 65308
rect 32776 65252 32832 65308
rect 32832 65252 32836 65308
rect 32772 65248 32836 65252
rect 32852 65308 32916 65312
rect 32852 65252 32856 65308
rect 32856 65252 32912 65308
rect 32912 65252 32916 65308
rect 32852 65248 32916 65252
rect 37612 65308 37676 65312
rect 37612 65252 37616 65308
rect 37616 65252 37672 65308
rect 37672 65252 37676 65308
rect 37612 65248 37676 65252
rect 37692 65308 37756 65312
rect 37692 65252 37696 65308
rect 37696 65252 37752 65308
rect 37752 65252 37756 65308
rect 37692 65248 37756 65252
rect 37772 65308 37836 65312
rect 37772 65252 37776 65308
rect 37776 65252 37832 65308
rect 37832 65252 37836 65308
rect 37772 65248 37836 65252
rect 37852 65308 37916 65312
rect 37852 65252 37856 65308
rect 37856 65252 37912 65308
rect 37912 65252 37916 65308
rect 37852 65248 37916 65252
rect 1952 64764 2016 64768
rect 1952 64708 1956 64764
rect 1956 64708 2012 64764
rect 2012 64708 2016 64764
rect 1952 64704 2016 64708
rect 2032 64764 2096 64768
rect 2032 64708 2036 64764
rect 2036 64708 2092 64764
rect 2092 64708 2096 64764
rect 2032 64704 2096 64708
rect 2112 64764 2176 64768
rect 2112 64708 2116 64764
rect 2116 64708 2172 64764
rect 2172 64708 2176 64764
rect 2112 64704 2176 64708
rect 2192 64764 2256 64768
rect 2192 64708 2196 64764
rect 2196 64708 2252 64764
rect 2252 64708 2256 64764
rect 2192 64704 2256 64708
rect 6952 64764 7016 64768
rect 6952 64708 6956 64764
rect 6956 64708 7012 64764
rect 7012 64708 7016 64764
rect 6952 64704 7016 64708
rect 7032 64764 7096 64768
rect 7032 64708 7036 64764
rect 7036 64708 7092 64764
rect 7092 64708 7096 64764
rect 7032 64704 7096 64708
rect 7112 64764 7176 64768
rect 7112 64708 7116 64764
rect 7116 64708 7172 64764
rect 7172 64708 7176 64764
rect 7112 64704 7176 64708
rect 7192 64764 7256 64768
rect 7192 64708 7196 64764
rect 7196 64708 7252 64764
rect 7252 64708 7256 64764
rect 7192 64704 7256 64708
rect 11952 64764 12016 64768
rect 11952 64708 11956 64764
rect 11956 64708 12012 64764
rect 12012 64708 12016 64764
rect 11952 64704 12016 64708
rect 12032 64764 12096 64768
rect 12032 64708 12036 64764
rect 12036 64708 12092 64764
rect 12092 64708 12096 64764
rect 12032 64704 12096 64708
rect 12112 64764 12176 64768
rect 12112 64708 12116 64764
rect 12116 64708 12172 64764
rect 12172 64708 12176 64764
rect 12112 64704 12176 64708
rect 12192 64764 12256 64768
rect 12192 64708 12196 64764
rect 12196 64708 12252 64764
rect 12252 64708 12256 64764
rect 12192 64704 12256 64708
rect 16952 64764 17016 64768
rect 16952 64708 16956 64764
rect 16956 64708 17012 64764
rect 17012 64708 17016 64764
rect 16952 64704 17016 64708
rect 17032 64764 17096 64768
rect 17032 64708 17036 64764
rect 17036 64708 17092 64764
rect 17092 64708 17096 64764
rect 17032 64704 17096 64708
rect 17112 64764 17176 64768
rect 17112 64708 17116 64764
rect 17116 64708 17172 64764
rect 17172 64708 17176 64764
rect 17112 64704 17176 64708
rect 17192 64764 17256 64768
rect 17192 64708 17196 64764
rect 17196 64708 17252 64764
rect 17252 64708 17256 64764
rect 17192 64704 17256 64708
rect 21952 64764 22016 64768
rect 21952 64708 21956 64764
rect 21956 64708 22012 64764
rect 22012 64708 22016 64764
rect 21952 64704 22016 64708
rect 22032 64764 22096 64768
rect 22032 64708 22036 64764
rect 22036 64708 22092 64764
rect 22092 64708 22096 64764
rect 22032 64704 22096 64708
rect 22112 64764 22176 64768
rect 22112 64708 22116 64764
rect 22116 64708 22172 64764
rect 22172 64708 22176 64764
rect 22112 64704 22176 64708
rect 22192 64764 22256 64768
rect 22192 64708 22196 64764
rect 22196 64708 22252 64764
rect 22252 64708 22256 64764
rect 22192 64704 22256 64708
rect 26952 64764 27016 64768
rect 26952 64708 26956 64764
rect 26956 64708 27012 64764
rect 27012 64708 27016 64764
rect 26952 64704 27016 64708
rect 27032 64764 27096 64768
rect 27032 64708 27036 64764
rect 27036 64708 27092 64764
rect 27092 64708 27096 64764
rect 27032 64704 27096 64708
rect 27112 64764 27176 64768
rect 27112 64708 27116 64764
rect 27116 64708 27172 64764
rect 27172 64708 27176 64764
rect 27112 64704 27176 64708
rect 27192 64764 27256 64768
rect 27192 64708 27196 64764
rect 27196 64708 27252 64764
rect 27252 64708 27256 64764
rect 27192 64704 27256 64708
rect 31952 64764 32016 64768
rect 31952 64708 31956 64764
rect 31956 64708 32012 64764
rect 32012 64708 32016 64764
rect 31952 64704 32016 64708
rect 32032 64764 32096 64768
rect 32032 64708 32036 64764
rect 32036 64708 32092 64764
rect 32092 64708 32096 64764
rect 32032 64704 32096 64708
rect 32112 64764 32176 64768
rect 32112 64708 32116 64764
rect 32116 64708 32172 64764
rect 32172 64708 32176 64764
rect 32112 64704 32176 64708
rect 32192 64764 32256 64768
rect 32192 64708 32196 64764
rect 32196 64708 32252 64764
rect 32252 64708 32256 64764
rect 32192 64704 32256 64708
rect 36952 64764 37016 64768
rect 36952 64708 36956 64764
rect 36956 64708 37012 64764
rect 37012 64708 37016 64764
rect 36952 64704 37016 64708
rect 37032 64764 37096 64768
rect 37032 64708 37036 64764
rect 37036 64708 37092 64764
rect 37092 64708 37096 64764
rect 37032 64704 37096 64708
rect 37112 64764 37176 64768
rect 37112 64708 37116 64764
rect 37116 64708 37172 64764
rect 37172 64708 37176 64764
rect 37112 64704 37176 64708
rect 37192 64764 37256 64768
rect 37192 64708 37196 64764
rect 37196 64708 37252 64764
rect 37252 64708 37256 64764
rect 37192 64704 37256 64708
rect 2612 64220 2676 64224
rect 2612 64164 2616 64220
rect 2616 64164 2672 64220
rect 2672 64164 2676 64220
rect 2612 64160 2676 64164
rect 2692 64220 2756 64224
rect 2692 64164 2696 64220
rect 2696 64164 2752 64220
rect 2752 64164 2756 64220
rect 2692 64160 2756 64164
rect 2772 64220 2836 64224
rect 2772 64164 2776 64220
rect 2776 64164 2832 64220
rect 2832 64164 2836 64220
rect 2772 64160 2836 64164
rect 2852 64220 2916 64224
rect 2852 64164 2856 64220
rect 2856 64164 2912 64220
rect 2912 64164 2916 64220
rect 2852 64160 2916 64164
rect 7612 64220 7676 64224
rect 7612 64164 7616 64220
rect 7616 64164 7672 64220
rect 7672 64164 7676 64220
rect 7612 64160 7676 64164
rect 7692 64220 7756 64224
rect 7692 64164 7696 64220
rect 7696 64164 7752 64220
rect 7752 64164 7756 64220
rect 7692 64160 7756 64164
rect 7772 64220 7836 64224
rect 7772 64164 7776 64220
rect 7776 64164 7832 64220
rect 7832 64164 7836 64220
rect 7772 64160 7836 64164
rect 7852 64220 7916 64224
rect 7852 64164 7856 64220
rect 7856 64164 7912 64220
rect 7912 64164 7916 64220
rect 7852 64160 7916 64164
rect 12612 64220 12676 64224
rect 12612 64164 12616 64220
rect 12616 64164 12672 64220
rect 12672 64164 12676 64220
rect 12612 64160 12676 64164
rect 12692 64220 12756 64224
rect 12692 64164 12696 64220
rect 12696 64164 12752 64220
rect 12752 64164 12756 64220
rect 12692 64160 12756 64164
rect 12772 64220 12836 64224
rect 12772 64164 12776 64220
rect 12776 64164 12832 64220
rect 12832 64164 12836 64220
rect 12772 64160 12836 64164
rect 12852 64220 12916 64224
rect 12852 64164 12856 64220
rect 12856 64164 12912 64220
rect 12912 64164 12916 64220
rect 12852 64160 12916 64164
rect 17612 64220 17676 64224
rect 17612 64164 17616 64220
rect 17616 64164 17672 64220
rect 17672 64164 17676 64220
rect 17612 64160 17676 64164
rect 17692 64220 17756 64224
rect 17692 64164 17696 64220
rect 17696 64164 17752 64220
rect 17752 64164 17756 64220
rect 17692 64160 17756 64164
rect 17772 64220 17836 64224
rect 17772 64164 17776 64220
rect 17776 64164 17832 64220
rect 17832 64164 17836 64220
rect 17772 64160 17836 64164
rect 17852 64220 17916 64224
rect 17852 64164 17856 64220
rect 17856 64164 17912 64220
rect 17912 64164 17916 64220
rect 17852 64160 17916 64164
rect 22612 64220 22676 64224
rect 22612 64164 22616 64220
rect 22616 64164 22672 64220
rect 22672 64164 22676 64220
rect 22612 64160 22676 64164
rect 22692 64220 22756 64224
rect 22692 64164 22696 64220
rect 22696 64164 22752 64220
rect 22752 64164 22756 64220
rect 22692 64160 22756 64164
rect 22772 64220 22836 64224
rect 22772 64164 22776 64220
rect 22776 64164 22832 64220
rect 22832 64164 22836 64220
rect 22772 64160 22836 64164
rect 22852 64220 22916 64224
rect 22852 64164 22856 64220
rect 22856 64164 22912 64220
rect 22912 64164 22916 64220
rect 22852 64160 22916 64164
rect 27612 64220 27676 64224
rect 27612 64164 27616 64220
rect 27616 64164 27672 64220
rect 27672 64164 27676 64220
rect 27612 64160 27676 64164
rect 27692 64220 27756 64224
rect 27692 64164 27696 64220
rect 27696 64164 27752 64220
rect 27752 64164 27756 64220
rect 27692 64160 27756 64164
rect 27772 64220 27836 64224
rect 27772 64164 27776 64220
rect 27776 64164 27832 64220
rect 27832 64164 27836 64220
rect 27772 64160 27836 64164
rect 27852 64220 27916 64224
rect 27852 64164 27856 64220
rect 27856 64164 27912 64220
rect 27912 64164 27916 64220
rect 27852 64160 27916 64164
rect 32612 64220 32676 64224
rect 32612 64164 32616 64220
rect 32616 64164 32672 64220
rect 32672 64164 32676 64220
rect 32612 64160 32676 64164
rect 32692 64220 32756 64224
rect 32692 64164 32696 64220
rect 32696 64164 32752 64220
rect 32752 64164 32756 64220
rect 32692 64160 32756 64164
rect 32772 64220 32836 64224
rect 32772 64164 32776 64220
rect 32776 64164 32832 64220
rect 32832 64164 32836 64220
rect 32772 64160 32836 64164
rect 32852 64220 32916 64224
rect 32852 64164 32856 64220
rect 32856 64164 32912 64220
rect 32912 64164 32916 64220
rect 32852 64160 32916 64164
rect 37612 64220 37676 64224
rect 37612 64164 37616 64220
rect 37616 64164 37672 64220
rect 37672 64164 37676 64220
rect 37612 64160 37676 64164
rect 37692 64220 37756 64224
rect 37692 64164 37696 64220
rect 37696 64164 37752 64220
rect 37752 64164 37756 64220
rect 37692 64160 37756 64164
rect 37772 64220 37836 64224
rect 37772 64164 37776 64220
rect 37776 64164 37832 64220
rect 37832 64164 37836 64220
rect 37772 64160 37836 64164
rect 37852 64220 37916 64224
rect 37852 64164 37856 64220
rect 37856 64164 37912 64220
rect 37912 64164 37916 64220
rect 37852 64160 37916 64164
rect 1952 63676 2016 63680
rect 1952 63620 1956 63676
rect 1956 63620 2012 63676
rect 2012 63620 2016 63676
rect 1952 63616 2016 63620
rect 2032 63676 2096 63680
rect 2032 63620 2036 63676
rect 2036 63620 2092 63676
rect 2092 63620 2096 63676
rect 2032 63616 2096 63620
rect 2112 63676 2176 63680
rect 2112 63620 2116 63676
rect 2116 63620 2172 63676
rect 2172 63620 2176 63676
rect 2112 63616 2176 63620
rect 2192 63676 2256 63680
rect 2192 63620 2196 63676
rect 2196 63620 2252 63676
rect 2252 63620 2256 63676
rect 2192 63616 2256 63620
rect 6952 63676 7016 63680
rect 6952 63620 6956 63676
rect 6956 63620 7012 63676
rect 7012 63620 7016 63676
rect 6952 63616 7016 63620
rect 7032 63676 7096 63680
rect 7032 63620 7036 63676
rect 7036 63620 7092 63676
rect 7092 63620 7096 63676
rect 7032 63616 7096 63620
rect 7112 63676 7176 63680
rect 7112 63620 7116 63676
rect 7116 63620 7172 63676
rect 7172 63620 7176 63676
rect 7112 63616 7176 63620
rect 7192 63676 7256 63680
rect 7192 63620 7196 63676
rect 7196 63620 7252 63676
rect 7252 63620 7256 63676
rect 7192 63616 7256 63620
rect 11952 63676 12016 63680
rect 11952 63620 11956 63676
rect 11956 63620 12012 63676
rect 12012 63620 12016 63676
rect 11952 63616 12016 63620
rect 12032 63676 12096 63680
rect 12032 63620 12036 63676
rect 12036 63620 12092 63676
rect 12092 63620 12096 63676
rect 12032 63616 12096 63620
rect 12112 63676 12176 63680
rect 12112 63620 12116 63676
rect 12116 63620 12172 63676
rect 12172 63620 12176 63676
rect 12112 63616 12176 63620
rect 12192 63676 12256 63680
rect 12192 63620 12196 63676
rect 12196 63620 12252 63676
rect 12252 63620 12256 63676
rect 12192 63616 12256 63620
rect 16952 63676 17016 63680
rect 16952 63620 16956 63676
rect 16956 63620 17012 63676
rect 17012 63620 17016 63676
rect 16952 63616 17016 63620
rect 17032 63676 17096 63680
rect 17032 63620 17036 63676
rect 17036 63620 17092 63676
rect 17092 63620 17096 63676
rect 17032 63616 17096 63620
rect 17112 63676 17176 63680
rect 17112 63620 17116 63676
rect 17116 63620 17172 63676
rect 17172 63620 17176 63676
rect 17112 63616 17176 63620
rect 17192 63676 17256 63680
rect 17192 63620 17196 63676
rect 17196 63620 17252 63676
rect 17252 63620 17256 63676
rect 17192 63616 17256 63620
rect 21952 63676 22016 63680
rect 21952 63620 21956 63676
rect 21956 63620 22012 63676
rect 22012 63620 22016 63676
rect 21952 63616 22016 63620
rect 22032 63676 22096 63680
rect 22032 63620 22036 63676
rect 22036 63620 22092 63676
rect 22092 63620 22096 63676
rect 22032 63616 22096 63620
rect 22112 63676 22176 63680
rect 22112 63620 22116 63676
rect 22116 63620 22172 63676
rect 22172 63620 22176 63676
rect 22112 63616 22176 63620
rect 22192 63676 22256 63680
rect 22192 63620 22196 63676
rect 22196 63620 22252 63676
rect 22252 63620 22256 63676
rect 22192 63616 22256 63620
rect 26952 63676 27016 63680
rect 26952 63620 26956 63676
rect 26956 63620 27012 63676
rect 27012 63620 27016 63676
rect 26952 63616 27016 63620
rect 27032 63676 27096 63680
rect 27032 63620 27036 63676
rect 27036 63620 27092 63676
rect 27092 63620 27096 63676
rect 27032 63616 27096 63620
rect 27112 63676 27176 63680
rect 27112 63620 27116 63676
rect 27116 63620 27172 63676
rect 27172 63620 27176 63676
rect 27112 63616 27176 63620
rect 27192 63676 27256 63680
rect 27192 63620 27196 63676
rect 27196 63620 27252 63676
rect 27252 63620 27256 63676
rect 27192 63616 27256 63620
rect 31952 63676 32016 63680
rect 31952 63620 31956 63676
rect 31956 63620 32012 63676
rect 32012 63620 32016 63676
rect 31952 63616 32016 63620
rect 32032 63676 32096 63680
rect 32032 63620 32036 63676
rect 32036 63620 32092 63676
rect 32092 63620 32096 63676
rect 32032 63616 32096 63620
rect 32112 63676 32176 63680
rect 32112 63620 32116 63676
rect 32116 63620 32172 63676
rect 32172 63620 32176 63676
rect 32112 63616 32176 63620
rect 32192 63676 32256 63680
rect 32192 63620 32196 63676
rect 32196 63620 32252 63676
rect 32252 63620 32256 63676
rect 32192 63616 32256 63620
rect 36952 63676 37016 63680
rect 36952 63620 36956 63676
rect 36956 63620 37012 63676
rect 37012 63620 37016 63676
rect 36952 63616 37016 63620
rect 37032 63676 37096 63680
rect 37032 63620 37036 63676
rect 37036 63620 37092 63676
rect 37092 63620 37096 63676
rect 37032 63616 37096 63620
rect 37112 63676 37176 63680
rect 37112 63620 37116 63676
rect 37116 63620 37172 63676
rect 37172 63620 37176 63676
rect 37112 63616 37176 63620
rect 37192 63676 37256 63680
rect 37192 63620 37196 63676
rect 37196 63620 37252 63676
rect 37252 63620 37256 63676
rect 37192 63616 37256 63620
rect 20484 63548 20548 63612
rect 21588 63548 21652 63612
rect 2612 63132 2676 63136
rect 2612 63076 2616 63132
rect 2616 63076 2672 63132
rect 2672 63076 2676 63132
rect 2612 63072 2676 63076
rect 2692 63132 2756 63136
rect 2692 63076 2696 63132
rect 2696 63076 2752 63132
rect 2752 63076 2756 63132
rect 2692 63072 2756 63076
rect 2772 63132 2836 63136
rect 2772 63076 2776 63132
rect 2776 63076 2832 63132
rect 2832 63076 2836 63132
rect 2772 63072 2836 63076
rect 2852 63132 2916 63136
rect 2852 63076 2856 63132
rect 2856 63076 2912 63132
rect 2912 63076 2916 63132
rect 2852 63072 2916 63076
rect 7612 63132 7676 63136
rect 7612 63076 7616 63132
rect 7616 63076 7672 63132
rect 7672 63076 7676 63132
rect 7612 63072 7676 63076
rect 7692 63132 7756 63136
rect 7692 63076 7696 63132
rect 7696 63076 7752 63132
rect 7752 63076 7756 63132
rect 7692 63072 7756 63076
rect 7772 63132 7836 63136
rect 7772 63076 7776 63132
rect 7776 63076 7832 63132
rect 7832 63076 7836 63132
rect 7772 63072 7836 63076
rect 7852 63132 7916 63136
rect 7852 63076 7856 63132
rect 7856 63076 7912 63132
rect 7912 63076 7916 63132
rect 7852 63072 7916 63076
rect 12612 63132 12676 63136
rect 12612 63076 12616 63132
rect 12616 63076 12672 63132
rect 12672 63076 12676 63132
rect 12612 63072 12676 63076
rect 12692 63132 12756 63136
rect 12692 63076 12696 63132
rect 12696 63076 12752 63132
rect 12752 63076 12756 63132
rect 12692 63072 12756 63076
rect 12772 63132 12836 63136
rect 12772 63076 12776 63132
rect 12776 63076 12832 63132
rect 12832 63076 12836 63132
rect 12772 63072 12836 63076
rect 12852 63132 12916 63136
rect 12852 63076 12856 63132
rect 12856 63076 12912 63132
rect 12912 63076 12916 63132
rect 12852 63072 12916 63076
rect 17612 63132 17676 63136
rect 17612 63076 17616 63132
rect 17616 63076 17672 63132
rect 17672 63076 17676 63132
rect 17612 63072 17676 63076
rect 17692 63132 17756 63136
rect 17692 63076 17696 63132
rect 17696 63076 17752 63132
rect 17752 63076 17756 63132
rect 17692 63072 17756 63076
rect 17772 63132 17836 63136
rect 17772 63076 17776 63132
rect 17776 63076 17832 63132
rect 17832 63076 17836 63132
rect 17772 63072 17836 63076
rect 17852 63132 17916 63136
rect 17852 63076 17856 63132
rect 17856 63076 17912 63132
rect 17912 63076 17916 63132
rect 17852 63072 17916 63076
rect 22612 63132 22676 63136
rect 22612 63076 22616 63132
rect 22616 63076 22672 63132
rect 22672 63076 22676 63132
rect 22612 63072 22676 63076
rect 22692 63132 22756 63136
rect 22692 63076 22696 63132
rect 22696 63076 22752 63132
rect 22752 63076 22756 63132
rect 22692 63072 22756 63076
rect 22772 63132 22836 63136
rect 22772 63076 22776 63132
rect 22776 63076 22832 63132
rect 22832 63076 22836 63132
rect 22772 63072 22836 63076
rect 22852 63132 22916 63136
rect 22852 63076 22856 63132
rect 22856 63076 22912 63132
rect 22912 63076 22916 63132
rect 22852 63072 22916 63076
rect 27612 63132 27676 63136
rect 27612 63076 27616 63132
rect 27616 63076 27672 63132
rect 27672 63076 27676 63132
rect 27612 63072 27676 63076
rect 27692 63132 27756 63136
rect 27692 63076 27696 63132
rect 27696 63076 27752 63132
rect 27752 63076 27756 63132
rect 27692 63072 27756 63076
rect 27772 63132 27836 63136
rect 27772 63076 27776 63132
rect 27776 63076 27832 63132
rect 27832 63076 27836 63132
rect 27772 63072 27836 63076
rect 27852 63132 27916 63136
rect 27852 63076 27856 63132
rect 27856 63076 27912 63132
rect 27912 63076 27916 63132
rect 27852 63072 27916 63076
rect 32612 63132 32676 63136
rect 32612 63076 32616 63132
rect 32616 63076 32672 63132
rect 32672 63076 32676 63132
rect 32612 63072 32676 63076
rect 32692 63132 32756 63136
rect 32692 63076 32696 63132
rect 32696 63076 32752 63132
rect 32752 63076 32756 63132
rect 32692 63072 32756 63076
rect 32772 63132 32836 63136
rect 32772 63076 32776 63132
rect 32776 63076 32832 63132
rect 32832 63076 32836 63132
rect 32772 63072 32836 63076
rect 32852 63132 32916 63136
rect 32852 63076 32856 63132
rect 32856 63076 32912 63132
rect 32912 63076 32916 63132
rect 32852 63072 32916 63076
rect 37612 63132 37676 63136
rect 37612 63076 37616 63132
rect 37616 63076 37672 63132
rect 37672 63076 37676 63132
rect 37612 63072 37676 63076
rect 37692 63132 37756 63136
rect 37692 63076 37696 63132
rect 37696 63076 37752 63132
rect 37752 63076 37756 63132
rect 37692 63072 37756 63076
rect 37772 63132 37836 63136
rect 37772 63076 37776 63132
rect 37776 63076 37832 63132
rect 37832 63076 37836 63132
rect 37772 63072 37836 63076
rect 37852 63132 37916 63136
rect 37852 63076 37856 63132
rect 37856 63076 37912 63132
rect 37912 63076 37916 63132
rect 37852 63072 37916 63076
rect 24716 62732 24780 62796
rect 1952 62588 2016 62592
rect 1952 62532 1956 62588
rect 1956 62532 2012 62588
rect 2012 62532 2016 62588
rect 1952 62528 2016 62532
rect 2032 62588 2096 62592
rect 2032 62532 2036 62588
rect 2036 62532 2092 62588
rect 2092 62532 2096 62588
rect 2032 62528 2096 62532
rect 2112 62588 2176 62592
rect 2112 62532 2116 62588
rect 2116 62532 2172 62588
rect 2172 62532 2176 62588
rect 2112 62528 2176 62532
rect 2192 62588 2256 62592
rect 2192 62532 2196 62588
rect 2196 62532 2252 62588
rect 2252 62532 2256 62588
rect 2192 62528 2256 62532
rect 6952 62588 7016 62592
rect 6952 62532 6956 62588
rect 6956 62532 7012 62588
rect 7012 62532 7016 62588
rect 6952 62528 7016 62532
rect 7032 62588 7096 62592
rect 7032 62532 7036 62588
rect 7036 62532 7092 62588
rect 7092 62532 7096 62588
rect 7032 62528 7096 62532
rect 7112 62588 7176 62592
rect 7112 62532 7116 62588
rect 7116 62532 7172 62588
rect 7172 62532 7176 62588
rect 7112 62528 7176 62532
rect 7192 62588 7256 62592
rect 7192 62532 7196 62588
rect 7196 62532 7252 62588
rect 7252 62532 7256 62588
rect 7192 62528 7256 62532
rect 11952 62588 12016 62592
rect 11952 62532 11956 62588
rect 11956 62532 12012 62588
rect 12012 62532 12016 62588
rect 11952 62528 12016 62532
rect 12032 62588 12096 62592
rect 12032 62532 12036 62588
rect 12036 62532 12092 62588
rect 12092 62532 12096 62588
rect 12032 62528 12096 62532
rect 12112 62588 12176 62592
rect 12112 62532 12116 62588
rect 12116 62532 12172 62588
rect 12172 62532 12176 62588
rect 12112 62528 12176 62532
rect 12192 62588 12256 62592
rect 12192 62532 12196 62588
rect 12196 62532 12252 62588
rect 12252 62532 12256 62588
rect 12192 62528 12256 62532
rect 16952 62588 17016 62592
rect 16952 62532 16956 62588
rect 16956 62532 17012 62588
rect 17012 62532 17016 62588
rect 16952 62528 17016 62532
rect 17032 62588 17096 62592
rect 17032 62532 17036 62588
rect 17036 62532 17092 62588
rect 17092 62532 17096 62588
rect 17032 62528 17096 62532
rect 17112 62588 17176 62592
rect 17112 62532 17116 62588
rect 17116 62532 17172 62588
rect 17172 62532 17176 62588
rect 17112 62528 17176 62532
rect 17192 62588 17256 62592
rect 17192 62532 17196 62588
rect 17196 62532 17252 62588
rect 17252 62532 17256 62588
rect 17192 62528 17256 62532
rect 21952 62588 22016 62592
rect 21952 62532 21956 62588
rect 21956 62532 22012 62588
rect 22012 62532 22016 62588
rect 21952 62528 22016 62532
rect 22032 62588 22096 62592
rect 22032 62532 22036 62588
rect 22036 62532 22092 62588
rect 22092 62532 22096 62588
rect 22032 62528 22096 62532
rect 22112 62588 22176 62592
rect 22112 62532 22116 62588
rect 22116 62532 22172 62588
rect 22172 62532 22176 62588
rect 22112 62528 22176 62532
rect 22192 62588 22256 62592
rect 22192 62532 22196 62588
rect 22196 62532 22252 62588
rect 22252 62532 22256 62588
rect 22192 62528 22256 62532
rect 26952 62588 27016 62592
rect 26952 62532 26956 62588
rect 26956 62532 27012 62588
rect 27012 62532 27016 62588
rect 26952 62528 27016 62532
rect 27032 62588 27096 62592
rect 27032 62532 27036 62588
rect 27036 62532 27092 62588
rect 27092 62532 27096 62588
rect 27032 62528 27096 62532
rect 27112 62588 27176 62592
rect 27112 62532 27116 62588
rect 27116 62532 27172 62588
rect 27172 62532 27176 62588
rect 27112 62528 27176 62532
rect 27192 62588 27256 62592
rect 27192 62532 27196 62588
rect 27196 62532 27252 62588
rect 27252 62532 27256 62588
rect 27192 62528 27256 62532
rect 31952 62588 32016 62592
rect 31952 62532 31956 62588
rect 31956 62532 32012 62588
rect 32012 62532 32016 62588
rect 31952 62528 32016 62532
rect 32032 62588 32096 62592
rect 32032 62532 32036 62588
rect 32036 62532 32092 62588
rect 32092 62532 32096 62588
rect 32032 62528 32096 62532
rect 32112 62588 32176 62592
rect 32112 62532 32116 62588
rect 32116 62532 32172 62588
rect 32172 62532 32176 62588
rect 32112 62528 32176 62532
rect 32192 62588 32256 62592
rect 32192 62532 32196 62588
rect 32196 62532 32252 62588
rect 32252 62532 32256 62588
rect 32192 62528 32256 62532
rect 36952 62588 37016 62592
rect 36952 62532 36956 62588
rect 36956 62532 37012 62588
rect 37012 62532 37016 62588
rect 36952 62528 37016 62532
rect 37032 62588 37096 62592
rect 37032 62532 37036 62588
rect 37036 62532 37092 62588
rect 37092 62532 37096 62588
rect 37032 62528 37096 62532
rect 37112 62588 37176 62592
rect 37112 62532 37116 62588
rect 37116 62532 37172 62588
rect 37172 62532 37176 62588
rect 37112 62528 37176 62532
rect 37192 62588 37256 62592
rect 37192 62532 37196 62588
rect 37196 62532 37252 62588
rect 37252 62532 37256 62588
rect 37192 62528 37256 62532
rect 2612 62044 2676 62048
rect 2612 61988 2616 62044
rect 2616 61988 2672 62044
rect 2672 61988 2676 62044
rect 2612 61984 2676 61988
rect 2692 62044 2756 62048
rect 2692 61988 2696 62044
rect 2696 61988 2752 62044
rect 2752 61988 2756 62044
rect 2692 61984 2756 61988
rect 2772 62044 2836 62048
rect 2772 61988 2776 62044
rect 2776 61988 2832 62044
rect 2832 61988 2836 62044
rect 2772 61984 2836 61988
rect 2852 62044 2916 62048
rect 2852 61988 2856 62044
rect 2856 61988 2912 62044
rect 2912 61988 2916 62044
rect 2852 61984 2916 61988
rect 7612 62044 7676 62048
rect 7612 61988 7616 62044
rect 7616 61988 7672 62044
rect 7672 61988 7676 62044
rect 7612 61984 7676 61988
rect 7692 62044 7756 62048
rect 7692 61988 7696 62044
rect 7696 61988 7752 62044
rect 7752 61988 7756 62044
rect 7692 61984 7756 61988
rect 7772 62044 7836 62048
rect 7772 61988 7776 62044
rect 7776 61988 7832 62044
rect 7832 61988 7836 62044
rect 7772 61984 7836 61988
rect 7852 62044 7916 62048
rect 7852 61988 7856 62044
rect 7856 61988 7912 62044
rect 7912 61988 7916 62044
rect 7852 61984 7916 61988
rect 12612 62044 12676 62048
rect 12612 61988 12616 62044
rect 12616 61988 12672 62044
rect 12672 61988 12676 62044
rect 12612 61984 12676 61988
rect 12692 62044 12756 62048
rect 12692 61988 12696 62044
rect 12696 61988 12752 62044
rect 12752 61988 12756 62044
rect 12692 61984 12756 61988
rect 12772 62044 12836 62048
rect 12772 61988 12776 62044
rect 12776 61988 12832 62044
rect 12832 61988 12836 62044
rect 12772 61984 12836 61988
rect 12852 62044 12916 62048
rect 12852 61988 12856 62044
rect 12856 61988 12912 62044
rect 12912 61988 12916 62044
rect 12852 61984 12916 61988
rect 17612 62044 17676 62048
rect 17612 61988 17616 62044
rect 17616 61988 17672 62044
rect 17672 61988 17676 62044
rect 17612 61984 17676 61988
rect 17692 62044 17756 62048
rect 17692 61988 17696 62044
rect 17696 61988 17752 62044
rect 17752 61988 17756 62044
rect 17692 61984 17756 61988
rect 17772 62044 17836 62048
rect 17772 61988 17776 62044
rect 17776 61988 17832 62044
rect 17832 61988 17836 62044
rect 17772 61984 17836 61988
rect 17852 62044 17916 62048
rect 17852 61988 17856 62044
rect 17856 61988 17912 62044
rect 17912 61988 17916 62044
rect 17852 61984 17916 61988
rect 22612 62044 22676 62048
rect 22612 61988 22616 62044
rect 22616 61988 22672 62044
rect 22672 61988 22676 62044
rect 22612 61984 22676 61988
rect 22692 62044 22756 62048
rect 22692 61988 22696 62044
rect 22696 61988 22752 62044
rect 22752 61988 22756 62044
rect 22692 61984 22756 61988
rect 22772 62044 22836 62048
rect 22772 61988 22776 62044
rect 22776 61988 22832 62044
rect 22832 61988 22836 62044
rect 22772 61984 22836 61988
rect 22852 62044 22916 62048
rect 22852 61988 22856 62044
rect 22856 61988 22912 62044
rect 22912 61988 22916 62044
rect 22852 61984 22916 61988
rect 27612 62044 27676 62048
rect 27612 61988 27616 62044
rect 27616 61988 27672 62044
rect 27672 61988 27676 62044
rect 27612 61984 27676 61988
rect 27692 62044 27756 62048
rect 27692 61988 27696 62044
rect 27696 61988 27752 62044
rect 27752 61988 27756 62044
rect 27692 61984 27756 61988
rect 27772 62044 27836 62048
rect 27772 61988 27776 62044
rect 27776 61988 27832 62044
rect 27832 61988 27836 62044
rect 27772 61984 27836 61988
rect 27852 62044 27916 62048
rect 27852 61988 27856 62044
rect 27856 61988 27912 62044
rect 27912 61988 27916 62044
rect 27852 61984 27916 61988
rect 32612 62044 32676 62048
rect 32612 61988 32616 62044
rect 32616 61988 32672 62044
rect 32672 61988 32676 62044
rect 32612 61984 32676 61988
rect 32692 62044 32756 62048
rect 32692 61988 32696 62044
rect 32696 61988 32752 62044
rect 32752 61988 32756 62044
rect 32692 61984 32756 61988
rect 32772 62044 32836 62048
rect 32772 61988 32776 62044
rect 32776 61988 32832 62044
rect 32832 61988 32836 62044
rect 32772 61984 32836 61988
rect 32852 62044 32916 62048
rect 32852 61988 32856 62044
rect 32856 61988 32912 62044
rect 32912 61988 32916 62044
rect 32852 61984 32916 61988
rect 37612 62044 37676 62048
rect 37612 61988 37616 62044
rect 37616 61988 37672 62044
rect 37672 61988 37676 62044
rect 37612 61984 37676 61988
rect 37692 62044 37756 62048
rect 37692 61988 37696 62044
rect 37696 61988 37752 62044
rect 37752 61988 37756 62044
rect 37692 61984 37756 61988
rect 37772 62044 37836 62048
rect 37772 61988 37776 62044
rect 37776 61988 37832 62044
rect 37832 61988 37836 62044
rect 37772 61984 37836 61988
rect 37852 62044 37916 62048
rect 37852 61988 37856 62044
rect 37856 61988 37912 62044
rect 37912 61988 37916 62044
rect 37852 61984 37916 61988
rect 25268 61644 25332 61708
rect 1952 61500 2016 61504
rect 1952 61444 1956 61500
rect 1956 61444 2012 61500
rect 2012 61444 2016 61500
rect 1952 61440 2016 61444
rect 2032 61500 2096 61504
rect 2032 61444 2036 61500
rect 2036 61444 2092 61500
rect 2092 61444 2096 61500
rect 2032 61440 2096 61444
rect 2112 61500 2176 61504
rect 2112 61444 2116 61500
rect 2116 61444 2172 61500
rect 2172 61444 2176 61500
rect 2112 61440 2176 61444
rect 2192 61500 2256 61504
rect 2192 61444 2196 61500
rect 2196 61444 2252 61500
rect 2252 61444 2256 61500
rect 2192 61440 2256 61444
rect 6952 61500 7016 61504
rect 6952 61444 6956 61500
rect 6956 61444 7012 61500
rect 7012 61444 7016 61500
rect 6952 61440 7016 61444
rect 7032 61500 7096 61504
rect 7032 61444 7036 61500
rect 7036 61444 7092 61500
rect 7092 61444 7096 61500
rect 7032 61440 7096 61444
rect 7112 61500 7176 61504
rect 7112 61444 7116 61500
rect 7116 61444 7172 61500
rect 7172 61444 7176 61500
rect 7112 61440 7176 61444
rect 7192 61500 7256 61504
rect 7192 61444 7196 61500
rect 7196 61444 7252 61500
rect 7252 61444 7256 61500
rect 7192 61440 7256 61444
rect 11952 61500 12016 61504
rect 11952 61444 11956 61500
rect 11956 61444 12012 61500
rect 12012 61444 12016 61500
rect 11952 61440 12016 61444
rect 12032 61500 12096 61504
rect 12032 61444 12036 61500
rect 12036 61444 12092 61500
rect 12092 61444 12096 61500
rect 12032 61440 12096 61444
rect 12112 61500 12176 61504
rect 12112 61444 12116 61500
rect 12116 61444 12172 61500
rect 12172 61444 12176 61500
rect 12112 61440 12176 61444
rect 12192 61500 12256 61504
rect 12192 61444 12196 61500
rect 12196 61444 12252 61500
rect 12252 61444 12256 61500
rect 12192 61440 12256 61444
rect 16952 61500 17016 61504
rect 16952 61444 16956 61500
rect 16956 61444 17012 61500
rect 17012 61444 17016 61500
rect 16952 61440 17016 61444
rect 17032 61500 17096 61504
rect 17032 61444 17036 61500
rect 17036 61444 17092 61500
rect 17092 61444 17096 61500
rect 17032 61440 17096 61444
rect 17112 61500 17176 61504
rect 17112 61444 17116 61500
rect 17116 61444 17172 61500
rect 17172 61444 17176 61500
rect 17112 61440 17176 61444
rect 17192 61500 17256 61504
rect 17192 61444 17196 61500
rect 17196 61444 17252 61500
rect 17252 61444 17256 61500
rect 17192 61440 17256 61444
rect 21952 61500 22016 61504
rect 21952 61444 21956 61500
rect 21956 61444 22012 61500
rect 22012 61444 22016 61500
rect 21952 61440 22016 61444
rect 22032 61500 22096 61504
rect 22032 61444 22036 61500
rect 22036 61444 22092 61500
rect 22092 61444 22096 61500
rect 22032 61440 22096 61444
rect 22112 61500 22176 61504
rect 22112 61444 22116 61500
rect 22116 61444 22172 61500
rect 22172 61444 22176 61500
rect 22112 61440 22176 61444
rect 22192 61500 22256 61504
rect 22192 61444 22196 61500
rect 22196 61444 22252 61500
rect 22252 61444 22256 61500
rect 22192 61440 22256 61444
rect 26952 61500 27016 61504
rect 26952 61444 26956 61500
rect 26956 61444 27012 61500
rect 27012 61444 27016 61500
rect 26952 61440 27016 61444
rect 27032 61500 27096 61504
rect 27032 61444 27036 61500
rect 27036 61444 27092 61500
rect 27092 61444 27096 61500
rect 27032 61440 27096 61444
rect 27112 61500 27176 61504
rect 27112 61444 27116 61500
rect 27116 61444 27172 61500
rect 27172 61444 27176 61500
rect 27112 61440 27176 61444
rect 27192 61500 27256 61504
rect 27192 61444 27196 61500
rect 27196 61444 27252 61500
rect 27252 61444 27256 61500
rect 27192 61440 27256 61444
rect 31952 61500 32016 61504
rect 31952 61444 31956 61500
rect 31956 61444 32012 61500
rect 32012 61444 32016 61500
rect 31952 61440 32016 61444
rect 32032 61500 32096 61504
rect 32032 61444 32036 61500
rect 32036 61444 32092 61500
rect 32092 61444 32096 61500
rect 32032 61440 32096 61444
rect 32112 61500 32176 61504
rect 32112 61444 32116 61500
rect 32116 61444 32172 61500
rect 32172 61444 32176 61500
rect 32112 61440 32176 61444
rect 32192 61500 32256 61504
rect 32192 61444 32196 61500
rect 32196 61444 32252 61500
rect 32252 61444 32256 61500
rect 32192 61440 32256 61444
rect 36952 61500 37016 61504
rect 36952 61444 36956 61500
rect 36956 61444 37012 61500
rect 37012 61444 37016 61500
rect 36952 61440 37016 61444
rect 37032 61500 37096 61504
rect 37032 61444 37036 61500
rect 37036 61444 37092 61500
rect 37092 61444 37096 61500
rect 37032 61440 37096 61444
rect 37112 61500 37176 61504
rect 37112 61444 37116 61500
rect 37116 61444 37172 61500
rect 37172 61444 37176 61500
rect 37112 61440 37176 61444
rect 37192 61500 37256 61504
rect 37192 61444 37196 61500
rect 37196 61444 37252 61500
rect 37252 61444 37256 61500
rect 37192 61440 37256 61444
rect 2612 60956 2676 60960
rect 2612 60900 2616 60956
rect 2616 60900 2672 60956
rect 2672 60900 2676 60956
rect 2612 60896 2676 60900
rect 2692 60956 2756 60960
rect 2692 60900 2696 60956
rect 2696 60900 2752 60956
rect 2752 60900 2756 60956
rect 2692 60896 2756 60900
rect 2772 60956 2836 60960
rect 2772 60900 2776 60956
rect 2776 60900 2832 60956
rect 2832 60900 2836 60956
rect 2772 60896 2836 60900
rect 2852 60956 2916 60960
rect 2852 60900 2856 60956
rect 2856 60900 2912 60956
rect 2912 60900 2916 60956
rect 2852 60896 2916 60900
rect 7612 60956 7676 60960
rect 7612 60900 7616 60956
rect 7616 60900 7672 60956
rect 7672 60900 7676 60956
rect 7612 60896 7676 60900
rect 7692 60956 7756 60960
rect 7692 60900 7696 60956
rect 7696 60900 7752 60956
rect 7752 60900 7756 60956
rect 7692 60896 7756 60900
rect 7772 60956 7836 60960
rect 7772 60900 7776 60956
rect 7776 60900 7832 60956
rect 7832 60900 7836 60956
rect 7772 60896 7836 60900
rect 7852 60956 7916 60960
rect 7852 60900 7856 60956
rect 7856 60900 7912 60956
rect 7912 60900 7916 60956
rect 7852 60896 7916 60900
rect 12612 60956 12676 60960
rect 12612 60900 12616 60956
rect 12616 60900 12672 60956
rect 12672 60900 12676 60956
rect 12612 60896 12676 60900
rect 12692 60956 12756 60960
rect 12692 60900 12696 60956
rect 12696 60900 12752 60956
rect 12752 60900 12756 60956
rect 12692 60896 12756 60900
rect 12772 60956 12836 60960
rect 12772 60900 12776 60956
rect 12776 60900 12832 60956
rect 12832 60900 12836 60956
rect 12772 60896 12836 60900
rect 12852 60956 12916 60960
rect 12852 60900 12856 60956
rect 12856 60900 12912 60956
rect 12912 60900 12916 60956
rect 12852 60896 12916 60900
rect 17612 60956 17676 60960
rect 17612 60900 17616 60956
rect 17616 60900 17672 60956
rect 17672 60900 17676 60956
rect 17612 60896 17676 60900
rect 17692 60956 17756 60960
rect 17692 60900 17696 60956
rect 17696 60900 17752 60956
rect 17752 60900 17756 60956
rect 17692 60896 17756 60900
rect 17772 60956 17836 60960
rect 17772 60900 17776 60956
rect 17776 60900 17832 60956
rect 17832 60900 17836 60956
rect 17772 60896 17836 60900
rect 17852 60956 17916 60960
rect 17852 60900 17856 60956
rect 17856 60900 17912 60956
rect 17912 60900 17916 60956
rect 17852 60896 17916 60900
rect 22612 60956 22676 60960
rect 22612 60900 22616 60956
rect 22616 60900 22672 60956
rect 22672 60900 22676 60956
rect 22612 60896 22676 60900
rect 22692 60956 22756 60960
rect 22692 60900 22696 60956
rect 22696 60900 22752 60956
rect 22752 60900 22756 60956
rect 22692 60896 22756 60900
rect 22772 60956 22836 60960
rect 22772 60900 22776 60956
rect 22776 60900 22832 60956
rect 22832 60900 22836 60956
rect 22772 60896 22836 60900
rect 22852 60956 22916 60960
rect 22852 60900 22856 60956
rect 22856 60900 22912 60956
rect 22912 60900 22916 60956
rect 22852 60896 22916 60900
rect 27612 60956 27676 60960
rect 27612 60900 27616 60956
rect 27616 60900 27672 60956
rect 27672 60900 27676 60956
rect 27612 60896 27676 60900
rect 27692 60956 27756 60960
rect 27692 60900 27696 60956
rect 27696 60900 27752 60956
rect 27752 60900 27756 60956
rect 27692 60896 27756 60900
rect 27772 60956 27836 60960
rect 27772 60900 27776 60956
rect 27776 60900 27832 60956
rect 27832 60900 27836 60956
rect 27772 60896 27836 60900
rect 27852 60956 27916 60960
rect 27852 60900 27856 60956
rect 27856 60900 27912 60956
rect 27912 60900 27916 60956
rect 27852 60896 27916 60900
rect 32612 60956 32676 60960
rect 32612 60900 32616 60956
rect 32616 60900 32672 60956
rect 32672 60900 32676 60956
rect 32612 60896 32676 60900
rect 32692 60956 32756 60960
rect 32692 60900 32696 60956
rect 32696 60900 32752 60956
rect 32752 60900 32756 60956
rect 32692 60896 32756 60900
rect 32772 60956 32836 60960
rect 32772 60900 32776 60956
rect 32776 60900 32832 60956
rect 32832 60900 32836 60956
rect 32772 60896 32836 60900
rect 32852 60956 32916 60960
rect 32852 60900 32856 60956
rect 32856 60900 32912 60956
rect 32912 60900 32916 60956
rect 32852 60896 32916 60900
rect 37612 60956 37676 60960
rect 37612 60900 37616 60956
rect 37616 60900 37672 60956
rect 37672 60900 37676 60956
rect 37612 60896 37676 60900
rect 37692 60956 37756 60960
rect 37692 60900 37696 60956
rect 37696 60900 37752 60956
rect 37752 60900 37756 60956
rect 37692 60896 37756 60900
rect 37772 60956 37836 60960
rect 37772 60900 37776 60956
rect 37776 60900 37832 60956
rect 37832 60900 37836 60956
rect 37772 60896 37836 60900
rect 37852 60956 37916 60960
rect 37852 60900 37856 60956
rect 37856 60900 37912 60956
rect 37912 60900 37916 60956
rect 37852 60896 37916 60900
rect 1952 60412 2016 60416
rect 1952 60356 1956 60412
rect 1956 60356 2012 60412
rect 2012 60356 2016 60412
rect 1952 60352 2016 60356
rect 2032 60412 2096 60416
rect 2032 60356 2036 60412
rect 2036 60356 2092 60412
rect 2092 60356 2096 60412
rect 2032 60352 2096 60356
rect 2112 60412 2176 60416
rect 2112 60356 2116 60412
rect 2116 60356 2172 60412
rect 2172 60356 2176 60412
rect 2112 60352 2176 60356
rect 2192 60412 2256 60416
rect 2192 60356 2196 60412
rect 2196 60356 2252 60412
rect 2252 60356 2256 60412
rect 2192 60352 2256 60356
rect 6952 60412 7016 60416
rect 6952 60356 6956 60412
rect 6956 60356 7012 60412
rect 7012 60356 7016 60412
rect 6952 60352 7016 60356
rect 7032 60412 7096 60416
rect 7032 60356 7036 60412
rect 7036 60356 7092 60412
rect 7092 60356 7096 60412
rect 7032 60352 7096 60356
rect 7112 60412 7176 60416
rect 7112 60356 7116 60412
rect 7116 60356 7172 60412
rect 7172 60356 7176 60412
rect 7112 60352 7176 60356
rect 7192 60412 7256 60416
rect 7192 60356 7196 60412
rect 7196 60356 7252 60412
rect 7252 60356 7256 60412
rect 7192 60352 7256 60356
rect 11952 60412 12016 60416
rect 11952 60356 11956 60412
rect 11956 60356 12012 60412
rect 12012 60356 12016 60412
rect 11952 60352 12016 60356
rect 12032 60412 12096 60416
rect 12032 60356 12036 60412
rect 12036 60356 12092 60412
rect 12092 60356 12096 60412
rect 12032 60352 12096 60356
rect 12112 60412 12176 60416
rect 12112 60356 12116 60412
rect 12116 60356 12172 60412
rect 12172 60356 12176 60412
rect 12112 60352 12176 60356
rect 12192 60412 12256 60416
rect 12192 60356 12196 60412
rect 12196 60356 12252 60412
rect 12252 60356 12256 60412
rect 12192 60352 12256 60356
rect 16952 60412 17016 60416
rect 16952 60356 16956 60412
rect 16956 60356 17012 60412
rect 17012 60356 17016 60412
rect 16952 60352 17016 60356
rect 17032 60412 17096 60416
rect 17032 60356 17036 60412
rect 17036 60356 17092 60412
rect 17092 60356 17096 60412
rect 17032 60352 17096 60356
rect 17112 60412 17176 60416
rect 17112 60356 17116 60412
rect 17116 60356 17172 60412
rect 17172 60356 17176 60412
rect 17112 60352 17176 60356
rect 17192 60412 17256 60416
rect 17192 60356 17196 60412
rect 17196 60356 17252 60412
rect 17252 60356 17256 60412
rect 17192 60352 17256 60356
rect 21952 60412 22016 60416
rect 21952 60356 21956 60412
rect 21956 60356 22012 60412
rect 22012 60356 22016 60412
rect 21952 60352 22016 60356
rect 22032 60412 22096 60416
rect 22032 60356 22036 60412
rect 22036 60356 22092 60412
rect 22092 60356 22096 60412
rect 22032 60352 22096 60356
rect 22112 60412 22176 60416
rect 22112 60356 22116 60412
rect 22116 60356 22172 60412
rect 22172 60356 22176 60412
rect 22112 60352 22176 60356
rect 22192 60412 22256 60416
rect 22192 60356 22196 60412
rect 22196 60356 22252 60412
rect 22252 60356 22256 60412
rect 22192 60352 22256 60356
rect 26952 60412 27016 60416
rect 26952 60356 26956 60412
rect 26956 60356 27012 60412
rect 27012 60356 27016 60412
rect 26952 60352 27016 60356
rect 27032 60412 27096 60416
rect 27032 60356 27036 60412
rect 27036 60356 27092 60412
rect 27092 60356 27096 60412
rect 27032 60352 27096 60356
rect 27112 60412 27176 60416
rect 27112 60356 27116 60412
rect 27116 60356 27172 60412
rect 27172 60356 27176 60412
rect 27112 60352 27176 60356
rect 27192 60412 27256 60416
rect 27192 60356 27196 60412
rect 27196 60356 27252 60412
rect 27252 60356 27256 60412
rect 27192 60352 27256 60356
rect 31952 60412 32016 60416
rect 31952 60356 31956 60412
rect 31956 60356 32012 60412
rect 32012 60356 32016 60412
rect 31952 60352 32016 60356
rect 32032 60412 32096 60416
rect 32032 60356 32036 60412
rect 32036 60356 32092 60412
rect 32092 60356 32096 60412
rect 32032 60352 32096 60356
rect 32112 60412 32176 60416
rect 32112 60356 32116 60412
rect 32116 60356 32172 60412
rect 32172 60356 32176 60412
rect 32112 60352 32176 60356
rect 32192 60412 32256 60416
rect 32192 60356 32196 60412
rect 32196 60356 32252 60412
rect 32252 60356 32256 60412
rect 32192 60352 32256 60356
rect 36952 60412 37016 60416
rect 36952 60356 36956 60412
rect 36956 60356 37012 60412
rect 37012 60356 37016 60412
rect 36952 60352 37016 60356
rect 37032 60412 37096 60416
rect 37032 60356 37036 60412
rect 37036 60356 37092 60412
rect 37092 60356 37096 60412
rect 37032 60352 37096 60356
rect 37112 60412 37176 60416
rect 37112 60356 37116 60412
rect 37116 60356 37172 60412
rect 37172 60356 37176 60412
rect 37112 60352 37176 60356
rect 37192 60412 37256 60416
rect 37192 60356 37196 60412
rect 37196 60356 37252 60412
rect 37252 60356 37256 60412
rect 37192 60352 37256 60356
rect 2612 59868 2676 59872
rect 2612 59812 2616 59868
rect 2616 59812 2672 59868
rect 2672 59812 2676 59868
rect 2612 59808 2676 59812
rect 2692 59868 2756 59872
rect 2692 59812 2696 59868
rect 2696 59812 2752 59868
rect 2752 59812 2756 59868
rect 2692 59808 2756 59812
rect 2772 59868 2836 59872
rect 2772 59812 2776 59868
rect 2776 59812 2832 59868
rect 2832 59812 2836 59868
rect 2772 59808 2836 59812
rect 2852 59868 2916 59872
rect 2852 59812 2856 59868
rect 2856 59812 2912 59868
rect 2912 59812 2916 59868
rect 2852 59808 2916 59812
rect 7612 59868 7676 59872
rect 7612 59812 7616 59868
rect 7616 59812 7672 59868
rect 7672 59812 7676 59868
rect 7612 59808 7676 59812
rect 7692 59868 7756 59872
rect 7692 59812 7696 59868
rect 7696 59812 7752 59868
rect 7752 59812 7756 59868
rect 7692 59808 7756 59812
rect 7772 59868 7836 59872
rect 7772 59812 7776 59868
rect 7776 59812 7832 59868
rect 7832 59812 7836 59868
rect 7772 59808 7836 59812
rect 7852 59868 7916 59872
rect 7852 59812 7856 59868
rect 7856 59812 7912 59868
rect 7912 59812 7916 59868
rect 7852 59808 7916 59812
rect 12612 59868 12676 59872
rect 12612 59812 12616 59868
rect 12616 59812 12672 59868
rect 12672 59812 12676 59868
rect 12612 59808 12676 59812
rect 12692 59868 12756 59872
rect 12692 59812 12696 59868
rect 12696 59812 12752 59868
rect 12752 59812 12756 59868
rect 12692 59808 12756 59812
rect 12772 59868 12836 59872
rect 12772 59812 12776 59868
rect 12776 59812 12832 59868
rect 12832 59812 12836 59868
rect 12772 59808 12836 59812
rect 12852 59868 12916 59872
rect 12852 59812 12856 59868
rect 12856 59812 12912 59868
rect 12912 59812 12916 59868
rect 12852 59808 12916 59812
rect 17612 59868 17676 59872
rect 17612 59812 17616 59868
rect 17616 59812 17672 59868
rect 17672 59812 17676 59868
rect 17612 59808 17676 59812
rect 17692 59868 17756 59872
rect 17692 59812 17696 59868
rect 17696 59812 17752 59868
rect 17752 59812 17756 59868
rect 17692 59808 17756 59812
rect 17772 59868 17836 59872
rect 17772 59812 17776 59868
rect 17776 59812 17832 59868
rect 17832 59812 17836 59868
rect 17772 59808 17836 59812
rect 17852 59868 17916 59872
rect 17852 59812 17856 59868
rect 17856 59812 17912 59868
rect 17912 59812 17916 59868
rect 17852 59808 17916 59812
rect 22612 59868 22676 59872
rect 22612 59812 22616 59868
rect 22616 59812 22672 59868
rect 22672 59812 22676 59868
rect 22612 59808 22676 59812
rect 22692 59868 22756 59872
rect 22692 59812 22696 59868
rect 22696 59812 22752 59868
rect 22752 59812 22756 59868
rect 22692 59808 22756 59812
rect 22772 59868 22836 59872
rect 22772 59812 22776 59868
rect 22776 59812 22832 59868
rect 22832 59812 22836 59868
rect 22772 59808 22836 59812
rect 22852 59868 22916 59872
rect 22852 59812 22856 59868
rect 22856 59812 22912 59868
rect 22912 59812 22916 59868
rect 22852 59808 22916 59812
rect 27612 59868 27676 59872
rect 27612 59812 27616 59868
rect 27616 59812 27672 59868
rect 27672 59812 27676 59868
rect 27612 59808 27676 59812
rect 27692 59868 27756 59872
rect 27692 59812 27696 59868
rect 27696 59812 27752 59868
rect 27752 59812 27756 59868
rect 27692 59808 27756 59812
rect 27772 59868 27836 59872
rect 27772 59812 27776 59868
rect 27776 59812 27832 59868
rect 27832 59812 27836 59868
rect 27772 59808 27836 59812
rect 27852 59868 27916 59872
rect 27852 59812 27856 59868
rect 27856 59812 27912 59868
rect 27912 59812 27916 59868
rect 27852 59808 27916 59812
rect 32612 59868 32676 59872
rect 32612 59812 32616 59868
rect 32616 59812 32672 59868
rect 32672 59812 32676 59868
rect 32612 59808 32676 59812
rect 32692 59868 32756 59872
rect 32692 59812 32696 59868
rect 32696 59812 32752 59868
rect 32752 59812 32756 59868
rect 32692 59808 32756 59812
rect 32772 59868 32836 59872
rect 32772 59812 32776 59868
rect 32776 59812 32832 59868
rect 32832 59812 32836 59868
rect 32772 59808 32836 59812
rect 32852 59868 32916 59872
rect 32852 59812 32856 59868
rect 32856 59812 32912 59868
rect 32912 59812 32916 59868
rect 32852 59808 32916 59812
rect 37612 59868 37676 59872
rect 37612 59812 37616 59868
rect 37616 59812 37672 59868
rect 37672 59812 37676 59868
rect 37612 59808 37676 59812
rect 37692 59868 37756 59872
rect 37692 59812 37696 59868
rect 37696 59812 37752 59868
rect 37752 59812 37756 59868
rect 37692 59808 37756 59812
rect 37772 59868 37836 59872
rect 37772 59812 37776 59868
rect 37776 59812 37832 59868
rect 37832 59812 37836 59868
rect 37772 59808 37836 59812
rect 37852 59868 37916 59872
rect 37852 59812 37856 59868
rect 37856 59812 37912 59868
rect 37912 59812 37916 59868
rect 37852 59808 37916 59812
rect 24900 59468 24964 59532
rect 1952 59324 2016 59328
rect 1952 59268 1956 59324
rect 1956 59268 2012 59324
rect 2012 59268 2016 59324
rect 1952 59264 2016 59268
rect 2032 59324 2096 59328
rect 2032 59268 2036 59324
rect 2036 59268 2092 59324
rect 2092 59268 2096 59324
rect 2032 59264 2096 59268
rect 2112 59324 2176 59328
rect 2112 59268 2116 59324
rect 2116 59268 2172 59324
rect 2172 59268 2176 59324
rect 2112 59264 2176 59268
rect 2192 59324 2256 59328
rect 2192 59268 2196 59324
rect 2196 59268 2252 59324
rect 2252 59268 2256 59324
rect 2192 59264 2256 59268
rect 6952 59324 7016 59328
rect 6952 59268 6956 59324
rect 6956 59268 7012 59324
rect 7012 59268 7016 59324
rect 6952 59264 7016 59268
rect 7032 59324 7096 59328
rect 7032 59268 7036 59324
rect 7036 59268 7092 59324
rect 7092 59268 7096 59324
rect 7032 59264 7096 59268
rect 7112 59324 7176 59328
rect 7112 59268 7116 59324
rect 7116 59268 7172 59324
rect 7172 59268 7176 59324
rect 7112 59264 7176 59268
rect 7192 59324 7256 59328
rect 7192 59268 7196 59324
rect 7196 59268 7252 59324
rect 7252 59268 7256 59324
rect 7192 59264 7256 59268
rect 11952 59324 12016 59328
rect 11952 59268 11956 59324
rect 11956 59268 12012 59324
rect 12012 59268 12016 59324
rect 11952 59264 12016 59268
rect 12032 59324 12096 59328
rect 12032 59268 12036 59324
rect 12036 59268 12092 59324
rect 12092 59268 12096 59324
rect 12032 59264 12096 59268
rect 12112 59324 12176 59328
rect 12112 59268 12116 59324
rect 12116 59268 12172 59324
rect 12172 59268 12176 59324
rect 12112 59264 12176 59268
rect 12192 59324 12256 59328
rect 12192 59268 12196 59324
rect 12196 59268 12252 59324
rect 12252 59268 12256 59324
rect 12192 59264 12256 59268
rect 16952 59324 17016 59328
rect 16952 59268 16956 59324
rect 16956 59268 17012 59324
rect 17012 59268 17016 59324
rect 16952 59264 17016 59268
rect 17032 59324 17096 59328
rect 17032 59268 17036 59324
rect 17036 59268 17092 59324
rect 17092 59268 17096 59324
rect 17032 59264 17096 59268
rect 17112 59324 17176 59328
rect 17112 59268 17116 59324
rect 17116 59268 17172 59324
rect 17172 59268 17176 59324
rect 17112 59264 17176 59268
rect 17192 59324 17256 59328
rect 17192 59268 17196 59324
rect 17196 59268 17252 59324
rect 17252 59268 17256 59324
rect 17192 59264 17256 59268
rect 21952 59324 22016 59328
rect 21952 59268 21956 59324
rect 21956 59268 22012 59324
rect 22012 59268 22016 59324
rect 21952 59264 22016 59268
rect 22032 59324 22096 59328
rect 22032 59268 22036 59324
rect 22036 59268 22092 59324
rect 22092 59268 22096 59324
rect 22032 59264 22096 59268
rect 22112 59324 22176 59328
rect 22112 59268 22116 59324
rect 22116 59268 22172 59324
rect 22172 59268 22176 59324
rect 22112 59264 22176 59268
rect 22192 59324 22256 59328
rect 22192 59268 22196 59324
rect 22196 59268 22252 59324
rect 22252 59268 22256 59324
rect 22192 59264 22256 59268
rect 26952 59324 27016 59328
rect 26952 59268 26956 59324
rect 26956 59268 27012 59324
rect 27012 59268 27016 59324
rect 26952 59264 27016 59268
rect 27032 59324 27096 59328
rect 27032 59268 27036 59324
rect 27036 59268 27092 59324
rect 27092 59268 27096 59324
rect 27032 59264 27096 59268
rect 27112 59324 27176 59328
rect 27112 59268 27116 59324
rect 27116 59268 27172 59324
rect 27172 59268 27176 59324
rect 27112 59264 27176 59268
rect 27192 59324 27256 59328
rect 27192 59268 27196 59324
rect 27196 59268 27252 59324
rect 27252 59268 27256 59324
rect 27192 59264 27256 59268
rect 31952 59324 32016 59328
rect 31952 59268 31956 59324
rect 31956 59268 32012 59324
rect 32012 59268 32016 59324
rect 31952 59264 32016 59268
rect 32032 59324 32096 59328
rect 32032 59268 32036 59324
rect 32036 59268 32092 59324
rect 32092 59268 32096 59324
rect 32032 59264 32096 59268
rect 32112 59324 32176 59328
rect 32112 59268 32116 59324
rect 32116 59268 32172 59324
rect 32172 59268 32176 59324
rect 32112 59264 32176 59268
rect 32192 59324 32256 59328
rect 32192 59268 32196 59324
rect 32196 59268 32252 59324
rect 32252 59268 32256 59324
rect 32192 59264 32256 59268
rect 36952 59324 37016 59328
rect 36952 59268 36956 59324
rect 36956 59268 37012 59324
rect 37012 59268 37016 59324
rect 36952 59264 37016 59268
rect 37032 59324 37096 59328
rect 37032 59268 37036 59324
rect 37036 59268 37092 59324
rect 37092 59268 37096 59324
rect 37032 59264 37096 59268
rect 37112 59324 37176 59328
rect 37112 59268 37116 59324
rect 37116 59268 37172 59324
rect 37172 59268 37176 59324
rect 37112 59264 37176 59268
rect 37192 59324 37256 59328
rect 37192 59268 37196 59324
rect 37196 59268 37252 59324
rect 37252 59268 37256 59324
rect 37192 59264 37256 59268
rect 2612 58780 2676 58784
rect 2612 58724 2616 58780
rect 2616 58724 2672 58780
rect 2672 58724 2676 58780
rect 2612 58720 2676 58724
rect 2692 58780 2756 58784
rect 2692 58724 2696 58780
rect 2696 58724 2752 58780
rect 2752 58724 2756 58780
rect 2692 58720 2756 58724
rect 2772 58780 2836 58784
rect 2772 58724 2776 58780
rect 2776 58724 2832 58780
rect 2832 58724 2836 58780
rect 2772 58720 2836 58724
rect 2852 58780 2916 58784
rect 2852 58724 2856 58780
rect 2856 58724 2912 58780
rect 2912 58724 2916 58780
rect 2852 58720 2916 58724
rect 7612 58780 7676 58784
rect 7612 58724 7616 58780
rect 7616 58724 7672 58780
rect 7672 58724 7676 58780
rect 7612 58720 7676 58724
rect 7692 58780 7756 58784
rect 7692 58724 7696 58780
rect 7696 58724 7752 58780
rect 7752 58724 7756 58780
rect 7692 58720 7756 58724
rect 7772 58780 7836 58784
rect 7772 58724 7776 58780
rect 7776 58724 7832 58780
rect 7832 58724 7836 58780
rect 7772 58720 7836 58724
rect 7852 58780 7916 58784
rect 7852 58724 7856 58780
rect 7856 58724 7912 58780
rect 7912 58724 7916 58780
rect 7852 58720 7916 58724
rect 12612 58780 12676 58784
rect 12612 58724 12616 58780
rect 12616 58724 12672 58780
rect 12672 58724 12676 58780
rect 12612 58720 12676 58724
rect 12692 58780 12756 58784
rect 12692 58724 12696 58780
rect 12696 58724 12752 58780
rect 12752 58724 12756 58780
rect 12692 58720 12756 58724
rect 12772 58780 12836 58784
rect 12772 58724 12776 58780
rect 12776 58724 12832 58780
rect 12832 58724 12836 58780
rect 12772 58720 12836 58724
rect 12852 58780 12916 58784
rect 12852 58724 12856 58780
rect 12856 58724 12912 58780
rect 12912 58724 12916 58780
rect 12852 58720 12916 58724
rect 17612 58780 17676 58784
rect 17612 58724 17616 58780
rect 17616 58724 17672 58780
rect 17672 58724 17676 58780
rect 17612 58720 17676 58724
rect 17692 58780 17756 58784
rect 17692 58724 17696 58780
rect 17696 58724 17752 58780
rect 17752 58724 17756 58780
rect 17692 58720 17756 58724
rect 17772 58780 17836 58784
rect 17772 58724 17776 58780
rect 17776 58724 17832 58780
rect 17832 58724 17836 58780
rect 17772 58720 17836 58724
rect 17852 58780 17916 58784
rect 17852 58724 17856 58780
rect 17856 58724 17912 58780
rect 17912 58724 17916 58780
rect 17852 58720 17916 58724
rect 22612 58780 22676 58784
rect 22612 58724 22616 58780
rect 22616 58724 22672 58780
rect 22672 58724 22676 58780
rect 22612 58720 22676 58724
rect 22692 58780 22756 58784
rect 22692 58724 22696 58780
rect 22696 58724 22752 58780
rect 22752 58724 22756 58780
rect 22692 58720 22756 58724
rect 22772 58780 22836 58784
rect 22772 58724 22776 58780
rect 22776 58724 22832 58780
rect 22832 58724 22836 58780
rect 22772 58720 22836 58724
rect 22852 58780 22916 58784
rect 22852 58724 22856 58780
rect 22856 58724 22912 58780
rect 22912 58724 22916 58780
rect 22852 58720 22916 58724
rect 27612 58780 27676 58784
rect 27612 58724 27616 58780
rect 27616 58724 27672 58780
rect 27672 58724 27676 58780
rect 27612 58720 27676 58724
rect 27692 58780 27756 58784
rect 27692 58724 27696 58780
rect 27696 58724 27752 58780
rect 27752 58724 27756 58780
rect 27692 58720 27756 58724
rect 27772 58780 27836 58784
rect 27772 58724 27776 58780
rect 27776 58724 27832 58780
rect 27832 58724 27836 58780
rect 27772 58720 27836 58724
rect 27852 58780 27916 58784
rect 27852 58724 27856 58780
rect 27856 58724 27912 58780
rect 27912 58724 27916 58780
rect 27852 58720 27916 58724
rect 32612 58780 32676 58784
rect 32612 58724 32616 58780
rect 32616 58724 32672 58780
rect 32672 58724 32676 58780
rect 32612 58720 32676 58724
rect 32692 58780 32756 58784
rect 32692 58724 32696 58780
rect 32696 58724 32752 58780
rect 32752 58724 32756 58780
rect 32692 58720 32756 58724
rect 32772 58780 32836 58784
rect 32772 58724 32776 58780
rect 32776 58724 32832 58780
rect 32832 58724 32836 58780
rect 32772 58720 32836 58724
rect 32852 58780 32916 58784
rect 32852 58724 32856 58780
rect 32856 58724 32912 58780
rect 32912 58724 32916 58780
rect 32852 58720 32916 58724
rect 37612 58780 37676 58784
rect 37612 58724 37616 58780
rect 37616 58724 37672 58780
rect 37672 58724 37676 58780
rect 37612 58720 37676 58724
rect 37692 58780 37756 58784
rect 37692 58724 37696 58780
rect 37696 58724 37752 58780
rect 37752 58724 37756 58780
rect 37692 58720 37756 58724
rect 37772 58780 37836 58784
rect 37772 58724 37776 58780
rect 37776 58724 37832 58780
rect 37832 58724 37836 58780
rect 37772 58720 37836 58724
rect 37852 58780 37916 58784
rect 37852 58724 37856 58780
rect 37856 58724 37912 58780
rect 37912 58724 37916 58780
rect 37852 58720 37916 58724
rect 1952 58236 2016 58240
rect 1952 58180 1956 58236
rect 1956 58180 2012 58236
rect 2012 58180 2016 58236
rect 1952 58176 2016 58180
rect 2032 58236 2096 58240
rect 2032 58180 2036 58236
rect 2036 58180 2092 58236
rect 2092 58180 2096 58236
rect 2032 58176 2096 58180
rect 2112 58236 2176 58240
rect 2112 58180 2116 58236
rect 2116 58180 2172 58236
rect 2172 58180 2176 58236
rect 2112 58176 2176 58180
rect 2192 58236 2256 58240
rect 2192 58180 2196 58236
rect 2196 58180 2252 58236
rect 2252 58180 2256 58236
rect 2192 58176 2256 58180
rect 6952 58236 7016 58240
rect 6952 58180 6956 58236
rect 6956 58180 7012 58236
rect 7012 58180 7016 58236
rect 6952 58176 7016 58180
rect 7032 58236 7096 58240
rect 7032 58180 7036 58236
rect 7036 58180 7092 58236
rect 7092 58180 7096 58236
rect 7032 58176 7096 58180
rect 7112 58236 7176 58240
rect 7112 58180 7116 58236
rect 7116 58180 7172 58236
rect 7172 58180 7176 58236
rect 7112 58176 7176 58180
rect 7192 58236 7256 58240
rect 7192 58180 7196 58236
rect 7196 58180 7252 58236
rect 7252 58180 7256 58236
rect 7192 58176 7256 58180
rect 11952 58236 12016 58240
rect 11952 58180 11956 58236
rect 11956 58180 12012 58236
rect 12012 58180 12016 58236
rect 11952 58176 12016 58180
rect 12032 58236 12096 58240
rect 12032 58180 12036 58236
rect 12036 58180 12092 58236
rect 12092 58180 12096 58236
rect 12032 58176 12096 58180
rect 12112 58236 12176 58240
rect 12112 58180 12116 58236
rect 12116 58180 12172 58236
rect 12172 58180 12176 58236
rect 12112 58176 12176 58180
rect 12192 58236 12256 58240
rect 12192 58180 12196 58236
rect 12196 58180 12252 58236
rect 12252 58180 12256 58236
rect 12192 58176 12256 58180
rect 16952 58236 17016 58240
rect 16952 58180 16956 58236
rect 16956 58180 17012 58236
rect 17012 58180 17016 58236
rect 16952 58176 17016 58180
rect 17032 58236 17096 58240
rect 17032 58180 17036 58236
rect 17036 58180 17092 58236
rect 17092 58180 17096 58236
rect 17032 58176 17096 58180
rect 17112 58236 17176 58240
rect 17112 58180 17116 58236
rect 17116 58180 17172 58236
rect 17172 58180 17176 58236
rect 17112 58176 17176 58180
rect 17192 58236 17256 58240
rect 17192 58180 17196 58236
rect 17196 58180 17252 58236
rect 17252 58180 17256 58236
rect 17192 58176 17256 58180
rect 21952 58236 22016 58240
rect 21952 58180 21956 58236
rect 21956 58180 22012 58236
rect 22012 58180 22016 58236
rect 21952 58176 22016 58180
rect 22032 58236 22096 58240
rect 22032 58180 22036 58236
rect 22036 58180 22092 58236
rect 22092 58180 22096 58236
rect 22032 58176 22096 58180
rect 22112 58236 22176 58240
rect 22112 58180 22116 58236
rect 22116 58180 22172 58236
rect 22172 58180 22176 58236
rect 22112 58176 22176 58180
rect 22192 58236 22256 58240
rect 22192 58180 22196 58236
rect 22196 58180 22252 58236
rect 22252 58180 22256 58236
rect 22192 58176 22256 58180
rect 26952 58236 27016 58240
rect 26952 58180 26956 58236
rect 26956 58180 27012 58236
rect 27012 58180 27016 58236
rect 26952 58176 27016 58180
rect 27032 58236 27096 58240
rect 27032 58180 27036 58236
rect 27036 58180 27092 58236
rect 27092 58180 27096 58236
rect 27032 58176 27096 58180
rect 27112 58236 27176 58240
rect 27112 58180 27116 58236
rect 27116 58180 27172 58236
rect 27172 58180 27176 58236
rect 27112 58176 27176 58180
rect 27192 58236 27256 58240
rect 27192 58180 27196 58236
rect 27196 58180 27252 58236
rect 27252 58180 27256 58236
rect 27192 58176 27256 58180
rect 31952 58236 32016 58240
rect 31952 58180 31956 58236
rect 31956 58180 32012 58236
rect 32012 58180 32016 58236
rect 31952 58176 32016 58180
rect 32032 58236 32096 58240
rect 32032 58180 32036 58236
rect 32036 58180 32092 58236
rect 32092 58180 32096 58236
rect 32032 58176 32096 58180
rect 32112 58236 32176 58240
rect 32112 58180 32116 58236
rect 32116 58180 32172 58236
rect 32172 58180 32176 58236
rect 32112 58176 32176 58180
rect 32192 58236 32256 58240
rect 32192 58180 32196 58236
rect 32196 58180 32252 58236
rect 32252 58180 32256 58236
rect 32192 58176 32256 58180
rect 36952 58236 37016 58240
rect 36952 58180 36956 58236
rect 36956 58180 37012 58236
rect 37012 58180 37016 58236
rect 36952 58176 37016 58180
rect 37032 58236 37096 58240
rect 37032 58180 37036 58236
rect 37036 58180 37092 58236
rect 37092 58180 37096 58236
rect 37032 58176 37096 58180
rect 37112 58236 37176 58240
rect 37112 58180 37116 58236
rect 37116 58180 37172 58236
rect 37172 58180 37176 58236
rect 37112 58176 37176 58180
rect 37192 58236 37256 58240
rect 37192 58180 37196 58236
rect 37196 58180 37252 58236
rect 37252 58180 37256 58236
rect 37192 58176 37256 58180
rect 2612 57692 2676 57696
rect 2612 57636 2616 57692
rect 2616 57636 2672 57692
rect 2672 57636 2676 57692
rect 2612 57632 2676 57636
rect 2692 57692 2756 57696
rect 2692 57636 2696 57692
rect 2696 57636 2752 57692
rect 2752 57636 2756 57692
rect 2692 57632 2756 57636
rect 2772 57692 2836 57696
rect 2772 57636 2776 57692
rect 2776 57636 2832 57692
rect 2832 57636 2836 57692
rect 2772 57632 2836 57636
rect 2852 57692 2916 57696
rect 2852 57636 2856 57692
rect 2856 57636 2912 57692
rect 2912 57636 2916 57692
rect 2852 57632 2916 57636
rect 7612 57692 7676 57696
rect 7612 57636 7616 57692
rect 7616 57636 7672 57692
rect 7672 57636 7676 57692
rect 7612 57632 7676 57636
rect 7692 57692 7756 57696
rect 7692 57636 7696 57692
rect 7696 57636 7752 57692
rect 7752 57636 7756 57692
rect 7692 57632 7756 57636
rect 7772 57692 7836 57696
rect 7772 57636 7776 57692
rect 7776 57636 7832 57692
rect 7832 57636 7836 57692
rect 7772 57632 7836 57636
rect 7852 57692 7916 57696
rect 7852 57636 7856 57692
rect 7856 57636 7912 57692
rect 7912 57636 7916 57692
rect 7852 57632 7916 57636
rect 12612 57692 12676 57696
rect 12612 57636 12616 57692
rect 12616 57636 12672 57692
rect 12672 57636 12676 57692
rect 12612 57632 12676 57636
rect 12692 57692 12756 57696
rect 12692 57636 12696 57692
rect 12696 57636 12752 57692
rect 12752 57636 12756 57692
rect 12692 57632 12756 57636
rect 12772 57692 12836 57696
rect 12772 57636 12776 57692
rect 12776 57636 12832 57692
rect 12832 57636 12836 57692
rect 12772 57632 12836 57636
rect 12852 57692 12916 57696
rect 12852 57636 12856 57692
rect 12856 57636 12912 57692
rect 12912 57636 12916 57692
rect 12852 57632 12916 57636
rect 17612 57692 17676 57696
rect 17612 57636 17616 57692
rect 17616 57636 17672 57692
rect 17672 57636 17676 57692
rect 17612 57632 17676 57636
rect 17692 57692 17756 57696
rect 17692 57636 17696 57692
rect 17696 57636 17752 57692
rect 17752 57636 17756 57692
rect 17692 57632 17756 57636
rect 17772 57692 17836 57696
rect 17772 57636 17776 57692
rect 17776 57636 17832 57692
rect 17832 57636 17836 57692
rect 17772 57632 17836 57636
rect 17852 57692 17916 57696
rect 17852 57636 17856 57692
rect 17856 57636 17912 57692
rect 17912 57636 17916 57692
rect 17852 57632 17916 57636
rect 22612 57692 22676 57696
rect 22612 57636 22616 57692
rect 22616 57636 22672 57692
rect 22672 57636 22676 57692
rect 22612 57632 22676 57636
rect 22692 57692 22756 57696
rect 22692 57636 22696 57692
rect 22696 57636 22752 57692
rect 22752 57636 22756 57692
rect 22692 57632 22756 57636
rect 22772 57692 22836 57696
rect 22772 57636 22776 57692
rect 22776 57636 22832 57692
rect 22832 57636 22836 57692
rect 22772 57632 22836 57636
rect 22852 57692 22916 57696
rect 22852 57636 22856 57692
rect 22856 57636 22912 57692
rect 22912 57636 22916 57692
rect 22852 57632 22916 57636
rect 27612 57692 27676 57696
rect 27612 57636 27616 57692
rect 27616 57636 27672 57692
rect 27672 57636 27676 57692
rect 27612 57632 27676 57636
rect 27692 57692 27756 57696
rect 27692 57636 27696 57692
rect 27696 57636 27752 57692
rect 27752 57636 27756 57692
rect 27692 57632 27756 57636
rect 27772 57692 27836 57696
rect 27772 57636 27776 57692
rect 27776 57636 27832 57692
rect 27832 57636 27836 57692
rect 27772 57632 27836 57636
rect 27852 57692 27916 57696
rect 27852 57636 27856 57692
rect 27856 57636 27912 57692
rect 27912 57636 27916 57692
rect 27852 57632 27916 57636
rect 32612 57692 32676 57696
rect 32612 57636 32616 57692
rect 32616 57636 32672 57692
rect 32672 57636 32676 57692
rect 32612 57632 32676 57636
rect 32692 57692 32756 57696
rect 32692 57636 32696 57692
rect 32696 57636 32752 57692
rect 32752 57636 32756 57692
rect 32692 57632 32756 57636
rect 32772 57692 32836 57696
rect 32772 57636 32776 57692
rect 32776 57636 32832 57692
rect 32832 57636 32836 57692
rect 32772 57632 32836 57636
rect 32852 57692 32916 57696
rect 32852 57636 32856 57692
rect 32856 57636 32912 57692
rect 32912 57636 32916 57692
rect 32852 57632 32916 57636
rect 37612 57692 37676 57696
rect 37612 57636 37616 57692
rect 37616 57636 37672 57692
rect 37672 57636 37676 57692
rect 37612 57632 37676 57636
rect 37692 57692 37756 57696
rect 37692 57636 37696 57692
rect 37696 57636 37752 57692
rect 37752 57636 37756 57692
rect 37692 57632 37756 57636
rect 37772 57692 37836 57696
rect 37772 57636 37776 57692
rect 37776 57636 37832 57692
rect 37832 57636 37836 57692
rect 37772 57632 37836 57636
rect 37852 57692 37916 57696
rect 37852 57636 37856 57692
rect 37856 57636 37912 57692
rect 37912 57636 37916 57692
rect 37852 57632 37916 57636
rect 1952 57148 2016 57152
rect 1952 57092 1956 57148
rect 1956 57092 2012 57148
rect 2012 57092 2016 57148
rect 1952 57088 2016 57092
rect 2032 57148 2096 57152
rect 2032 57092 2036 57148
rect 2036 57092 2092 57148
rect 2092 57092 2096 57148
rect 2032 57088 2096 57092
rect 2112 57148 2176 57152
rect 2112 57092 2116 57148
rect 2116 57092 2172 57148
rect 2172 57092 2176 57148
rect 2112 57088 2176 57092
rect 2192 57148 2256 57152
rect 2192 57092 2196 57148
rect 2196 57092 2252 57148
rect 2252 57092 2256 57148
rect 2192 57088 2256 57092
rect 6952 57148 7016 57152
rect 6952 57092 6956 57148
rect 6956 57092 7012 57148
rect 7012 57092 7016 57148
rect 6952 57088 7016 57092
rect 7032 57148 7096 57152
rect 7032 57092 7036 57148
rect 7036 57092 7092 57148
rect 7092 57092 7096 57148
rect 7032 57088 7096 57092
rect 7112 57148 7176 57152
rect 7112 57092 7116 57148
rect 7116 57092 7172 57148
rect 7172 57092 7176 57148
rect 7112 57088 7176 57092
rect 7192 57148 7256 57152
rect 7192 57092 7196 57148
rect 7196 57092 7252 57148
rect 7252 57092 7256 57148
rect 7192 57088 7256 57092
rect 11952 57148 12016 57152
rect 11952 57092 11956 57148
rect 11956 57092 12012 57148
rect 12012 57092 12016 57148
rect 11952 57088 12016 57092
rect 12032 57148 12096 57152
rect 12032 57092 12036 57148
rect 12036 57092 12092 57148
rect 12092 57092 12096 57148
rect 12032 57088 12096 57092
rect 12112 57148 12176 57152
rect 12112 57092 12116 57148
rect 12116 57092 12172 57148
rect 12172 57092 12176 57148
rect 12112 57088 12176 57092
rect 12192 57148 12256 57152
rect 12192 57092 12196 57148
rect 12196 57092 12252 57148
rect 12252 57092 12256 57148
rect 12192 57088 12256 57092
rect 16952 57148 17016 57152
rect 16952 57092 16956 57148
rect 16956 57092 17012 57148
rect 17012 57092 17016 57148
rect 16952 57088 17016 57092
rect 17032 57148 17096 57152
rect 17032 57092 17036 57148
rect 17036 57092 17092 57148
rect 17092 57092 17096 57148
rect 17032 57088 17096 57092
rect 17112 57148 17176 57152
rect 17112 57092 17116 57148
rect 17116 57092 17172 57148
rect 17172 57092 17176 57148
rect 17112 57088 17176 57092
rect 17192 57148 17256 57152
rect 17192 57092 17196 57148
rect 17196 57092 17252 57148
rect 17252 57092 17256 57148
rect 17192 57088 17256 57092
rect 21952 57148 22016 57152
rect 21952 57092 21956 57148
rect 21956 57092 22012 57148
rect 22012 57092 22016 57148
rect 21952 57088 22016 57092
rect 22032 57148 22096 57152
rect 22032 57092 22036 57148
rect 22036 57092 22092 57148
rect 22092 57092 22096 57148
rect 22032 57088 22096 57092
rect 22112 57148 22176 57152
rect 22112 57092 22116 57148
rect 22116 57092 22172 57148
rect 22172 57092 22176 57148
rect 22112 57088 22176 57092
rect 22192 57148 22256 57152
rect 22192 57092 22196 57148
rect 22196 57092 22252 57148
rect 22252 57092 22256 57148
rect 22192 57088 22256 57092
rect 26952 57148 27016 57152
rect 26952 57092 26956 57148
rect 26956 57092 27012 57148
rect 27012 57092 27016 57148
rect 26952 57088 27016 57092
rect 27032 57148 27096 57152
rect 27032 57092 27036 57148
rect 27036 57092 27092 57148
rect 27092 57092 27096 57148
rect 27032 57088 27096 57092
rect 27112 57148 27176 57152
rect 27112 57092 27116 57148
rect 27116 57092 27172 57148
rect 27172 57092 27176 57148
rect 27112 57088 27176 57092
rect 27192 57148 27256 57152
rect 27192 57092 27196 57148
rect 27196 57092 27252 57148
rect 27252 57092 27256 57148
rect 27192 57088 27256 57092
rect 31952 57148 32016 57152
rect 31952 57092 31956 57148
rect 31956 57092 32012 57148
rect 32012 57092 32016 57148
rect 31952 57088 32016 57092
rect 32032 57148 32096 57152
rect 32032 57092 32036 57148
rect 32036 57092 32092 57148
rect 32092 57092 32096 57148
rect 32032 57088 32096 57092
rect 32112 57148 32176 57152
rect 32112 57092 32116 57148
rect 32116 57092 32172 57148
rect 32172 57092 32176 57148
rect 32112 57088 32176 57092
rect 32192 57148 32256 57152
rect 32192 57092 32196 57148
rect 32196 57092 32252 57148
rect 32252 57092 32256 57148
rect 32192 57088 32256 57092
rect 36952 57148 37016 57152
rect 36952 57092 36956 57148
rect 36956 57092 37012 57148
rect 37012 57092 37016 57148
rect 36952 57088 37016 57092
rect 37032 57148 37096 57152
rect 37032 57092 37036 57148
rect 37036 57092 37092 57148
rect 37092 57092 37096 57148
rect 37032 57088 37096 57092
rect 37112 57148 37176 57152
rect 37112 57092 37116 57148
rect 37116 57092 37172 57148
rect 37172 57092 37176 57148
rect 37112 57088 37176 57092
rect 37192 57148 37256 57152
rect 37192 57092 37196 57148
rect 37196 57092 37252 57148
rect 37252 57092 37256 57148
rect 37192 57088 37256 57092
rect 18460 56748 18524 56812
rect 2612 56604 2676 56608
rect 2612 56548 2616 56604
rect 2616 56548 2672 56604
rect 2672 56548 2676 56604
rect 2612 56544 2676 56548
rect 2692 56604 2756 56608
rect 2692 56548 2696 56604
rect 2696 56548 2752 56604
rect 2752 56548 2756 56604
rect 2692 56544 2756 56548
rect 2772 56604 2836 56608
rect 2772 56548 2776 56604
rect 2776 56548 2832 56604
rect 2832 56548 2836 56604
rect 2772 56544 2836 56548
rect 2852 56604 2916 56608
rect 2852 56548 2856 56604
rect 2856 56548 2912 56604
rect 2912 56548 2916 56604
rect 2852 56544 2916 56548
rect 7612 56604 7676 56608
rect 7612 56548 7616 56604
rect 7616 56548 7672 56604
rect 7672 56548 7676 56604
rect 7612 56544 7676 56548
rect 7692 56604 7756 56608
rect 7692 56548 7696 56604
rect 7696 56548 7752 56604
rect 7752 56548 7756 56604
rect 7692 56544 7756 56548
rect 7772 56604 7836 56608
rect 7772 56548 7776 56604
rect 7776 56548 7832 56604
rect 7832 56548 7836 56604
rect 7772 56544 7836 56548
rect 7852 56604 7916 56608
rect 7852 56548 7856 56604
rect 7856 56548 7912 56604
rect 7912 56548 7916 56604
rect 7852 56544 7916 56548
rect 12612 56604 12676 56608
rect 12612 56548 12616 56604
rect 12616 56548 12672 56604
rect 12672 56548 12676 56604
rect 12612 56544 12676 56548
rect 12692 56604 12756 56608
rect 12692 56548 12696 56604
rect 12696 56548 12752 56604
rect 12752 56548 12756 56604
rect 12692 56544 12756 56548
rect 12772 56604 12836 56608
rect 12772 56548 12776 56604
rect 12776 56548 12832 56604
rect 12832 56548 12836 56604
rect 12772 56544 12836 56548
rect 12852 56604 12916 56608
rect 12852 56548 12856 56604
rect 12856 56548 12912 56604
rect 12912 56548 12916 56604
rect 12852 56544 12916 56548
rect 17612 56604 17676 56608
rect 17612 56548 17616 56604
rect 17616 56548 17672 56604
rect 17672 56548 17676 56604
rect 17612 56544 17676 56548
rect 17692 56604 17756 56608
rect 17692 56548 17696 56604
rect 17696 56548 17752 56604
rect 17752 56548 17756 56604
rect 17692 56544 17756 56548
rect 17772 56604 17836 56608
rect 17772 56548 17776 56604
rect 17776 56548 17832 56604
rect 17832 56548 17836 56604
rect 17772 56544 17836 56548
rect 17852 56604 17916 56608
rect 17852 56548 17856 56604
rect 17856 56548 17912 56604
rect 17912 56548 17916 56604
rect 17852 56544 17916 56548
rect 22612 56604 22676 56608
rect 22612 56548 22616 56604
rect 22616 56548 22672 56604
rect 22672 56548 22676 56604
rect 22612 56544 22676 56548
rect 22692 56604 22756 56608
rect 22692 56548 22696 56604
rect 22696 56548 22752 56604
rect 22752 56548 22756 56604
rect 22692 56544 22756 56548
rect 22772 56604 22836 56608
rect 22772 56548 22776 56604
rect 22776 56548 22832 56604
rect 22832 56548 22836 56604
rect 22772 56544 22836 56548
rect 22852 56604 22916 56608
rect 22852 56548 22856 56604
rect 22856 56548 22912 56604
rect 22912 56548 22916 56604
rect 22852 56544 22916 56548
rect 27612 56604 27676 56608
rect 27612 56548 27616 56604
rect 27616 56548 27672 56604
rect 27672 56548 27676 56604
rect 27612 56544 27676 56548
rect 27692 56604 27756 56608
rect 27692 56548 27696 56604
rect 27696 56548 27752 56604
rect 27752 56548 27756 56604
rect 27692 56544 27756 56548
rect 27772 56604 27836 56608
rect 27772 56548 27776 56604
rect 27776 56548 27832 56604
rect 27832 56548 27836 56604
rect 27772 56544 27836 56548
rect 27852 56604 27916 56608
rect 27852 56548 27856 56604
rect 27856 56548 27912 56604
rect 27912 56548 27916 56604
rect 27852 56544 27916 56548
rect 32612 56604 32676 56608
rect 32612 56548 32616 56604
rect 32616 56548 32672 56604
rect 32672 56548 32676 56604
rect 32612 56544 32676 56548
rect 32692 56604 32756 56608
rect 32692 56548 32696 56604
rect 32696 56548 32752 56604
rect 32752 56548 32756 56604
rect 32692 56544 32756 56548
rect 32772 56604 32836 56608
rect 32772 56548 32776 56604
rect 32776 56548 32832 56604
rect 32832 56548 32836 56604
rect 32772 56544 32836 56548
rect 32852 56604 32916 56608
rect 32852 56548 32856 56604
rect 32856 56548 32912 56604
rect 32912 56548 32916 56604
rect 32852 56544 32916 56548
rect 37612 56604 37676 56608
rect 37612 56548 37616 56604
rect 37616 56548 37672 56604
rect 37672 56548 37676 56604
rect 37612 56544 37676 56548
rect 37692 56604 37756 56608
rect 37692 56548 37696 56604
rect 37696 56548 37752 56604
rect 37752 56548 37756 56604
rect 37692 56544 37756 56548
rect 37772 56604 37836 56608
rect 37772 56548 37776 56604
rect 37776 56548 37832 56604
rect 37832 56548 37836 56604
rect 37772 56544 37836 56548
rect 37852 56604 37916 56608
rect 37852 56548 37856 56604
rect 37856 56548 37912 56604
rect 37912 56548 37916 56604
rect 37852 56544 37916 56548
rect 1952 56060 2016 56064
rect 1952 56004 1956 56060
rect 1956 56004 2012 56060
rect 2012 56004 2016 56060
rect 1952 56000 2016 56004
rect 2032 56060 2096 56064
rect 2032 56004 2036 56060
rect 2036 56004 2092 56060
rect 2092 56004 2096 56060
rect 2032 56000 2096 56004
rect 2112 56060 2176 56064
rect 2112 56004 2116 56060
rect 2116 56004 2172 56060
rect 2172 56004 2176 56060
rect 2112 56000 2176 56004
rect 2192 56060 2256 56064
rect 2192 56004 2196 56060
rect 2196 56004 2252 56060
rect 2252 56004 2256 56060
rect 2192 56000 2256 56004
rect 6952 56060 7016 56064
rect 6952 56004 6956 56060
rect 6956 56004 7012 56060
rect 7012 56004 7016 56060
rect 6952 56000 7016 56004
rect 7032 56060 7096 56064
rect 7032 56004 7036 56060
rect 7036 56004 7092 56060
rect 7092 56004 7096 56060
rect 7032 56000 7096 56004
rect 7112 56060 7176 56064
rect 7112 56004 7116 56060
rect 7116 56004 7172 56060
rect 7172 56004 7176 56060
rect 7112 56000 7176 56004
rect 7192 56060 7256 56064
rect 7192 56004 7196 56060
rect 7196 56004 7252 56060
rect 7252 56004 7256 56060
rect 7192 56000 7256 56004
rect 11952 56060 12016 56064
rect 11952 56004 11956 56060
rect 11956 56004 12012 56060
rect 12012 56004 12016 56060
rect 11952 56000 12016 56004
rect 12032 56060 12096 56064
rect 12032 56004 12036 56060
rect 12036 56004 12092 56060
rect 12092 56004 12096 56060
rect 12032 56000 12096 56004
rect 12112 56060 12176 56064
rect 12112 56004 12116 56060
rect 12116 56004 12172 56060
rect 12172 56004 12176 56060
rect 12112 56000 12176 56004
rect 12192 56060 12256 56064
rect 12192 56004 12196 56060
rect 12196 56004 12252 56060
rect 12252 56004 12256 56060
rect 12192 56000 12256 56004
rect 16952 56060 17016 56064
rect 16952 56004 16956 56060
rect 16956 56004 17012 56060
rect 17012 56004 17016 56060
rect 16952 56000 17016 56004
rect 17032 56060 17096 56064
rect 17032 56004 17036 56060
rect 17036 56004 17092 56060
rect 17092 56004 17096 56060
rect 17032 56000 17096 56004
rect 17112 56060 17176 56064
rect 17112 56004 17116 56060
rect 17116 56004 17172 56060
rect 17172 56004 17176 56060
rect 17112 56000 17176 56004
rect 17192 56060 17256 56064
rect 17192 56004 17196 56060
rect 17196 56004 17252 56060
rect 17252 56004 17256 56060
rect 17192 56000 17256 56004
rect 21952 56060 22016 56064
rect 21952 56004 21956 56060
rect 21956 56004 22012 56060
rect 22012 56004 22016 56060
rect 21952 56000 22016 56004
rect 22032 56060 22096 56064
rect 22032 56004 22036 56060
rect 22036 56004 22092 56060
rect 22092 56004 22096 56060
rect 22032 56000 22096 56004
rect 22112 56060 22176 56064
rect 22112 56004 22116 56060
rect 22116 56004 22172 56060
rect 22172 56004 22176 56060
rect 22112 56000 22176 56004
rect 22192 56060 22256 56064
rect 22192 56004 22196 56060
rect 22196 56004 22252 56060
rect 22252 56004 22256 56060
rect 22192 56000 22256 56004
rect 26952 56060 27016 56064
rect 26952 56004 26956 56060
rect 26956 56004 27012 56060
rect 27012 56004 27016 56060
rect 26952 56000 27016 56004
rect 27032 56060 27096 56064
rect 27032 56004 27036 56060
rect 27036 56004 27092 56060
rect 27092 56004 27096 56060
rect 27032 56000 27096 56004
rect 27112 56060 27176 56064
rect 27112 56004 27116 56060
rect 27116 56004 27172 56060
rect 27172 56004 27176 56060
rect 27112 56000 27176 56004
rect 27192 56060 27256 56064
rect 27192 56004 27196 56060
rect 27196 56004 27252 56060
rect 27252 56004 27256 56060
rect 27192 56000 27256 56004
rect 31952 56060 32016 56064
rect 31952 56004 31956 56060
rect 31956 56004 32012 56060
rect 32012 56004 32016 56060
rect 31952 56000 32016 56004
rect 32032 56060 32096 56064
rect 32032 56004 32036 56060
rect 32036 56004 32092 56060
rect 32092 56004 32096 56060
rect 32032 56000 32096 56004
rect 32112 56060 32176 56064
rect 32112 56004 32116 56060
rect 32116 56004 32172 56060
rect 32172 56004 32176 56060
rect 32112 56000 32176 56004
rect 32192 56060 32256 56064
rect 32192 56004 32196 56060
rect 32196 56004 32252 56060
rect 32252 56004 32256 56060
rect 32192 56000 32256 56004
rect 36952 56060 37016 56064
rect 36952 56004 36956 56060
rect 36956 56004 37012 56060
rect 37012 56004 37016 56060
rect 36952 56000 37016 56004
rect 37032 56060 37096 56064
rect 37032 56004 37036 56060
rect 37036 56004 37092 56060
rect 37092 56004 37096 56060
rect 37032 56000 37096 56004
rect 37112 56060 37176 56064
rect 37112 56004 37116 56060
rect 37116 56004 37172 56060
rect 37172 56004 37176 56060
rect 37112 56000 37176 56004
rect 37192 56060 37256 56064
rect 37192 56004 37196 56060
rect 37196 56004 37252 56060
rect 37252 56004 37256 56060
rect 37192 56000 37256 56004
rect 2612 55516 2676 55520
rect 2612 55460 2616 55516
rect 2616 55460 2672 55516
rect 2672 55460 2676 55516
rect 2612 55456 2676 55460
rect 2692 55516 2756 55520
rect 2692 55460 2696 55516
rect 2696 55460 2752 55516
rect 2752 55460 2756 55516
rect 2692 55456 2756 55460
rect 2772 55516 2836 55520
rect 2772 55460 2776 55516
rect 2776 55460 2832 55516
rect 2832 55460 2836 55516
rect 2772 55456 2836 55460
rect 2852 55516 2916 55520
rect 2852 55460 2856 55516
rect 2856 55460 2912 55516
rect 2912 55460 2916 55516
rect 2852 55456 2916 55460
rect 7612 55516 7676 55520
rect 7612 55460 7616 55516
rect 7616 55460 7672 55516
rect 7672 55460 7676 55516
rect 7612 55456 7676 55460
rect 7692 55516 7756 55520
rect 7692 55460 7696 55516
rect 7696 55460 7752 55516
rect 7752 55460 7756 55516
rect 7692 55456 7756 55460
rect 7772 55516 7836 55520
rect 7772 55460 7776 55516
rect 7776 55460 7832 55516
rect 7832 55460 7836 55516
rect 7772 55456 7836 55460
rect 7852 55516 7916 55520
rect 7852 55460 7856 55516
rect 7856 55460 7912 55516
rect 7912 55460 7916 55516
rect 7852 55456 7916 55460
rect 12612 55516 12676 55520
rect 12612 55460 12616 55516
rect 12616 55460 12672 55516
rect 12672 55460 12676 55516
rect 12612 55456 12676 55460
rect 12692 55516 12756 55520
rect 12692 55460 12696 55516
rect 12696 55460 12752 55516
rect 12752 55460 12756 55516
rect 12692 55456 12756 55460
rect 12772 55516 12836 55520
rect 12772 55460 12776 55516
rect 12776 55460 12832 55516
rect 12832 55460 12836 55516
rect 12772 55456 12836 55460
rect 12852 55516 12916 55520
rect 12852 55460 12856 55516
rect 12856 55460 12912 55516
rect 12912 55460 12916 55516
rect 12852 55456 12916 55460
rect 17612 55516 17676 55520
rect 17612 55460 17616 55516
rect 17616 55460 17672 55516
rect 17672 55460 17676 55516
rect 17612 55456 17676 55460
rect 17692 55516 17756 55520
rect 17692 55460 17696 55516
rect 17696 55460 17752 55516
rect 17752 55460 17756 55516
rect 17692 55456 17756 55460
rect 17772 55516 17836 55520
rect 17772 55460 17776 55516
rect 17776 55460 17832 55516
rect 17832 55460 17836 55516
rect 17772 55456 17836 55460
rect 17852 55516 17916 55520
rect 17852 55460 17856 55516
rect 17856 55460 17912 55516
rect 17912 55460 17916 55516
rect 17852 55456 17916 55460
rect 22612 55516 22676 55520
rect 22612 55460 22616 55516
rect 22616 55460 22672 55516
rect 22672 55460 22676 55516
rect 22612 55456 22676 55460
rect 22692 55516 22756 55520
rect 22692 55460 22696 55516
rect 22696 55460 22752 55516
rect 22752 55460 22756 55516
rect 22692 55456 22756 55460
rect 22772 55516 22836 55520
rect 22772 55460 22776 55516
rect 22776 55460 22832 55516
rect 22832 55460 22836 55516
rect 22772 55456 22836 55460
rect 22852 55516 22916 55520
rect 22852 55460 22856 55516
rect 22856 55460 22912 55516
rect 22912 55460 22916 55516
rect 22852 55456 22916 55460
rect 27612 55516 27676 55520
rect 27612 55460 27616 55516
rect 27616 55460 27672 55516
rect 27672 55460 27676 55516
rect 27612 55456 27676 55460
rect 27692 55516 27756 55520
rect 27692 55460 27696 55516
rect 27696 55460 27752 55516
rect 27752 55460 27756 55516
rect 27692 55456 27756 55460
rect 27772 55516 27836 55520
rect 27772 55460 27776 55516
rect 27776 55460 27832 55516
rect 27832 55460 27836 55516
rect 27772 55456 27836 55460
rect 27852 55516 27916 55520
rect 27852 55460 27856 55516
rect 27856 55460 27912 55516
rect 27912 55460 27916 55516
rect 27852 55456 27916 55460
rect 32612 55516 32676 55520
rect 32612 55460 32616 55516
rect 32616 55460 32672 55516
rect 32672 55460 32676 55516
rect 32612 55456 32676 55460
rect 32692 55516 32756 55520
rect 32692 55460 32696 55516
rect 32696 55460 32752 55516
rect 32752 55460 32756 55516
rect 32692 55456 32756 55460
rect 32772 55516 32836 55520
rect 32772 55460 32776 55516
rect 32776 55460 32832 55516
rect 32832 55460 32836 55516
rect 32772 55456 32836 55460
rect 32852 55516 32916 55520
rect 32852 55460 32856 55516
rect 32856 55460 32912 55516
rect 32912 55460 32916 55516
rect 32852 55456 32916 55460
rect 37612 55516 37676 55520
rect 37612 55460 37616 55516
rect 37616 55460 37672 55516
rect 37672 55460 37676 55516
rect 37612 55456 37676 55460
rect 37692 55516 37756 55520
rect 37692 55460 37696 55516
rect 37696 55460 37752 55516
rect 37752 55460 37756 55516
rect 37692 55456 37756 55460
rect 37772 55516 37836 55520
rect 37772 55460 37776 55516
rect 37776 55460 37832 55516
rect 37832 55460 37836 55516
rect 37772 55456 37836 55460
rect 37852 55516 37916 55520
rect 37852 55460 37856 55516
rect 37856 55460 37912 55516
rect 37912 55460 37916 55516
rect 37852 55456 37916 55460
rect 16436 55312 16500 55316
rect 16436 55256 16486 55312
rect 16486 55256 16500 55312
rect 16436 55252 16500 55256
rect 1952 54972 2016 54976
rect 1952 54916 1956 54972
rect 1956 54916 2012 54972
rect 2012 54916 2016 54972
rect 1952 54912 2016 54916
rect 2032 54972 2096 54976
rect 2032 54916 2036 54972
rect 2036 54916 2092 54972
rect 2092 54916 2096 54972
rect 2032 54912 2096 54916
rect 2112 54972 2176 54976
rect 2112 54916 2116 54972
rect 2116 54916 2172 54972
rect 2172 54916 2176 54972
rect 2112 54912 2176 54916
rect 2192 54972 2256 54976
rect 2192 54916 2196 54972
rect 2196 54916 2252 54972
rect 2252 54916 2256 54972
rect 2192 54912 2256 54916
rect 6952 54972 7016 54976
rect 6952 54916 6956 54972
rect 6956 54916 7012 54972
rect 7012 54916 7016 54972
rect 6952 54912 7016 54916
rect 7032 54972 7096 54976
rect 7032 54916 7036 54972
rect 7036 54916 7092 54972
rect 7092 54916 7096 54972
rect 7032 54912 7096 54916
rect 7112 54972 7176 54976
rect 7112 54916 7116 54972
rect 7116 54916 7172 54972
rect 7172 54916 7176 54972
rect 7112 54912 7176 54916
rect 7192 54972 7256 54976
rect 7192 54916 7196 54972
rect 7196 54916 7252 54972
rect 7252 54916 7256 54972
rect 7192 54912 7256 54916
rect 11952 54972 12016 54976
rect 11952 54916 11956 54972
rect 11956 54916 12012 54972
rect 12012 54916 12016 54972
rect 11952 54912 12016 54916
rect 12032 54972 12096 54976
rect 12032 54916 12036 54972
rect 12036 54916 12092 54972
rect 12092 54916 12096 54972
rect 12032 54912 12096 54916
rect 12112 54972 12176 54976
rect 12112 54916 12116 54972
rect 12116 54916 12172 54972
rect 12172 54916 12176 54972
rect 12112 54912 12176 54916
rect 12192 54972 12256 54976
rect 12192 54916 12196 54972
rect 12196 54916 12252 54972
rect 12252 54916 12256 54972
rect 12192 54912 12256 54916
rect 16952 54972 17016 54976
rect 16952 54916 16956 54972
rect 16956 54916 17012 54972
rect 17012 54916 17016 54972
rect 16952 54912 17016 54916
rect 17032 54972 17096 54976
rect 17032 54916 17036 54972
rect 17036 54916 17092 54972
rect 17092 54916 17096 54972
rect 17032 54912 17096 54916
rect 17112 54972 17176 54976
rect 17112 54916 17116 54972
rect 17116 54916 17172 54972
rect 17172 54916 17176 54972
rect 17112 54912 17176 54916
rect 17192 54972 17256 54976
rect 17192 54916 17196 54972
rect 17196 54916 17252 54972
rect 17252 54916 17256 54972
rect 17192 54912 17256 54916
rect 21952 54972 22016 54976
rect 21952 54916 21956 54972
rect 21956 54916 22012 54972
rect 22012 54916 22016 54972
rect 21952 54912 22016 54916
rect 22032 54972 22096 54976
rect 22032 54916 22036 54972
rect 22036 54916 22092 54972
rect 22092 54916 22096 54972
rect 22032 54912 22096 54916
rect 22112 54972 22176 54976
rect 22112 54916 22116 54972
rect 22116 54916 22172 54972
rect 22172 54916 22176 54972
rect 22112 54912 22176 54916
rect 22192 54972 22256 54976
rect 22192 54916 22196 54972
rect 22196 54916 22252 54972
rect 22252 54916 22256 54972
rect 22192 54912 22256 54916
rect 26952 54972 27016 54976
rect 26952 54916 26956 54972
rect 26956 54916 27012 54972
rect 27012 54916 27016 54972
rect 26952 54912 27016 54916
rect 27032 54972 27096 54976
rect 27032 54916 27036 54972
rect 27036 54916 27092 54972
rect 27092 54916 27096 54972
rect 27032 54912 27096 54916
rect 27112 54972 27176 54976
rect 27112 54916 27116 54972
rect 27116 54916 27172 54972
rect 27172 54916 27176 54972
rect 27112 54912 27176 54916
rect 27192 54972 27256 54976
rect 27192 54916 27196 54972
rect 27196 54916 27252 54972
rect 27252 54916 27256 54972
rect 27192 54912 27256 54916
rect 31952 54972 32016 54976
rect 31952 54916 31956 54972
rect 31956 54916 32012 54972
rect 32012 54916 32016 54972
rect 31952 54912 32016 54916
rect 32032 54972 32096 54976
rect 32032 54916 32036 54972
rect 32036 54916 32092 54972
rect 32092 54916 32096 54972
rect 32032 54912 32096 54916
rect 32112 54972 32176 54976
rect 32112 54916 32116 54972
rect 32116 54916 32172 54972
rect 32172 54916 32176 54972
rect 32112 54912 32176 54916
rect 32192 54972 32256 54976
rect 32192 54916 32196 54972
rect 32196 54916 32252 54972
rect 32252 54916 32256 54972
rect 32192 54912 32256 54916
rect 36952 54972 37016 54976
rect 36952 54916 36956 54972
rect 36956 54916 37012 54972
rect 37012 54916 37016 54972
rect 36952 54912 37016 54916
rect 37032 54972 37096 54976
rect 37032 54916 37036 54972
rect 37036 54916 37092 54972
rect 37092 54916 37096 54972
rect 37032 54912 37096 54916
rect 37112 54972 37176 54976
rect 37112 54916 37116 54972
rect 37116 54916 37172 54972
rect 37172 54916 37176 54972
rect 37112 54912 37176 54916
rect 37192 54972 37256 54976
rect 37192 54916 37196 54972
rect 37196 54916 37252 54972
rect 37252 54916 37256 54972
rect 37192 54912 37256 54916
rect 2612 54428 2676 54432
rect 2612 54372 2616 54428
rect 2616 54372 2672 54428
rect 2672 54372 2676 54428
rect 2612 54368 2676 54372
rect 2692 54428 2756 54432
rect 2692 54372 2696 54428
rect 2696 54372 2752 54428
rect 2752 54372 2756 54428
rect 2692 54368 2756 54372
rect 2772 54428 2836 54432
rect 2772 54372 2776 54428
rect 2776 54372 2832 54428
rect 2832 54372 2836 54428
rect 2772 54368 2836 54372
rect 2852 54428 2916 54432
rect 2852 54372 2856 54428
rect 2856 54372 2912 54428
rect 2912 54372 2916 54428
rect 2852 54368 2916 54372
rect 7612 54428 7676 54432
rect 7612 54372 7616 54428
rect 7616 54372 7672 54428
rect 7672 54372 7676 54428
rect 7612 54368 7676 54372
rect 7692 54428 7756 54432
rect 7692 54372 7696 54428
rect 7696 54372 7752 54428
rect 7752 54372 7756 54428
rect 7692 54368 7756 54372
rect 7772 54428 7836 54432
rect 7772 54372 7776 54428
rect 7776 54372 7832 54428
rect 7832 54372 7836 54428
rect 7772 54368 7836 54372
rect 7852 54428 7916 54432
rect 7852 54372 7856 54428
rect 7856 54372 7912 54428
rect 7912 54372 7916 54428
rect 7852 54368 7916 54372
rect 12612 54428 12676 54432
rect 12612 54372 12616 54428
rect 12616 54372 12672 54428
rect 12672 54372 12676 54428
rect 12612 54368 12676 54372
rect 12692 54428 12756 54432
rect 12692 54372 12696 54428
rect 12696 54372 12752 54428
rect 12752 54372 12756 54428
rect 12692 54368 12756 54372
rect 12772 54428 12836 54432
rect 12772 54372 12776 54428
rect 12776 54372 12832 54428
rect 12832 54372 12836 54428
rect 12772 54368 12836 54372
rect 12852 54428 12916 54432
rect 12852 54372 12856 54428
rect 12856 54372 12912 54428
rect 12912 54372 12916 54428
rect 12852 54368 12916 54372
rect 17612 54428 17676 54432
rect 17612 54372 17616 54428
rect 17616 54372 17672 54428
rect 17672 54372 17676 54428
rect 17612 54368 17676 54372
rect 17692 54428 17756 54432
rect 17692 54372 17696 54428
rect 17696 54372 17752 54428
rect 17752 54372 17756 54428
rect 17692 54368 17756 54372
rect 17772 54428 17836 54432
rect 17772 54372 17776 54428
rect 17776 54372 17832 54428
rect 17832 54372 17836 54428
rect 17772 54368 17836 54372
rect 17852 54428 17916 54432
rect 17852 54372 17856 54428
rect 17856 54372 17912 54428
rect 17912 54372 17916 54428
rect 17852 54368 17916 54372
rect 22612 54428 22676 54432
rect 22612 54372 22616 54428
rect 22616 54372 22672 54428
rect 22672 54372 22676 54428
rect 22612 54368 22676 54372
rect 22692 54428 22756 54432
rect 22692 54372 22696 54428
rect 22696 54372 22752 54428
rect 22752 54372 22756 54428
rect 22692 54368 22756 54372
rect 22772 54428 22836 54432
rect 22772 54372 22776 54428
rect 22776 54372 22832 54428
rect 22832 54372 22836 54428
rect 22772 54368 22836 54372
rect 22852 54428 22916 54432
rect 22852 54372 22856 54428
rect 22856 54372 22912 54428
rect 22912 54372 22916 54428
rect 22852 54368 22916 54372
rect 27612 54428 27676 54432
rect 27612 54372 27616 54428
rect 27616 54372 27672 54428
rect 27672 54372 27676 54428
rect 27612 54368 27676 54372
rect 27692 54428 27756 54432
rect 27692 54372 27696 54428
rect 27696 54372 27752 54428
rect 27752 54372 27756 54428
rect 27692 54368 27756 54372
rect 27772 54428 27836 54432
rect 27772 54372 27776 54428
rect 27776 54372 27832 54428
rect 27832 54372 27836 54428
rect 27772 54368 27836 54372
rect 27852 54428 27916 54432
rect 27852 54372 27856 54428
rect 27856 54372 27912 54428
rect 27912 54372 27916 54428
rect 27852 54368 27916 54372
rect 32612 54428 32676 54432
rect 32612 54372 32616 54428
rect 32616 54372 32672 54428
rect 32672 54372 32676 54428
rect 32612 54368 32676 54372
rect 32692 54428 32756 54432
rect 32692 54372 32696 54428
rect 32696 54372 32752 54428
rect 32752 54372 32756 54428
rect 32692 54368 32756 54372
rect 32772 54428 32836 54432
rect 32772 54372 32776 54428
rect 32776 54372 32832 54428
rect 32832 54372 32836 54428
rect 32772 54368 32836 54372
rect 32852 54428 32916 54432
rect 32852 54372 32856 54428
rect 32856 54372 32912 54428
rect 32912 54372 32916 54428
rect 32852 54368 32916 54372
rect 37612 54428 37676 54432
rect 37612 54372 37616 54428
rect 37616 54372 37672 54428
rect 37672 54372 37676 54428
rect 37612 54368 37676 54372
rect 37692 54428 37756 54432
rect 37692 54372 37696 54428
rect 37696 54372 37752 54428
rect 37752 54372 37756 54428
rect 37692 54368 37756 54372
rect 37772 54428 37836 54432
rect 37772 54372 37776 54428
rect 37776 54372 37832 54428
rect 37832 54372 37836 54428
rect 37772 54368 37836 54372
rect 37852 54428 37916 54432
rect 37852 54372 37856 54428
rect 37856 54372 37912 54428
rect 37912 54372 37916 54428
rect 37852 54368 37916 54372
rect 1952 53884 2016 53888
rect 1952 53828 1956 53884
rect 1956 53828 2012 53884
rect 2012 53828 2016 53884
rect 1952 53824 2016 53828
rect 2032 53884 2096 53888
rect 2032 53828 2036 53884
rect 2036 53828 2092 53884
rect 2092 53828 2096 53884
rect 2032 53824 2096 53828
rect 2112 53884 2176 53888
rect 2112 53828 2116 53884
rect 2116 53828 2172 53884
rect 2172 53828 2176 53884
rect 2112 53824 2176 53828
rect 2192 53884 2256 53888
rect 2192 53828 2196 53884
rect 2196 53828 2252 53884
rect 2252 53828 2256 53884
rect 2192 53824 2256 53828
rect 6952 53884 7016 53888
rect 6952 53828 6956 53884
rect 6956 53828 7012 53884
rect 7012 53828 7016 53884
rect 6952 53824 7016 53828
rect 7032 53884 7096 53888
rect 7032 53828 7036 53884
rect 7036 53828 7092 53884
rect 7092 53828 7096 53884
rect 7032 53824 7096 53828
rect 7112 53884 7176 53888
rect 7112 53828 7116 53884
rect 7116 53828 7172 53884
rect 7172 53828 7176 53884
rect 7112 53824 7176 53828
rect 7192 53884 7256 53888
rect 7192 53828 7196 53884
rect 7196 53828 7252 53884
rect 7252 53828 7256 53884
rect 7192 53824 7256 53828
rect 11952 53884 12016 53888
rect 11952 53828 11956 53884
rect 11956 53828 12012 53884
rect 12012 53828 12016 53884
rect 11952 53824 12016 53828
rect 12032 53884 12096 53888
rect 12032 53828 12036 53884
rect 12036 53828 12092 53884
rect 12092 53828 12096 53884
rect 12032 53824 12096 53828
rect 12112 53884 12176 53888
rect 12112 53828 12116 53884
rect 12116 53828 12172 53884
rect 12172 53828 12176 53884
rect 12112 53824 12176 53828
rect 12192 53884 12256 53888
rect 12192 53828 12196 53884
rect 12196 53828 12252 53884
rect 12252 53828 12256 53884
rect 12192 53824 12256 53828
rect 16952 53884 17016 53888
rect 16952 53828 16956 53884
rect 16956 53828 17012 53884
rect 17012 53828 17016 53884
rect 16952 53824 17016 53828
rect 17032 53884 17096 53888
rect 17032 53828 17036 53884
rect 17036 53828 17092 53884
rect 17092 53828 17096 53884
rect 17032 53824 17096 53828
rect 17112 53884 17176 53888
rect 17112 53828 17116 53884
rect 17116 53828 17172 53884
rect 17172 53828 17176 53884
rect 17112 53824 17176 53828
rect 17192 53884 17256 53888
rect 17192 53828 17196 53884
rect 17196 53828 17252 53884
rect 17252 53828 17256 53884
rect 17192 53824 17256 53828
rect 21952 53884 22016 53888
rect 21952 53828 21956 53884
rect 21956 53828 22012 53884
rect 22012 53828 22016 53884
rect 21952 53824 22016 53828
rect 22032 53884 22096 53888
rect 22032 53828 22036 53884
rect 22036 53828 22092 53884
rect 22092 53828 22096 53884
rect 22032 53824 22096 53828
rect 22112 53884 22176 53888
rect 22112 53828 22116 53884
rect 22116 53828 22172 53884
rect 22172 53828 22176 53884
rect 22112 53824 22176 53828
rect 22192 53884 22256 53888
rect 22192 53828 22196 53884
rect 22196 53828 22252 53884
rect 22252 53828 22256 53884
rect 22192 53824 22256 53828
rect 26952 53884 27016 53888
rect 26952 53828 26956 53884
rect 26956 53828 27012 53884
rect 27012 53828 27016 53884
rect 26952 53824 27016 53828
rect 27032 53884 27096 53888
rect 27032 53828 27036 53884
rect 27036 53828 27092 53884
rect 27092 53828 27096 53884
rect 27032 53824 27096 53828
rect 27112 53884 27176 53888
rect 27112 53828 27116 53884
rect 27116 53828 27172 53884
rect 27172 53828 27176 53884
rect 27112 53824 27176 53828
rect 27192 53884 27256 53888
rect 27192 53828 27196 53884
rect 27196 53828 27252 53884
rect 27252 53828 27256 53884
rect 27192 53824 27256 53828
rect 31952 53884 32016 53888
rect 31952 53828 31956 53884
rect 31956 53828 32012 53884
rect 32012 53828 32016 53884
rect 31952 53824 32016 53828
rect 32032 53884 32096 53888
rect 32032 53828 32036 53884
rect 32036 53828 32092 53884
rect 32092 53828 32096 53884
rect 32032 53824 32096 53828
rect 32112 53884 32176 53888
rect 32112 53828 32116 53884
rect 32116 53828 32172 53884
rect 32172 53828 32176 53884
rect 32112 53824 32176 53828
rect 32192 53884 32256 53888
rect 32192 53828 32196 53884
rect 32196 53828 32252 53884
rect 32252 53828 32256 53884
rect 32192 53824 32256 53828
rect 36952 53884 37016 53888
rect 36952 53828 36956 53884
rect 36956 53828 37012 53884
rect 37012 53828 37016 53884
rect 36952 53824 37016 53828
rect 37032 53884 37096 53888
rect 37032 53828 37036 53884
rect 37036 53828 37092 53884
rect 37092 53828 37096 53884
rect 37032 53824 37096 53828
rect 37112 53884 37176 53888
rect 37112 53828 37116 53884
rect 37116 53828 37172 53884
rect 37172 53828 37176 53884
rect 37112 53824 37176 53828
rect 37192 53884 37256 53888
rect 37192 53828 37196 53884
rect 37196 53828 37252 53884
rect 37252 53828 37256 53884
rect 37192 53824 37256 53828
rect 2612 53340 2676 53344
rect 2612 53284 2616 53340
rect 2616 53284 2672 53340
rect 2672 53284 2676 53340
rect 2612 53280 2676 53284
rect 2692 53340 2756 53344
rect 2692 53284 2696 53340
rect 2696 53284 2752 53340
rect 2752 53284 2756 53340
rect 2692 53280 2756 53284
rect 2772 53340 2836 53344
rect 2772 53284 2776 53340
rect 2776 53284 2832 53340
rect 2832 53284 2836 53340
rect 2772 53280 2836 53284
rect 2852 53340 2916 53344
rect 2852 53284 2856 53340
rect 2856 53284 2912 53340
rect 2912 53284 2916 53340
rect 2852 53280 2916 53284
rect 7612 53340 7676 53344
rect 7612 53284 7616 53340
rect 7616 53284 7672 53340
rect 7672 53284 7676 53340
rect 7612 53280 7676 53284
rect 7692 53340 7756 53344
rect 7692 53284 7696 53340
rect 7696 53284 7752 53340
rect 7752 53284 7756 53340
rect 7692 53280 7756 53284
rect 7772 53340 7836 53344
rect 7772 53284 7776 53340
rect 7776 53284 7832 53340
rect 7832 53284 7836 53340
rect 7772 53280 7836 53284
rect 7852 53340 7916 53344
rect 7852 53284 7856 53340
rect 7856 53284 7912 53340
rect 7912 53284 7916 53340
rect 7852 53280 7916 53284
rect 12612 53340 12676 53344
rect 12612 53284 12616 53340
rect 12616 53284 12672 53340
rect 12672 53284 12676 53340
rect 12612 53280 12676 53284
rect 12692 53340 12756 53344
rect 12692 53284 12696 53340
rect 12696 53284 12752 53340
rect 12752 53284 12756 53340
rect 12692 53280 12756 53284
rect 12772 53340 12836 53344
rect 12772 53284 12776 53340
rect 12776 53284 12832 53340
rect 12832 53284 12836 53340
rect 12772 53280 12836 53284
rect 12852 53340 12916 53344
rect 12852 53284 12856 53340
rect 12856 53284 12912 53340
rect 12912 53284 12916 53340
rect 12852 53280 12916 53284
rect 17612 53340 17676 53344
rect 17612 53284 17616 53340
rect 17616 53284 17672 53340
rect 17672 53284 17676 53340
rect 17612 53280 17676 53284
rect 17692 53340 17756 53344
rect 17692 53284 17696 53340
rect 17696 53284 17752 53340
rect 17752 53284 17756 53340
rect 17692 53280 17756 53284
rect 17772 53340 17836 53344
rect 17772 53284 17776 53340
rect 17776 53284 17832 53340
rect 17832 53284 17836 53340
rect 17772 53280 17836 53284
rect 17852 53340 17916 53344
rect 17852 53284 17856 53340
rect 17856 53284 17912 53340
rect 17912 53284 17916 53340
rect 17852 53280 17916 53284
rect 22612 53340 22676 53344
rect 22612 53284 22616 53340
rect 22616 53284 22672 53340
rect 22672 53284 22676 53340
rect 22612 53280 22676 53284
rect 22692 53340 22756 53344
rect 22692 53284 22696 53340
rect 22696 53284 22752 53340
rect 22752 53284 22756 53340
rect 22692 53280 22756 53284
rect 22772 53340 22836 53344
rect 22772 53284 22776 53340
rect 22776 53284 22832 53340
rect 22832 53284 22836 53340
rect 22772 53280 22836 53284
rect 22852 53340 22916 53344
rect 22852 53284 22856 53340
rect 22856 53284 22912 53340
rect 22912 53284 22916 53340
rect 22852 53280 22916 53284
rect 27612 53340 27676 53344
rect 27612 53284 27616 53340
rect 27616 53284 27672 53340
rect 27672 53284 27676 53340
rect 27612 53280 27676 53284
rect 27692 53340 27756 53344
rect 27692 53284 27696 53340
rect 27696 53284 27752 53340
rect 27752 53284 27756 53340
rect 27692 53280 27756 53284
rect 27772 53340 27836 53344
rect 27772 53284 27776 53340
rect 27776 53284 27832 53340
rect 27832 53284 27836 53340
rect 27772 53280 27836 53284
rect 27852 53340 27916 53344
rect 27852 53284 27856 53340
rect 27856 53284 27912 53340
rect 27912 53284 27916 53340
rect 27852 53280 27916 53284
rect 32612 53340 32676 53344
rect 32612 53284 32616 53340
rect 32616 53284 32672 53340
rect 32672 53284 32676 53340
rect 32612 53280 32676 53284
rect 32692 53340 32756 53344
rect 32692 53284 32696 53340
rect 32696 53284 32752 53340
rect 32752 53284 32756 53340
rect 32692 53280 32756 53284
rect 32772 53340 32836 53344
rect 32772 53284 32776 53340
rect 32776 53284 32832 53340
rect 32832 53284 32836 53340
rect 32772 53280 32836 53284
rect 32852 53340 32916 53344
rect 32852 53284 32856 53340
rect 32856 53284 32912 53340
rect 32912 53284 32916 53340
rect 32852 53280 32916 53284
rect 37612 53340 37676 53344
rect 37612 53284 37616 53340
rect 37616 53284 37672 53340
rect 37672 53284 37676 53340
rect 37612 53280 37676 53284
rect 37692 53340 37756 53344
rect 37692 53284 37696 53340
rect 37696 53284 37752 53340
rect 37752 53284 37756 53340
rect 37692 53280 37756 53284
rect 37772 53340 37836 53344
rect 37772 53284 37776 53340
rect 37776 53284 37832 53340
rect 37832 53284 37836 53340
rect 37772 53280 37836 53284
rect 37852 53340 37916 53344
rect 37852 53284 37856 53340
rect 37856 53284 37912 53340
rect 37912 53284 37916 53340
rect 37852 53280 37916 53284
rect 1952 52796 2016 52800
rect 1952 52740 1956 52796
rect 1956 52740 2012 52796
rect 2012 52740 2016 52796
rect 1952 52736 2016 52740
rect 2032 52796 2096 52800
rect 2032 52740 2036 52796
rect 2036 52740 2092 52796
rect 2092 52740 2096 52796
rect 2032 52736 2096 52740
rect 2112 52796 2176 52800
rect 2112 52740 2116 52796
rect 2116 52740 2172 52796
rect 2172 52740 2176 52796
rect 2112 52736 2176 52740
rect 2192 52796 2256 52800
rect 2192 52740 2196 52796
rect 2196 52740 2252 52796
rect 2252 52740 2256 52796
rect 2192 52736 2256 52740
rect 6952 52796 7016 52800
rect 6952 52740 6956 52796
rect 6956 52740 7012 52796
rect 7012 52740 7016 52796
rect 6952 52736 7016 52740
rect 7032 52796 7096 52800
rect 7032 52740 7036 52796
rect 7036 52740 7092 52796
rect 7092 52740 7096 52796
rect 7032 52736 7096 52740
rect 7112 52796 7176 52800
rect 7112 52740 7116 52796
rect 7116 52740 7172 52796
rect 7172 52740 7176 52796
rect 7112 52736 7176 52740
rect 7192 52796 7256 52800
rect 7192 52740 7196 52796
rect 7196 52740 7252 52796
rect 7252 52740 7256 52796
rect 7192 52736 7256 52740
rect 11952 52796 12016 52800
rect 11952 52740 11956 52796
rect 11956 52740 12012 52796
rect 12012 52740 12016 52796
rect 11952 52736 12016 52740
rect 12032 52796 12096 52800
rect 12032 52740 12036 52796
rect 12036 52740 12092 52796
rect 12092 52740 12096 52796
rect 12032 52736 12096 52740
rect 12112 52796 12176 52800
rect 12112 52740 12116 52796
rect 12116 52740 12172 52796
rect 12172 52740 12176 52796
rect 12112 52736 12176 52740
rect 12192 52796 12256 52800
rect 12192 52740 12196 52796
rect 12196 52740 12252 52796
rect 12252 52740 12256 52796
rect 12192 52736 12256 52740
rect 16952 52796 17016 52800
rect 16952 52740 16956 52796
rect 16956 52740 17012 52796
rect 17012 52740 17016 52796
rect 16952 52736 17016 52740
rect 17032 52796 17096 52800
rect 17032 52740 17036 52796
rect 17036 52740 17092 52796
rect 17092 52740 17096 52796
rect 17032 52736 17096 52740
rect 17112 52796 17176 52800
rect 17112 52740 17116 52796
rect 17116 52740 17172 52796
rect 17172 52740 17176 52796
rect 17112 52736 17176 52740
rect 17192 52796 17256 52800
rect 17192 52740 17196 52796
rect 17196 52740 17252 52796
rect 17252 52740 17256 52796
rect 17192 52736 17256 52740
rect 21952 52796 22016 52800
rect 21952 52740 21956 52796
rect 21956 52740 22012 52796
rect 22012 52740 22016 52796
rect 21952 52736 22016 52740
rect 22032 52796 22096 52800
rect 22032 52740 22036 52796
rect 22036 52740 22092 52796
rect 22092 52740 22096 52796
rect 22032 52736 22096 52740
rect 22112 52796 22176 52800
rect 22112 52740 22116 52796
rect 22116 52740 22172 52796
rect 22172 52740 22176 52796
rect 22112 52736 22176 52740
rect 22192 52796 22256 52800
rect 22192 52740 22196 52796
rect 22196 52740 22252 52796
rect 22252 52740 22256 52796
rect 22192 52736 22256 52740
rect 26952 52796 27016 52800
rect 26952 52740 26956 52796
rect 26956 52740 27012 52796
rect 27012 52740 27016 52796
rect 26952 52736 27016 52740
rect 27032 52796 27096 52800
rect 27032 52740 27036 52796
rect 27036 52740 27092 52796
rect 27092 52740 27096 52796
rect 27032 52736 27096 52740
rect 27112 52796 27176 52800
rect 27112 52740 27116 52796
rect 27116 52740 27172 52796
rect 27172 52740 27176 52796
rect 27112 52736 27176 52740
rect 27192 52796 27256 52800
rect 27192 52740 27196 52796
rect 27196 52740 27252 52796
rect 27252 52740 27256 52796
rect 27192 52736 27256 52740
rect 31952 52796 32016 52800
rect 31952 52740 31956 52796
rect 31956 52740 32012 52796
rect 32012 52740 32016 52796
rect 31952 52736 32016 52740
rect 32032 52796 32096 52800
rect 32032 52740 32036 52796
rect 32036 52740 32092 52796
rect 32092 52740 32096 52796
rect 32032 52736 32096 52740
rect 32112 52796 32176 52800
rect 32112 52740 32116 52796
rect 32116 52740 32172 52796
rect 32172 52740 32176 52796
rect 32112 52736 32176 52740
rect 32192 52796 32256 52800
rect 32192 52740 32196 52796
rect 32196 52740 32252 52796
rect 32252 52740 32256 52796
rect 32192 52736 32256 52740
rect 36952 52796 37016 52800
rect 36952 52740 36956 52796
rect 36956 52740 37012 52796
rect 37012 52740 37016 52796
rect 36952 52736 37016 52740
rect 37032 52796 37096 52800
rect 37032 52740 37036 52796
rect 37036 52740 37092 52796
rect 37092 52740 37096 52796
rect 37032 52736 37096 52740
rect 37112 52796 37176 52800
rect 37112 52740 37116 52796
rect 37116 52740 37172 52796
rect 37172 52740 37176 52796
rect 37112 52736 37176 52740
rect 37192 52796 37256 52800
rect 37192 52740 37196 52796
rect 37196 52740 37252 52796
rect 37252 52740 37256 52796
rect 37192 52736 37256 52740
rect 2612 52252 2676 52256
rect 2612 52196 2616 52252
rect 2616 52196 2672 52252
rect 2672 52196 2676 52252
rect 2612 52192 2676 52196
rect 2692 52252 2756 52256
rect 2692 52196 2696 52252
rect 2696 52196 2752 52252
rect 2752 52196 2756 52252
rect 2692 52192 2756 52196
rect 2772 52252 2836 52256
rect 2772 52196 2776 52252
rect 2776 52196 2832 52252
rect 2832 52196 2836 52252
rect 2772 52192 2836 52196
rect 2852 52252 2916 52256
rect 2852 52196 2856 52252
rect 2856 52196 2912 52252
rect 2912 52196 2916 52252
rect 2852 52192 2916 52196
rect 7612 52252 7676 52256
rect 7612 52196 7616 52252
rect 7616 52196 7672 52252
rect 7672 52196 7676 52252
rect 7612 52192 7676 52196
rect 7692 52252 7756 52256
rect 7692 52196 7696 52252
rect 7696 52196 7752 52252
rect 7752 52196 7756 52252
rect 7692 52192 7756 52196
rect 7772 52252 7836 52256
rect 7772 52196 7776 52252
rect 7776 52196 7832 52252
rect 7832 52196 7836 52252
rect 7772 52192 7836 52196
rect 7852 52252 7916 52256
rect 7852 52196 7856 52252
rect 7856 52196 7912 52252
rect 7912 52196 7916 52252
rect 7852 52192 7916 52196
rect 12612 52252 12676 52256
rect 12612 52196 12616 52252
rect 12616 52196 12672 52252
rect 12672 52196 12676 52252
rect 12612 52192 12676 52196
rect 12692 52252 12756 52256
rect 12692 52196 12696 52252
rect 12696 52196 12752 52252
rect 12752 52196 12756 52252
rect 12692 52192 12756 52196
rect 12772 52252 12836 52256
rect 12772 52196 12776 52252
rect 12776 52196 12832 52252
rect 12832 52196 12836 52252
rect 12772 52192 12836 52196
rect 12852 52252 12916 52256
rect 12852 52196 12856 52252
rect 12856 52196 12912 52252
rect 12912 52196 12916 52252
rect 12852 52192 12916 52196
rect 17612 52252 17676 52256
rect 17612 52196 17616 52252
rect 17616 52196 17672 52252
rect 17672 52196 17676 52252
rect 17612 52192 17676 52196
rect 17692 52252 17756 52256
rect 17692 52196 17696 52252
rect 17696 52196 17752 52252
rect 17752 52196 17756 52252
rect 17692 52192 17756 52196
rect 17772 52252 17836 52256
rect 17772 52196 17776 52252
rect 17776 52196 17832 52252
rect 17832 52196 17836 52252
rect 17772 52192 17836 52196
rect 17852 52252 17916 52256
rect 17852 52196 17856 52252
rect 17856 52196 17912 52252
rect 17912 52196 17916 52252
rect 17852 52192 17916 52196
rect 22612 52252 22676 52256
rect 22612 52196 22616 52252
rect 22616 52196 22672 52252
rect 22672 52196 22676 52252
rect 22612 52192 22676 52196
rect 22692 52252 22756 52256
rect 22692 52196 22696 52252
rect 22696 52196 22752 52252
rect 22752 52196 22756 52252
rect 22692 52192 22756 52196
rect 22772 52252 22836 52256
rect 22772 52196 22776 52252
rect 22776 52196 22832 52252
rect 22832 52196 22836 52252
rect 22772 52192 22836 52196
rect 22852 52252 22916 52256
rect 22852 52196 22856 52252
rect 22856 52196 22912 52252
rect 22912 52196 22916 52252
rect 22852 52192 22916 52196
rect 27612 52252 27676 52256
rect 27612 52196 27616 52252
rect 27616 52196 27672 52252
rect 27672 52196 27676 52252
rect 27612 52192 27676 52196
rect 27692 52252 27756 52256
rect 27692 52196 27696 52252
rect 27696 52196 27752 52252
rect 27752 52196 27756 52252
rect 27692 52192 27756 52196
rect 27772 52252 27836 52256
rect 27772 52196 27776 52252
rect 27776 52196 27832 52252
rect 27832 52196 27836 52252
rect 27772 52192 27836 52196
rect 27852 52252 27916 52256
rect 27852 52196 27856 52252
rect 27856 52196 27912 52252
rect 27912 52196 27916 52252
rect 27852 52192 27916 52196
rect 32612 52252 32676 52256
rect 32612 52196 32616 52252
rect 32616 52196 32672 52252
rect 32672 52196 32676 52252
rect 32612 52192 32676 52196
rect 32692 52252 32756 52256
rect 32692 52196 32696 52252
rect 32696 52196 32752 52252
rect 32752 52196 32756 52252
rect 32692 52192 32756 52196
rect 32772 52252 32836 52256
rect 32772 52196 32776 52252
rect 32776 52196 32832 52252
rect 32832 52196 32836 52252
rect 32772 52192 32836 52196
rect 32852 52252 32916 52256
rect 32852 52196 32856 52252
rect 32856 52196 32912 52252
rect 32912 52196 32916 52252
rect 32852 52192 32916 52196
rect 37612 52252 37676 52256
rect 37612 52196 37616 52252
rect 37616 52196 37672 52252
rect 37672 52196 37676 52252
rect 37612 52192 37676 52196
rect 37692 52252 37756 52256
rect 37692 52196 37696 52252
rect 37696 52196 37752 52252
rect 37752 52196 37756 52252
rect 37692 52192 37756 52196
rect 37772 52252 37836 52256
rect 37772 52196 37776 52252
rect 37776 52196 37832 52252
rect 37832 52196 37836 52252
rect 37772 52192 37836 52196
rect 37852 52252 37916 52256
rect 37852 52196 37856 52252
rect 37856 52196 37912 52252
rect 37912 52196 37916 52252
rect 37852 52192 37916 52196
rect 1952 51708 2016 51712
rect 1952 51652 1956 51708
rect 1956 51652 2012 51708
rect 2012 51652 2016 51708
rect 1952 51648 2016 51652
rect 2032 51708 2096 51712
rect 2032 51652 2036 51708
rect 2036 51652 2092 51708
rect 2092 51652 2096 51708
rect 2032 51648 2096 51652
rect 2112 51708 2176 51712
rect 2112 51652 2116 51708
rect 2116 51652 2172 51708
rect 2172 51652 2176 51708
rect 2112 51648 2176 51652
rect 2192 51708 2256 51712
rect 2192 51652 2196 51708
rect 2196 51652 2252 51708
rect 2252 51652 2256 51708
rect 2192 51648 2256 51652
rect 6952 51708 7016 51712
rect 6952 51652 6956 51708
rect 6956 51652 7012 51708
rect 7012 51652 7016 51708
rect 6952 51648 7016 51652
rect 7032 51708 7096 51712
rect 7032 51652 7036 51708
rect 7036 51652 7092 51708
rect 7092 51652 7096 51708
rect 7032 51648 7096 51652
rect 7112 51708 7176 51712
rect 7112 51652 7116 51708
rect 7116 51652 7172 51708
rect 7172 51652 7176 51708
rect 7112 51648 7176 51652
rect 7192 51708 7256 51712
rect 7192 51652 7196 51708
rect 7196 51652 7252 51708
rect 7252 51652 7256 51708
rect 7192 51648 7256 51652
rect 11952 51708 12016 51712
rect 11952 51652 11956 51708
rect 11956 51652 12012 51708
rect 12012 51652 12016 51708
rect 11952 51648 12016 51652
rect 12032 51708 12096 51712
rect 12032 51652 12036 51708
rect 12036 51652 12092 51708
rect 12092 51652 12096 51708
rect 12032 51648 12096 51652
rect 12112 51708 12176 51712
rect 12112 51652 12116 51708
rect 12116 51652 12172 51708
rect 12172 51652 12176 51708
rect 12112 51648 12176 51652
rect 12192 51708 12256 51712
rect 12192 51652 12196 51708
rect 12196 51652 12252 51708
rect 12252 51652 12256 51708
rect 12192 51648 12256 51652
rect 16952 51708 17016 51712
rect 16952 51652 16956 51708
rect 16956 51652 17012 51708
rect 17012 51652 17016 51708
rect 16952 51648 17016 51652
rect 17032 51708 17096 51712
rect 17032 51652 17036 51708
rect 17036 51652 17092 51708
rect 17092 51652 17096 51708
rect 17032 51648 17096 51652
rect 17112 51708 17176 51712
rect 17112 51652 17116 51708
rect 17116 51652 17172 51708
rect 17172 51652 17176 51708
rect 17112 51648 17176 51652
rect 17192 51708 17256 51712
rect 17192 51652 17196 51708
rect 17196 51652 17252 51708
rect 17252 51652 17256 51708
rect 17192 51648 17256 51652
rect 21952 51708 22016 51712
rect 21952 51652 21956 51708
rect 21956 51652 22012 51708
rect 22012 51652 22016 51708
rect 21952 51648 22016 51652
rect 22032 51708 22096 51712
rect 22032 51652 22036 51708
rect 22036 51652 22092 51708
rect 22092 51652 22096 51708
rect 22032 51648 22096 51652
rect 22112 51708 22176 51712
rect 22112 51652 22116 51708
rect 22116 51652 22172 51708
rect 22172 51652 22176 51708
rect 22112 51648 22176 51652
rect 22192 51708 22256 51712
rect 22192 51652 22196 51708
rect 22196 51652 22252 51708
rect 22252 51652 22256 51708
rect 22192 51648 22256 51652
rect 26952 51708 27016 51712
rect 26952 51652 26956 51708
rect 26956 51652 27012 51708
rect 27012 51652 27016 51708
rect 26952 51648 27016 51652
rect 27032 51708 27096 51712
rect 27032 51652 27036 51708
rect 27036 51652 27092 51708
rect 27092 51652 27096 51708
rect 27032 51648 27096 51652
rect 27112 51708 27176 51712
rect 27112 51652 27116 51708
rect 27116 51652 27172 51708
rect 27172 51652 27176 51708
rect 27112 51648 27176 51652
rect 27192 51708 27256 51712
rect 27192 51652 27196 51708
rect 27196 51652 27252 51708
rect 27252 51652 27256 51708
rect 27192 51648 27256 51652
rect 31952 51708 32016 51712
rect 31952 51652 31956 51708
rect 31956 51652 32012 51708
rect 32012 51652 32016 51708
rect 31952 51648 32016 51652
rect 32032 51708 32096 51712
rect 32032 51652 32036 51708
rect 32036 51652 32092 51708
rect 32092 51652 32096 51708
rect 32032 51648 32096 51652
rect 32112 51708 32176 51712
rect 32112 51652 32116 51708
rect 32116 51652 32172 51708
rect 32172 51652 32176 51708
rect 32112 51648 32176 51652
rect 32192 51708 32256 51712
rect 32192 51652 32196 51708
rect 32196 51652 32252 51708
rect 32252 51652 32256 51708
rect 32192 51648 32256 51652
rect 36952 51708 37016 51712
rect 36952 51652 36956 51708
rect 36956 51652 37012 51708
rect 37012 51652 37016 51708
rect 36952 51648 37016 51652
rect 37032 51708 37096 51712
rect 37032 51652 37036 51708
rect 37036 51652 37092 51708
rect 37092 51652 37096 51708
rect 37032 51648 37096 51652
rect 37112 51708 37176 51712
rect 37112 51652 37116 51708
rect 37116 51652 37172 51708
rect 37172 51652 37176 51708
rect 37112 51648 37176 51652
rect 37192 51708 37256 51712
rect 37192 51652 37196 51708
rect 37196 51652 37252 51708
rect 37252 51652 37256 51708
rect 37192 51648 37256 51652
rect 2612 51164 2676 51168
rect 2612 51108 2616 51164
rect 2616 51108 2672 51164
rect 2672 51108 2676 51164
rect 2612 51104 2676 51108
rect 2692 51164 2756 51168
rect 2692 51108 2696 51164
rect 2696 51108 2752 51164
rect 2752 51108 2756 51164
rect 2692 51104 2756 51108
rect 2772 51164 2836 51168
rect 2772 51108 2776 51164
rect 2776 51108 2832 51164
rect 2832 51108 2836 51164
rect 2772 51104 2836 51108
rect 2852 51164 2916 51168
rect 2852 51108 2856 51164
rect 2856 51108 2912 51164
rect 2912 51108 2916 51164
rect 2852 51104 2916 51108
rect 7612 51164 7676 51168
rect 7612 51108 7616 51164
rect 7616 51108 7672 51164
rect 7672 51108 7676 51164
rect 7612 51104 7676 51108
rect 7692 51164 7756 51168
rect 7692 51108 7696 51164
rect 7696 51108 7752 51164
rect 7752 51108 7756 51164
rect 7692 51104 7756 51108
rect 7772 51164 7836 51168
rect 7772 51108 7776 51164
rect 7776 51108 7832 51164
rect 7832 51108 7836 51164
rect 7772 51104 7836 51108
rect 7852 51164 7916 51168
rect 7852 51108 7856 51164
rect 7856 51108 7912 51164
rect 7912 51108 7916 51164
rect 7852 51104 7916 51108
rect 12612 51164 12676 51168
rect 12612 51108 12616 51164
rect 12616 51108 12672 51164
rect 12672 51108 12676 51164
rect 12612 51104 12676 51108
rect 12692 51164 12756 51168
rect 12692 51108 12696 51164
rect 12696 51108 12752 51164
rect 12752 51108 12756 51164
rect 12692 51104 12756 51108
rect 12772 51164 12836 51168
rect 12772 51108 12776 51164
rect 12776 51108 12832 51164
rect 12832 51108 12836 51164
rect 12772 51104 12836 51108
rect 12852 51164 12916 51168
rect 12852 51108 12856 51164
rect 12856 51108 12912 51164
rect 12912 51108 12916 51164
rect 12852 51104 12916 51108
rect 17612 51164 17676 51168
rect 17612 51108 17616 51164
rect 17616 51108 17672 51164
rect 17672 51108 17676 51164
rect 17612 51104 17676 51108
rect 17692 51164 17756 51168
rect 17692 51108 17696 51164
rect 17696 51108 17752 51164
rect 17752 51108 17756 51164
rect 17692 51104 17756 51108
rect 17772 51164 17836 51168
rect 17772 51108 17776 51164
rect 17776 51108 17832 51164
rect 17832 51108 17836 51164
rect 17772 51104 17836 51108
rect 17852 51164 17916 51168
rect 17852 51108 17856 51164
rect 17856 51108 17912 51164
rect 17912 51108 17916 51164
rect 17852 51104 17916 51108
rect 22612 51164 22676 51168
rect 22612 51108 22616 51164
rect 22616 51108 22672 51164
rect 22672 51108 22676 51164
rect 22612 51104 22676 51108
rect 22692 51164 22756 51168
rect 22692 51108 22696 51164
rect 22696 51108 22752 51164
rect 22752 51108 22756 51164
rect 22692 51104 22756 51108
rect 22772 51164 22836 51168
rect 22772 51108 22776 51164
rect 22776 51108 22832 51164
rect 22832 51108 22836 51164
rect 22772 51104 22836 51108
rect 22852 51164 22916 51168
rect 22852 51108 22856 51164
rect 22856 51108 22912 51164
rect 22912 51108 22916 51164
rect 22852 51104 22916 51108
rect 27612 51164 27676 51168
rect 27612 51108 27616 51164
rect 27616 51108 27672 51164
rect 27672 51108 27676 51164
rect 27612 51104 27676 51108
rect 27692 51164 27756 51168
rect 27692 51108 27696 51164
rect 27696 51108 27752 51164
rect 27752 51108 27756 51164
rect 27692 51104 27756 51108
rect 27772 51164 27836 51168
rect 27772 51108 27776 51164
rect 27776 51108 27832 51164
rect 27832 51108 27836 51164
rect 27772 51104 27836 51108
rect 27852 51164 27916 51168
rect 27852 51108 27856 51164
rect 27856 51108 27912 51164
rect 27912 51108 27916 51164
rect 27852 51104 27916 51108
rect 32612 51164 32676 51168
rect 32612 51108 32616 51164
rect 32616 51108 32672 51164
rect 32672 51108 32676 51164
rect 32612 51104 32676 51108
rect 32692 51164 32756 51168
rect 32692 51108 32696 51164
rect 32696 51108 32752 51164
rect 32752 51108 32756 51164
rect 32692 51104 32756 51108
rect 32772 51164 32836 51168
rect 32772 51108 32776 51164
rect 32776 51108 32832 51164
rect 32832 51108 32836 51164
rect 32772 51104 32836 51108
rect 32852 51164 32916 51168
rect 32852 51108 32856 51164
rect 32856 51108 32912 51164
rect 32912 51108 32916 51164
rect 32852 51104 32916 51108
rect 37612 51164 37676 51168
rect 37612 51108 37616 51164
rect 37616 51108 37672 51164
rect 37672 51108 37676 51164
rect 37612 51104 37676 51108
rect 37692 51164 37756 51168
rect 37692 51108 37696 51164
rect 37696 51108 37752 51164
rect 37752 51108 37756 51164
rect 37692 51104 37756 51108
rect 37772 51164 37836 51168
rect 37772 51108 37776 51164
rect 37776 51108 37832 51164
rect 37832 51108 37836 51164
rect 37772 51104 37836 51108
rect 37852 51164 37916 51168
rect 37852 51108 37856 51164
rect 37856 51108 37912 51164
rect 37912 51108 37916 51164
rect 37852 51104 37916 51108
rect 34836 51036 34900 51100
rect 1952 50620 2016 50624
rect 1952 50564 1956 50620
rect 1956 50564 2012 50620
rect 2012 50564 2016 50620
rect 1952 50560 2016 50564
rect 2032 50620 2096 50624
rect 2032 50564 2036 50620
rect 2036 50564 2092 50620
rect 2092 50564 2096 50620
rect 2032 50560 2096 50564
rect 2112 50620 2176 50624
rect 2112 50564 2116 50620
rect 2116 50564 2172 50620
rect 2172 50564 2176 50620
rect 2112 50560 2176 50564
rect 2192 50620 2256 50624
rect 2192 50564 2196 50620
rect 2196 50564 2252 50620
rect 2252 50564 2256 50620
rect 2192 50560 2256 50564
rect 6952 50620 7016 50624
rect 6952 50564 6956 50620
rect 6956 50564 7012 50620
rect 7012 50564 7016 50620
rect 6952 50560 7016 50564
rect 7032 50620 7096 50624
rect 7032 50564 7036 50620
rect 7036 50564 7092 50620
rect 7092 50564 7096 50620
rect 7032 50560 7096 50564
rect 7112 50620 7176 50624
rect 7112 50564 7116 50620
rect 7116 50564 7172 50620
rect 7172 50564 7176 50620
rect 7112 50560 7176 50564
rect 7192 50620 7256 50624
rect 7192 50564 7196 50620
rect 7196 50564 7252 50620
rect 7252 50564 7256 50620
rect 7192 50560 7256 50564
rect 11952 50620 12016 50624
rect 11952 50564 11956 50620
rect 11956 50564 12012 50620
rect 12012 50564 12016 50620
rect 11952 50560 12016 50564
rect 12032 50620 12096 50624
rect 12032 50564 12036 50620
rect 12036 50564 12092 50620
rect 12092 50564 12096 50620
rect 12032 50560 12096 50564
rect 12112 50620 12176 50624
rect 12112 50564 12116 50620
rect 12116 50564 12172 50620
rect 12172 50564 12176 50620
rect 12112 50560 12176 50564
rect 12192 50620 12256 50624
rect 12192 50564 12196 50620
rect 12196 50564 12252 50620
rect 12252 50564 12256 50620
rect 12192 50560 12256 50564
rect 16952 50620 17016 50624
rect 16952 50564 16956 50620
rect 16956 50564 17012 50620
rect 17012 50564 17016 50620
rect 16952 50560 17016 50564
rect 17032 50620 17096 50624
rect 17032 50564 17036 50620
rect 17036 50564 17092 50620
rect 17092 50564 17096 50620
rect 17032 50560 17096 50564
rect 17112 50620 17176 50624
rect 17112 50564 17116 50620
rect 17116 50564 17172 50620
rect 17172 50564 17176 50620
rect 17112 50560 17176 50564
rect 17192 50620 17256 50624
rect 17192 50564 17196 50620
rect 17196 50564 17252 50620
rect 17252 50564 17256 50620
rect 17192 50560 17256 50564
rect 21952 50620 22016 50624
rect 21952 50564 21956 50620
rect 21956 50564 22012 50620
rect 22012 50564 22016 50620
rect 21952 50560 22016 50564
rect 22032 50620 22096 50624
rect 22032 50564 22036 50620
rect 22036 50564 22092 50620
rect 22092 50564 22096 50620
rect 22032 50560 22096 50564
rect 22112 50620 22176 50624
rect 22112 50564 22116 50620
rect 22116 50564 22172 50620
rect 22172 50564 22176 50620
rect 22112 50560 22176 50564
rect 22192 50620 22256 50624
rect 22192 50564 22196 50620
rect 22196 50564 22252 50620
rect 22252 50564 22256 50620
rect 22192 50560 22256 50564
rect 26952 50620 27016 50624
rect 26952 50564 26956 50620
rect 26956 50564 27012 50620
rect 27012 50564 27016 50620
rect 26952 50560 27016 50564
rect 27032 50620 27096 50624
rect 27032 50564 27036 50620
rect 27036 50564 27092 50620
rect 27092 50564 27096 50620
rect 27032 50560 27096 50564
rect 27112 50620 27176 50624
rect 27112 50564 27116 50620
rect 27116 50564 27172 50620
rect 27172 50564 27176 50620
rect 27112 50560 27176 50564
rect 27192 50620 27256 50624
rect 27192 50564 27196 50620
rect 27196 50564 27252 50620
rect 27252 50564 27256 50620
rect 27192 50560 27256 50564
rect 31952 50620 32016 50624
rect 31952 50564 31956 50620
rect 31956 50564 32012 50620
rect 32012 50564 32016 50620
rect 31952 50560 32016 50564
rect 32032 50620 32096 50624
rect 32032 50564 32036 50620
rect 32036 50564 32092 50620
rect 32092 50564 32096 50620
rect 32032 50560 32096 50564
rect 32112 50620 32176 50624
rect 32112 50564 32116 50620
rect 32116 50564 32172 50620
rect 32172 50564 32176 50620
rect 32112 50560 32176 50564
rect 32192 50620 32256 50624
rect 32192 50564 32196 50620
rect 32196 50564 32252 50620
rect 32252 50564 32256 50620
rect 32192 50560 32256 50564
rect 36952 50620 37016 50624
rect 36952 50564 36956 50620
rect 36956 50564 37012 50620
rect 37012 50564 37016 50620
rect 36952 50560 37016 50564
rect 37032 50620 37096 50624
rect 37032 50564 37036 50620
rect 37036 50564 37092 50620
rect 37092 50564 37096 50620
rect 37032 50560 37096 50564
rect 37112 50620 37176 50624
rect 37112 50564 37116 50620
rect 37116 50564 37172 50620
rect 37172 50564 37176 50620
rect 37112 50560 37176 50564
rect 37192 50620 37256 50624
rect 37192 50564 37196 50620
rect 37196 50564 37252 50620
rect 37252 50564 37256 50620
rect 37192 50560 37256 50564
rect 2612 50076 2676 50080
rect 2612 50020 2616 50076
rect 2616 50020 2672 50076
rect 2672 50020 2676 50076
rect 2612 50016 2676 50020
rect 2692 50076 2756 50080
rect 2692 50020 2696 50076
rect 2696 50020 2752 50076
rect 2752 50020 2756 50076
rect 2692 50016 2756 50020
rect 2772 50076 2836 50080
rect 2772 50020 2776 50076
rect 2776 50020 2832 50076
rect 2832 50020 2836 50076
rect 2772 50016 2836 50020
rect 2852 50076 2916 50080
rect 2852 50020 2856 50076
rect 2856 50020 2912 50076
rect 2912 50020 2916 50076
rect 2852 50016 2916 50020
rect 7612 50076 7676 50080
rect 7612 50020 7616 50076
rect 7616 50020 7672 50076
rect 7672 50020 7676 50076
rect 7612 50016 7676 50020
rect 7692 50076 7756 50080
rect 7692 50020 7696 50076
rect 7696 50020 7752 50076
rect 7752 50020 7756 50076
rect 7692 50016 7756 50020
rect 7772 50076 7836 50080
rect 7772 50020 7776 50076
rect 7776 50020 7832 50076
rect 7832 50020 7836 50076
rect 7772 50016 7836 50020
rect 7852 50076 7916 50080
rect 7852 50020 7856 50076
rect 7856 50020 7912 50076
rect 7912 50020 7916 50076
rect 7852 50016 7916 50020
rect 12612 50076 12676 50080
rect 12612 50020 12616 50076
rect 12616 50020 12672 50076
rect 12672 50020 12676 50076
rect 12612 50016 12676 50020
rect 12692 50076 12756 50080
rect 12692 50020 12696 50076
rect 12696 50020 12752 50076
rect 12752 50020 12756 50076
rect 12692 50016 12756 50020
rect 12772 50076 12836 50080
rect 12772 50020 12776 50076
rect 12776 50020 12832 50076
rect 12832 50020 12836 50076
rect 12772 50016 12836 50020
rect 12852 50076 12916 50080
rect 12852 50020 12856 50076
rect 12856 50020 12912 50076
rect 12912 50020 12916 50076
rect 12852 50016 12916 50020
rect 17612 50076 17676 50080
rect 17612 50020 17616 50076
rect 17616 50020 17672 50076
rect 17672 50020 17676 50076
rect 17612 50016 17676 50020
rect 17692 50076 17756 50080
rect 17692 50020 17696 50076
rect 17696 50020 17752 50076
rect 17752 50020 17756 50076
rect 17692 50016 17756 50020
rect 17772 50076 17836 50080
rect 17772 50020 17776 50076
rect 17776 50020 17832 50076
rect 17832 50020 17836 50076
rect 17772 50016 17836 50020
rect 17852 50076 17916 50080
rect 17852 50020 17856 50076
rect 17856 50020 17912 50076
rect 17912 50020 17916 50076
rect 17852 50016 17916 50020
rect 22612 50076 22676 50080
rect 22612 50020 22616 50076
rect 22616 50020 22672 50076
rect 22672 50020 22676 50076
rect 22612 50016 22676 50020
rect 22692 50076 22756 50080
rect 22692 50020 22696 50076
rect 22696 50020 22752 50076
rect 22752 50020 22756 50076
rect 22692 50016 22756 50020
rect 22772 50076 22836 50080
rect 22772 50020 22776 50076
rect 22776 50020 22832 50076
rect 22832 50020 22836 50076
rect 22772 50016 22836 50020
rect 22852 50076 22916 50080
rect 22852 50020 22856 50076
rect 22856 50020 22912 50076
rect 22912 50020 22916 50076
rect 22852 50016 22916 50020
rect 27612 50076 27676 50080
rect 27612 50020 27616 50076
rect 27616 50020 27672 50076
rect 27672 50020 27676 50076
rect 27612 50016 27676 50020
rect 27692 50076 27756 50080
rect 27692 50020 27696 50076
rect 27696 50020 27752 50076
rect 27752 50020 27756 50076
rect 27692 50016 27756 50020
rect 27772 50076 27836 50080
rect 27772 50020 27776 50076
rect 27776 50020 27832 50076
rect 27832 50020 27836 50076
rect 27772 50016 27836 50020
rect 27852 50076 27916 50080
rect 27852 50020 27856 50076
rect 27856 50020 27912 50076
rect 27912 50020 27916 50076
rect 27852 50016 27916 50020
rect 32612 50076 32676 50080
rect 32612 50020 32616 50076
rect 32616 50020 32672 50076
rect 32672 50020 32676 50076
rect 32612 50016 32676 50020
rect 32692 50076 32756 50080
rect 32692 50020 32696 50076
rect 32696 50020 32752 50076
rect 32752 50020 32756 50076
rect 32692 50016 32756 50020
rect 32772 50076 32836 50080
rect 32772 50020 32776 50076
rect 32776 50020 32832 50076
rect 32832 50020 32836 50076
rect 32772 50016 32836 50020
rect 32852 50076 32916 50080
rect 32852 50020 32856 50076
rect 32856 50020 32912 50076
rect 32912 50020 32916 50076
rect 32852 50016 32916 50020
rect 37612 50076 37676 50080
rect 37612 50020 37616 50076
rect 37616 50020 37672 50076
rect 37672 50020 37676 50076
rect 37612 50016 37676 50020
rect 37692 50076 37756 50080
rect 37692 50020 37696 50076
rect 37696 50020 37752 50076
rect 37752 50020 37756 50076
rect 37692 50016 37756 50020
rect 37772 50076 37836 50080
rect 37772 50020 37776 50076
rect 37776 50020 37832 50076
rect 37832 50020 37836 50076
rect 37772 50016 37836 50020
rect 37852 50076 37916 50080
rect 37852 50020 37856 50076
rect 37856 50020 37912 50076
rect 37912 50020 37916 50076
rect 37852 50016 37916 50020
rect 1952 49532 2016 49536
rect 1952 49476 1956 49532
rect 1956 49476 2012 49532
rect 2012 49476 2016 49532
rect 1952 49472 2016 49476
rect 2032 49532 2096 49536
rect 2032 49476 2036 49532
rect 2036 49476 2092 49532
rect 2092 49476 2096 49532
rect 2032 49472 2096 49476
rect 2112 49532 2176 49536
rect 2112 49476 2116 49532
rect 2116 49476 2172 49532
rect 2172 49476 2176 49532
rect 2112 49472 2176 49476
rect 2192 49532 2256 49536
rect 2192 49476 2196 49532
rect 2196 49476 2252 49532
rect 2252 49476 2256 49532
rect 2192 49472 2256 49476
rect 6952 49532 7016 49536
rect 6952 49476 6956 49532
rect 6956 49476 7012 49532
rect 7012 49476 7016 49532
rect 6952 49472 7016 49476
rect 7032 49532 7096 49536
rect 7032 49476 7036 49532
rect 7036 49476 7092 49532
rect 7092 49476 7096 49532
rect 7032 49472 7096 49476
rect 7112 49532 7176 49536
rect 7112 49476 7116 49532
rect 7116 49476 7172 49532
rect 7172 49476 7176 49532
rect 7112 49472 7176 49476
rect 7192 49532 7256 49536
rect 7192 49476 7196 49532
rect 7196 49476 7252 49532
rect 7252 49476 7256 49532
rect 7192 49472 7256 49476
rect 11952 49532 12016 49536
rect 11952 49476 11956 49532
rect 11956 49476 12012 49532
rect 12012 49476 12016 49532
rect 11952 49472 12016 49476
rect 12032 49532 12096 49536
rect 12032 49476 12036 49532
rect 12036 49476 12092 49532
rect 12092 49476 12096 49532
rect 12032 49472 12096 49476
rect 12112 49532 12176 49536
rect 12112 49476 12116 49532
rect 12116 49476 12172 49532
rect 12172 49476 12176 49532
rect 12112 49472 12176 49476
rect 12192 49532 12256 49536
rect 12192 49476 12196 49532
rect 12196 49476 12252 49532
rect 12252 49476 12256 49532
rect 12192 49472 12256 49476
rect 16952 49532 17016 49536
rect 16952 49476 16956 49532
rect 16956 49476 17012 49532
rect 17012 49476 17016 49532
rect 16952 49472 17016 49476
rect 17032 49532 17096 49536
rect 17032 49476 17036 49532
rect 17036 49476 17092 49532
rect 17092 49476 17096 49532
rect 17032 49472 17096 49476
rect 17112 49532 17176 49536
rect 17112 49476 17116 49532
rect 17116 49476 17172 49532
rect 17172 49476 17176 49532
rect 17112 49472 17176 49476
rect 17192 49532 17256 49536
rect 17192 49476 17196 49532
rect 17196 49476 17252 49532
rect 17252 49476 17256 49532
rect 17192 49472 17256 49476
rect 21952 49532 22016 49536
rect 21952 49476 21956 49532
rect 21956 49476 22012 49532
rect 22012 49476 22016 49532
rect 21952 49472 22016 49476
rect 22032 49532 22096 49536
rect 22032 49476 22036 49532
rect 22036 49476 22092 49532
rect 22092 49476 22096 49532
rect 22032 49472 22096 49476
rect 22112 49532 22176 49536
rect 22112 49476 22116 49532
rect 22116 49476 22172 49532
rect 22172 49476 22176 49532
rect 22112 49472 22176 49476
rect 22192 49532 22256 49536
rect 22192 49476 22196 49532
rect 22196 49476 22252 49532
rect 22252 49476 22256 49532
rect 22192 49472 22256 49476
rect 26952 49532 27016 49536
rect 26952 49476 26956 49532
rect 26956 49476 27012 49532
rect 27012 49476 27016 49532
rect 26952 49472 27016 49476
rect 27032 49532 27096 49536
rect 27032 49476 27036 49532
rect 27036 49476 27092 49532
rect 27092 49476 27096 49532
rect 27032 49472 27096 49476
rect 27112 49532 27176 49536
rect 27112 49476 27116 49532
rect 27116 49476 27172 49532
rect 27172 49476 27176 49532
rect 27112 49472 27176 49476
rect 27192 49532 27256 49536
rect 27192 49476 27196 49532
rect 27196 49476 27252 49532
rect 27252 49476 27256 49532
rect 27192 49472 27256 49476
rect 31952 49532 32016 49536
rect 31952 49476 31956 49532
rect 31956 49476 32012 49532
rect 32012 49476 32016 49532
rect 31952 49472 32016 49476
rect 32032 49532 32096 49536
rect 32032 49476 32036 49532
rect 32036 49476 32092 49532
rect 32092 49476 32096 49532
rect 32032 49472 32096 49476
rect 32112 49532 32176 49536
rect 32112 49476 32116 49532
rect 32116 49476 32172 49532
rect 32172 49476 32176 49532
rect 32112 49472 32176 49476
rect 32192 49532 32256 49536
rect 32192 49476 32196 49532
rect 32196 49476 32252 49532
rect 32252 49476 32256 49532
rect 32192 49472 32256 49476
rect 36952 49532 37016 49536
rect 36952 49476 36956 49532
rect 36956 49476 37012 49532
rect 37012 49476 37016 49532
rect 36952 49472 37016 49476
rect 37032 49532 37096 49536
rect 37032 49476 37036 49532
rect 37036 49476 37092 49532
rect 37092 49476 37096 49532
rect 37032 49472 37096 49476
rect 37112 49532 37176 49536
rect 37112 49476 37116 49532
rect 37116 49476 37172 49532
rect 37172 49476 37176 49532
rect 37112 49472 37176 49476
rect 37192 49532 37256 49536
rect 37192 49476 37196 49532
rect 37196 49476 37252 49532
rect 37252 49476 37256 49532
rect 37192 49472 37256 49476
rect 2612 48988 2676 48992
rect 2612 48932 2616 48988
rect 2616 48932 2672 48988
rect 2672 48932 2676 48988
rect 2612 48928 2676 48932
rect 2692 48988 2756 48992
rect 2692 48932 2696 48988
rect 2696 48932 2752 48988
rect 2752 48932 2756 48988
rect 2692 48928 2756 48932
rect 2772 48988 2836 48992
rect 2772 48932 2776 48988
rect 2776 48932 2832 48988
rect 2832 48932 2836 48988
rect 2772 48928 2836 48932
rect 2852 48988 2916 48992
rect 2852 48932 2856 48988
rect 2856 48932 2912 48988
rect 2912 48932 2916 48988
rect 2852 48928 2916 48932
rect 7612 48988 7676 48992
rect 7612 48932 7616 48988
rect 7616 48932 7672 48988
rect 7672 48932 7676 48988
rect 7612 48928 7676 48932
rect 7692 48988 7756 48992
rect 7692 48932 7696 48988
rect 7696 48932 7752 48988
rect 7752 48932 7756 48988
rect 7692 48928 7756 48932
rect 7772 48988 7836 48992
rect 7772 48932 7776 48988
rect 7776 48932 7832 48988
rect 7832 48932 7836 48988
rect 7772 48928 7836 48932
rect 7852 48988 7916 48992
rect 7852 48932 7856 48988
rect 7856 48932 7912 48988
rect 7912 48932 7916 48988
rect 7852 48928 7916 48932
rect 12612 48988 12676 48992
rect 12612 48932 12616 48988
rect 12616 48932 12672 48988
rect 12672 48932 12676 48988
rect 12612 48928 12676 48932
rect 12692 48988 12756 48992
rect 12692 48932 12696 48988
rect 12696 48932 12752 48988
rect 12752 48932 12756 48988
rect 12692 48928 12756 48932
rect 12772 48988 12836 48992
rect 12772 48932 12776 48988
rect 12776 48932 12832 48988
rect 12832 48932 12836 48988
rect 12772 48928 12836 48932
rect 12852 48988 12916 48992
rect 12852 48932 12856 48988
rect 12856 48932 12912 48988
rect 12912 48932 12916 48988
rect 12852 48928 12916 48932
rect 17612 48988 17676 48992
rect 17612 48932 17616 48988
rect 17616 48932 17672 48988
rect 17672 48932 17676 48988
rect 17612 48928 17676 48932
rect 17692 48988 17756 48992
rect 17692 48932 17696 48988
rect 17696 48932 17752 48988
rect 17752 48932 17756 48988
rect 17692 48928 17756 48932
rect 17772 48988 17836 48992
rect 17772 48932 17776 48988
rect 17776 48932 17832 48988
rect 17832 48932 17836 48988
rect 17772 48928 17836 48932
rect 17852 48988 17916 48992
rect 17852 48932 17856 48988
rect 17856 48932 17912 48988
rect 17912 48932 17916 48988
rect 17852 48928 17916 48932
rect 22612 48988 22676 48992
rect 22612 48932 22616 48988
rect 22616 48932 22672 48988
rect 22672 48932 22676 48988
rect 22612 48928 22676 48932
rect 22692 48988 22756 48992
rect 22692 48932 22696 48988
rect 22696 48932 22752 48988
rect 22752 48932 22756 48988
rect 22692 48928 22756 48932
rect 22772 48988 22836 48992
rect 22772 48932 22776 48988
rect 22776 48932 22832 48988
rect 22832 48932 22836 48988
rect 22772 48928 22836 48932
rect 22852 48988 22916 48992
rect 22852 48932 22856 48988
rect 22856 48932 22912 48988
rect 22912 48932 22916 48988
rect 22852 48928 22916 48932
rect 27612 48988 27676 48992
rect 27612 48932 27616 48988
rect 27616 48932 27672 48988
rect 27672 48932 27676 48988
rect 27612 48928 27676 48932
rect 27692 48988 27756 48992
rect 27692 48932 27696 48988
rect 27696 48932 27752 48988
rect 27752 48932 27756 48988
rect 27692 48928 27756 48932
rect 27772 48988 27836 48992
rect 27772 48932 27776 48988
rect 27776 48932 27832 48988
rect 27832 48932 27836 48988
rect 27772 48928 27836 48932
rect 27852 48988 27916 48992
rect 27852 48932 27856 48988
rect 27856 48932 27912 48988
rect 27912 48932 27916 48988
rect 27852 48928 27916 48932
rect 32612 48988 32676 48992
rect 32612 48932 32616 48988
rect 32616 48932 32672 48988
rect 32672 48932 32676 48988
rect 32612 48928 32676 48932
rect 32692 48988 32756 48992
rect 32692 48932 32696 48988
rect 32696 48932 32752 48988
rect 32752 48932 32756 48988
rect 32692 48928 32756 48932
rect 32772 48988 32836 48992
rect 32772 48932 32776 48988
rect 32776 48932 32832 48988
rect 32832 48932 32836 48988
rect 32772 48928 32836 48932
rect 32852 48988 32916 48992
rect 32852 48932 32856 48988
rect 32856 48932 32912 48988
rect 32912 48932 32916 48988
rect 32852 48928 32916 48932
rect 37612 48988 37676 48992
rect 37612 48932 37616 48988
rect 37616 48932 37672 48988
rect 37672 48932 37676 48988
rect 37612 48928 37676 48932
rect 37692 48988 37756 48992
rect 37692 48932 37696 48988
rect 37696 48932 37752 48988
rect 37752 48932 37756 48988
rect 37692 48928 37756 48932
rect 37772 48988 37836 48992
rect 37772 48932 37776 48988
rect 37776 48932 37832 48988
rect 37832 48932 37836 48988
rect 37772 48928 37836 48932
rect 37852 48988 37916 48992
rect 37852 48932 37856 48988
rect 37856 48932 37912 48988
rect 37912 48932 37916 48988
rect 37852 48928 37916 48932
rect 1952 48444 2016 48448
rect 1952 48388 1956 48444
rect 1956 48388 2012 48444
rect 2012 48388 2016 48444
rect 1952 48384 2016 48388
rect 2032 48444 2096 48448
rect 2032 48388 2036 48444
rect 2036 48388 2092 48444
rect 2092 48388 2096 48444
rect 2032 48384 2096 48388
rect 2112 48444 2176 48448
rect 2112 48388 2116 48444
rect 2116 48388 2172 48444
rect 2172 48388 2176 48444
rect 2112 48384 2176 48388
rect 2192 48444 2256 48448
rect 2192 48388 2196 48444
rect 2196 48388 2252 48444
rect 2252 48388 2256 48444
rect 2192 48384 2256 48388
rect 6952 48444 7016 48448
rect 6952 48388 6956 48444
rect 6956 48388 7012 48444
rect 7012 48388 7016 48444
rect 6952 48384 7016 48388
rect 7032 48444 7096 48448
rect 7032 48388 7036 48444
rect 7036 48388 7092 48444
rect 7092 48388 7096 48444
rect 7032 48384 7096 48388
rect 7112 48444 7176 48448
rect 7112 48388 7116 48444
rect 7116 48388 7172 48444
rect 7172 48388 7176 48444
rect 7112 48384 7176 48388
rect 7192 48444 7256 48448
rect 7192 48388 7196 48444
rect 7196 48388 7252 48444
rect 7252 48388 7256 48444
rect 7192 48384 7256 48388
rect 11952 48444 12016 48448
rect 11952 48388 11956 48444
rect 11956 48388 12012 48444
rect 12012 48388 12016 48444
rect 11952 48384 12016 48388
rect 12032 48444 12096 48448
rect 12032 48388 12036 48444
rect 12036 48388 12092 48444
rect 12092 48388 12096 48444
rect 12032 48384 12096 48388
rect 12112 48444 12176 48448
rect 12112 48388 12116 48444
rect 12116 48388 12172 48444
rect 12172 48388 12176 48444
rect 12112 48384 12176 48388
rect 12192 48444 12256 48448
rect 12192 48388 12196 48444
rect 12196 48388 12252 48444
rect 12252 48388 12256 48444
rect 12192 48384 12256 48388
rect 16952 48444 17016 48448
rect 16952 48388 16956 48444
rect 16956 48388 17012 48444
rect 17012 48388 17016 48444
rect 16952 48384 17016 48388
rect 17032 48444 17096 48448
rect 17032 48388 17036 48444
rect 17036 48388 17092 48444
rect 17092 48388 17096 48444
rect 17032 48384 17096 48388
rect 17112 48444 17176 48448
rect 17112 48388 17116 48444
rect 17116 48388 17172 48444
rect 17172 48388 17176 48444
rect 17112 48384 17176 48388
rect 17192 48444 17256 48448
rect 17192 48388 17196 48444
rect 17196 48388 17252 48444
rect 17252 48388 17256 48444
rect 17192 48384 17256 48388
rect 21952 48444 22016 48448
rect 21952 48388 21956 48444
rect 21956 48388 22012 48444
rect 22012 48388 22016 48444
rect 21952 48384 22016 48388
rect 22032 48444 22096 48448
rect 22032 48388 22036 48444
rect 22036 48388 22092 48444
rect 22092 48388 22096 48444
rect 22032 48384 22096 48388
rect 22112 48444 22176 48448
rect 22112 48388 22116 48444
rect 22116 48388 22172 48444
rect 22172 48388 22176 48444
rect 22112 48384 22176 48388
rect 22192 48444 22256 48448
rect 22192 48388 22196 48444
rect 22196 48388 22252 48444
rect 22252 48388 22256 48444
rect 22192 48384 22256 48388
rect 26952 48444 27016 48448
rect 26952 48388 26956 48444
rect 26956 48388 27012 48444
rect 27012 48388 27016 48444
rect 26952 48384 27016 48388
rect 27032 48444 27096 48448
rect 27032 48388 27036 48444
rect 27036 48388 27092 48444
rect 27092 48388 27096 48444
rect 27032 48384 27096 48388
rect 27112 48444 27176 48448
rect 27112 48388 27116 48444
rect 27116 48388 27172 48444
rect 27172 48388 27176 48444
rect 27112 48384 27176 48388
rect 27192 48444 27256 48448
rect 27192 48388 27196 48444
rect 27196 48388 27252 48444
rect 27252 48388 27256 48444
rect 27192 48384 27256 48388
rect 31952 48444 32016 48448
rect 31952 48388 31956 48444
rect 31956 48388 32012 48444
rect 32012 48388 32016 48444
rect 31952 48384 32016 48388
rect 32032 48444 32096 48448
rect 32032 48388 32036 48444
rect 32036 48388 32092 48444
rect 32092 48388 32096 48444
rect 32032 48384 32096 48388
rect 32112 48444 32176 48448
rect 32112 48388 32116 48444
rect 32116 48388 32172 48444
rect 32172 48388 32176 48444
rect 32112 48384 32176 48388
rect 32192 48444 32256 48448
rect 32192 48388 32196 48444
rect 32196 48388 32252 48444
rect 32252 48388 32256 48444
rect 32192 48384 32256 48388
rect 36952 48444 37016 48448
rect 36952 48388 36956 48444
rect 36956 48388 37012 48444
rect 37012 48388 37016 48444
rect 36952 48384 37016 48388
rect 37032 48444 37096 48448
rect 37032 48388 37036 48444
rect 37036 48388 37092 48444
rect 37092 48388 37096 48444
rect 37032 48384 37096 48388
rect 37112 48444 37176 48448
rect 37112 48388 37116 48444
rect 37116 48388 37172 48444
rect 37172 48388 37176 48444
rect 37112 48384 37176 48388
rect 37192 48444 37256 48448
rect 37192 48388 37196 48444
rect 37196 48388 37252 48444
rect 37252 48388 37256 48444
rect 37192 48384 37256 48388
rect 2612 47900 2676 47904
rect 2612 47844 2616 47900
rect 2616 47844 2672 47900
rect 2672 47844 2676 47900
rect 2612 47840 2676 47844
rect 2692 47900 2756 47904
rect 2692 47844 2696 47900
rect 2696 47844 2752 47900
rect 2752 47844 2756 47900
rect 2692 47840 2756 47844
rect 2772 47900 2836 47904
rect 2772 47844 2776 47900
rect 2776 47844 2832 47900
rect 2832 47844 2836 47900
rect 2772 47840 2836 47844
rect 2852 47900 2916 47904
rect 2852 47844 2856 47900
rect 2856 47844 2912 47900
rect 2912 47844 2916 47900
rect 2852 47840 2916 47844
rect 7612 47900 7676 47904
rect 7612 47844 7616 47900
rect 7616 47844 7672 47900
rect 7672 47844 7676 47900
rect 7612 47840 7676 47844
rect 7692 47900 7756 47904
rect 7692 47844 7696 47900
rect 7696 47844 7752 47900
rect 7752 47844 7756 47900
rect 7692 47840 7756 47844
rect 7772 47900 7836 47904
rect 7772 47844 7776 47900
rect 7776 47844 7832 47900
rect 7832 47844 7836 47900
rect 7772 47840 7836 47844
rect 7852 47900 7916 47904
rect 7852 47844 7856 47900
rect 7856 47844 7912 47900
rect 7912 47844 7916 47900
rect 7852 47840 7916 47844
rect 12612 47900 12676 47904
rect 12612 47844 12616 47900
rect 12616 47844 12672 47900
rect 12672 47844 12676 47900
rect 12612 47840 12676 47844
rect 12692 47900 12756 47904
rect 12692 47844 12696 47900
rect 12696 47844 12752 47900
rect 12752 47844 12756 47900
rect 12692 47840 12756 47844
rect 12772 47900 12836 47904
rect 12772 47844 12776 47900
rect 12776 47844 12832 47900
rect 12832 47844 12836 47900
rect 12772 47840 12836 47844
rect 12852 47900 12916 47904
rect 12852 47844 12856 47900
rect 12856 47844 12912 47900
rect 12912 47844 12916 47900
rect 12852 47840 12916 47844
rect 17612 47900 17676 47904
rect 17612 47844 17616 47900
rect 17616 47844 17672 47900
rect 17672 47844 17676 47900
rect 17612 47840 17676 47844
rect 17692 47900 17756 47904
rect 17692 47844 17696 47900
rect 17696 47844 17752 47900
rect 17752 47844 17756 47900
rect 17692 47840 17756 47844
rect 17772 47900 17836 47904
rect 17772 47844 17776 47900
rect 17776 47844 17832 47900
rect 17832 47844 17836 47900
rect 17772 47840 17836 47844
rect 17852 47900 17916 47904
rect 17852 47844 17856 47900
rect 17856 47844 17912 47900
rect 17912 47844 17916 47900
rect 17852 47840 17916 47844
rect 22612 47900 22676 47904
rect 22612 47844 22616 47900
rect 22616 47844 22672 47900
rect 22672 47844 22676 47900
rect 22612 47840 22676 47844
rect 22692 47900 22756 47904
rect 22692 47844 22696 47900
rect 22696 47844 22752 47900
rect 22752 47844 22756 47900
rect 22692 47840 22756 47844
rect 22772 47900 22836 47904
rect 22772 47844 22776 47900
rect 22776 47844 22832 47900
rect 22832 47844 22836 47900
rect 22772 47840 22836 47844
rect 22852 47900 22916 47904
rect 22852 47844 22856 47900
rect 22856 47844 22912 47900
rect 22912 47844 22916 47900
rect 22852 47840 22916 47844
rect 27612 47900 27676 47904
rect 27612 47844 27616 47900
rect 27616 47844 27672 47900
rect 27672 47844 27676 47900
rect 27612 47840 27676 47844
rect 27692 47900 27756 47904
rect 27692 47844 27696 47900
rect 27696 47844 27752 47900
rect 27752 47844 27756 47900
rect 27692 47840 27756 47844
rect 27772 47900 27836 47904
rect 27772 47844 27776 47900
rect 27776 47844 27832 47900
rect 27832 47844 27836 47900
rect 27772 47840 27836 47844
rect 27852 47900 27916 47904
rect 27852 47844 27856 47900
rect 27856 47844 27912 47900
rect 27912 47844 27916 47900
rect 27852 47840 27916 47844
rect 32612 47900 32676 47904
rect 32612 47844 32616 47900
rect 32616 47844 32672 47900
rect 32672 47844 32676 47900
rect 32612 47840 32676 47844
rect 32692 47900 32756 47904
rect 32692 47844 32696 47900
rect 32696 47844 32752 47900
rect 32752 47844 32756 47900
rect 32692 47840 32756 47844
rect 32772 47900 32836 47904
rect 32772 47844 32776 47900
rect 32776 47844 32832 47900
rect 32832 47844 32836 47900
rect 32772 47840 32836 47844
rect 32852 47900 32916 47904
rect 32852 47844 32856 47900
rect 32856 47844 32912 47900
rect 32912 47844 32916 47900
rect 32852 47840 32916 47844
rect 37612 47900 37676 47904
rect 37612 47844 37616 47900
rect 37616 47844 37672 47900
rect 37672 47844 37676 47900
rect 37612 47840 37676 47844
rect 37692 47900 37756 47904
rect 37692 47844 37696 47900
rect 37696 47844 37752 47900
rect 37752 47844 37756 47900
rect 37692 47840 37756 47844
rect 37772 47900 37836 47904
rect 37772 47844 37776 47900
rect 37776 47844 37832 47900
rect 37832 47844 37836 47900
rect 37772 47840 37836 47844
rect 37852 47900 37916 47904
rect 37852 47844 37856 47900
rect 37856 47844 37912 47900
rect 37912 47844 37916 47900
rect 37852 47840 37916 47844
rect 1952 47356 2016 47360
rect 1952 47300 1956 47356
rect 1956 47300 2012 47356
rect 2012 47300 2016 47356
rect 1952 47296 2016 47300
rect 2032 47356 2096 47360
rect 2032 47300 2036 47356
rect 2036 47300 2092 47356
rect 2092 47300 2096 47356
rect 2032 47296 2096 47300
rect 2112 47356 2176 47360
rect 2112 47300 2116 47356
rect 2116 47300 2172 47356
rect 2172 47300 2176 47356
rect 2112 47296 2176 47300
rect 2192 47356 2256 47360
rect 2192 47300 2196 47356
rect 2196 47300 2252 47356
rect 2252 47300 2256 47356
rect 2192 47296 2256 47300
rect 6952 47356 7016 47360
rect 6952 47300 6956 47356
rect 6956 47300 7012 47356
rect 7012 47300 7016 47356
rect 6952 47296 7016 47300
rect 7032 47356 7096 47360
rect 7032 47300 7036 47356
rect 7036 47300 7092 47356
rect 7092 47300 7096 47356
rect 7032 47296 7096 47300
rect 7112 47356 7176 47360
rect 7112 47300 7116 47356
rect 7116 47300 7172 47356
rect 7172 47300 7176 47356
rect 7112 47296 7176 47300
rect 7192 47356 7256 47360
rect 7192 47300 7196 47356
rect 7196 47300 7252 47356
rect 7252 47300 7256 47356
rect 7192 47296 7256 47300
rect 11952 47356 12016 47360
rect 11952 47300 11956 47356
rect 11956 47300 12012 47356
rect 12012 47300 12016 47356
rect 11952 47296 12016 47300
rect 12032 47356 12096 47360
rect 12032 47300 12036 47356
rect 12036 47300 12092 47356
rect 12092 47300 12096 47356
rect 12032 47296 12096 47300
rect 12112 47356 12176 47360
rect 12112 47300 12116 47356
rect 12116 47300 12172 47356
rect 12172 47300 12176 47356
rect 12112 47296 12176 47300
rect 12192 47356 12256 47360
rect 12192 47300 12196 47356
rect 12196 47300 12252 47356
rect 12252 47300 12256 47356
rect 12192 47296 12256 47300
rect 16952 47356 17016 47360
rect 16952 47300 16956 47356
rect 16956 47300 17012 47356
rect 17012 47300 17016 47356
rect 16952 47296 17016 47300
rect 17032 47356 17096 47360
rect 17032 47300 17036 47356
rect 17036 47300 17092 47356
rect 17092 47300 17096 47356
rect 17032 47296 17096 47300
rect 17112 47356 17176 47360
rect 17112 47300 17116 47356
rect 17116 47300 17172 47356
rect 17172 47300 17176 47356
rect 17112 47296 17176 47300
rect 17192 47356 17256 47360
rect 17192 47300 17196 47356
rect 17196 47300 17252 47356
rect 17252 47300 17256 47356
rect 17192 47296 17256 47300
rect 21952 47356 22016 47360
rect 21952 47300 21956 47356
rect 21956 47300 22012 47356
rect 22012 47300 22016 47356
rect 21952 47296 22016 47300
rect 22032 47356 22096 47360
rect 22032 47300 22036 47356
rect 22036 47300 22092 47356
rect 22092 47300 22096 47356
rect 22032 47296 22096 47300
rect 22112 47356 22176 47360
rect 22112 47300 22116 47356
rect 22116 47300 22172 47356
rect 22172 47300 22176 47356
rect 22112 47296 22176 47300
rect 22192 47356 22256 47360
rect 22192 47300 22196 47356
rect 22196 47300 22252 47356
rect 22252 47300 22256 47356
rect 22192 47296 22256 47300
rect 26952 47356 27016 47360
rect 26952 47300 26956 47356
rect 26956 47300 27012 47356
rect 27012 47300 27016 47356
rect 26952 47296 27016 47300
rect 27032 47356 27096 47360
rect 27032 47300 27036 47356
rect 27036 47300 27092 47356
rect 27092 47300 27096 47356
rect 27032 47296 27096 47300
rect 27112 47356 27176 47360
rect 27112 47300 27116 47356
rect 27116 47300 27172 47356
rect 27172 47300 27176 47356
rect 27112 47296 27176 47300
rect 27192 47356 27256 47360
rect 27192 47300 27196 47356
rect 27196 47300 27252 47356
rect 27252 47300 27256 47356
rect 27192 47296 27256 47300
rect 31952 47356 32016 47360
rect 31952 47300 31956 47356
rect 31956 47300 32012 47356
rect 32012 47300 32016 47356
rect 31952 47296 32016 47300
rect 32032 47356 32096 47360
rect 32032 47300 32036 47356
rect 32036 47300 32092 47356
rect 32092 47300 32096 47356
rect 32032 47296 32096 47300
rect 32112 47356 32176 47360
rect 32112 47300 32116 47356
rect 32116 47300 32172 47356
rect 32172 47300 32176 47356
rect 32112 47296 32176 47300
rect 32192 47356 32256 47360
rect 32192 47300 32196 47356
rect 32196 47300 32252 47356
rect 32252 47300 32256 47356
rect 32192 47296 32256 47300
rect 36952 47356 37016 47360
rect 36952 47300 36956 47356
rect 36956 47300 37012 47356
rect 37012 47300 37016 47356
rect 36952 47296 37016 47300
rect 37032 47356 37096 47360
rect 37032 47300 37036 47356
rect 37036 47300 37092 47356
rect 37092 47300 37096 47356
rect 37032 47296 37096 47300
rect 37112 47356 37176 47360
rect 37112 47300 37116 47356
rect 37116 47300 37172 47356
rect 37172 47300 37176 47356
rect 37112 47296 37176 47300
rect 37192 47356 37256 47360
rect 37192 47300 37196 47356
rect 37196 47300 37252 47356
rect 37252 47300 37256 47356
rect 37192 47296 37256 47300
rect 2612 46812 2676 46816
rect 2612 46756 2616 46812
rect 2616 46756 2672 46812
rect 2672 46756 2676 46812
rect 2612 46752 2676 46756
rect 2692 46812 2756 46816
rect 2692 46756 2696 46812
rect 2696 46756 2752 46812
rect 2752 46756 2756 46812
rect 2692 46752 2756 46756
rect 2772 46812 2836 46816
rect 2772 46756 2776 46812
rect 2776 46756 2832 46812
rect 2832 46756 2836 46812
rect 2772 46752 2836 46756
rect 2852 46812 2916 46816
rect 2852 46756 2856 46812
rect 2856 46756 2912 46812
rect 2912 46756 2916 46812
rect 2852 46752 2916 46756
rect 7612 46812 7676 46816
rect 7612 46756 7616 46812
rect 7616 46756 7672 46812
rect 7672 46756 7676 46812
rect 7612 46752 7676 46756
rect 7692 46812 7756 46816
rect 7692 46756 7696 46812
rect 7696 46756 7752 46812
rect 7752 46756 7756 46812
rect 7692 46752 7756 46756
rect 7772 46812 7836 46816
rect 7772 46756 7776 46812
rect 7776 46756 7832 46812
rect 7832 46756 7836 46812
rect 7772 46752 7836 46756
rect 7852 46812 7916 46816
rect 7852 46756 7856 46812
rect 7856 46756 7912 46812
rect 7912 46756 7916 46812
rect 7852 46752 7916 46756
rect 12612 46812 12676 46816
rect 12612 46756 12616 46812
rect 12616 46756 12672 46812
rect 12672 46756 12676 46812
rect 12612 46752 12676 46756
rect 12692 46812 12756 46816
rect 12692 46756 12696 46812
rect 12696 46756 12752 46812
rect 12752 46756 12756 46812
rect 12692 46752 12756 46756
rect 12772 46812 12836 46816
rect 12772 46756 12776 46812
rect 12776 46756 12832 46812
rect 12832 46756 12836 46812
rect 12772 46752 12836 46756
rect 12852 46812 12916 46816
rect 12852 46756 12856 46812
rect 12856 46756 12912 46812
rect 12912 46756 12916 46812
rect 12852 46752 12916 46756
rect 17612 46812 17676 46816
rect 17612 46756 17616 46812
rect 17616 46756 17672 46812
rect 17672 46756 17676 46812
rect 17612 46752 17676 46756
rect 17692 46812 17756 46816
rect 17692 46756 17696 46812
rect 17696 46756 17752 46812
rect 17752 46756 17756 46812
rect 17692 46752 17756 46756
rect 17772 46812 17836 46816
rect 17772 46756 17776 46812
rect 17776 46756 17832 46812
rect 17832 46756 17836 46812
rect 17772 46752 17836 46756
rect 17852 46812 17916 46816
rect 17852 46756 17856 46812
rect 17856 46756 17912 46812
rect 17912 46756 17916 46812
rect 17852 46752 17916 46756
rect 22612 46812 22676 46816
rect 22612 46756 22616 46812
rect 22616 46756 22672 46812
rect 22672 46756 22676 46812
rect 22612 46752 22676 46756
rect 22692 46812 22756 46816
rect 22692 46756 22696 46812
rect 22696 46756 22752 46812
rect 22752 46756 22756 46812
rect 22692 46752 22756 46756
rect 22772 46812 22836 46816
rect 22772 46756 22776 46812
rect 22776 46756 22832 46812
rect 22832 46756 22836 46812
rect 22772 46752 22836 46756
rect 22852 46812 22916 46816
rect 22852 46756 22856 46812
rect 22856 46756 22912 46812
rect 22912 46756 22916 46812
rect 22852 46752 22916 46756
rect 27612 46812 27676 46816
rect 27612 46756 27616 46812
rect 27616 46756 27672 46812
rect 27672 46756 27676 46812
rect 27612 46752 27676 46756
rect 27692 46812 27756 46816
rect 27692 46756 27696 46812
rect 27696 46756 27752 46812
rect 27752 46756 27756 46812
rect 27692 46752 27756 46756
rect 27772 46812 27836 46816
rect 27772 46756 27776 46812
rect 27776 46756 27832 46812
rect 27832 46756 27836 46812
rect 27772 46752 27836 46756
rect 27852 46812 27916 46816
rect 27852 46756 27856 46812
rect 27856 46756 27912 46812
rect 27912 46756 27916 46812
rect 27852 46752 27916 46756
rect 32612 46812 32676 46816
rect 32612 46756 32616 46812
rect 32616 46756 32672 46812
rect 32672 46756 32676 46812
rect 32612 46752 32676 46756
rect 32692 46812 32756 46816
rect 32692 46756 32696 46812
rect 32696 46756 32752 46812
rect 32752 46756 32756 46812
rect 32692 46752 32756 46756
rect 32772 46812 32836 46816
rect 32772 46756 32776 46812
rect 32776 46756 32832 46812
rect 32832 46756 32836 46812
rect 32772 46752 32836 46756
rect 32852 46812 32916 46816
rect 32852 46756 32856 46812
rect 32856 46756 32912 46812
rect 32912 46756 32916 46812
rect 32852 46752 32916 46756
rect 37612 46812 37676 46816
rect 37612 46756 37616 46812
rect 37616 46756 37672 46812
rect 37672 46756 37676 46812
rect 37612 46752 37676 46756
rect 37692 46812 37756 46816
rect 37692 46756 37696 46812
rect 37696 46756 37752 46812
rect 37752 46756 37756 46812
rect 37692 46752 37756 46756
rect 37772 46812 37836 46816
rect 37772 46756 37776 46812
rect 37776 46756 37832 46812
rect 37832 46756 37836 46812
rect 37772 46752 37836 46756
rect 37852 46812 37916 46816
rect 37852 46756 37856 46812
rect 37856 46756 37912 46812
rect 37912 46756 37916 46812
rect 37852 46752 37916 46756
rect 1952 46268 2016 46272
rect 1952 46212 1956 46268
rect 1956 46212 2012 46268
rect 2012 46212 2016 46268
rect 1952 46208 2016 46212
rect 2032 46268 2096 46272
rect 2032 46212 2036 46268
rect 2036 46212 2092 46268
rect 2092 46212 2096 46268
rect 2032 46208 2096 46212
rect 2112 46268 2176 46272
rect 2112 46212 2116 46268
rect 2116 46212 2172 46268
rect 2172 46212 2176 46268
rect 2112 46208 2176 46212
rect 2192 46268 2256 46272
rect 2192 46212 2196 46268
rect 2196 46212 2252 46268
rect 2252 46212 2256 46268
rect 2192 46208 2256 46212
rect 6952 46268 7016 46272
rect 6952 46212 6956 46268
rect 6956 46212 7012 46268
rect 7012 46212 7016 46268
rect 6952 46208 7016 46212
rect 7032 46268 7096 46272
rect 7032 46212 7036 46268
rect 7036 46212 7092 46268
rect 7092 46212 7096 46268
rect 7032 46208 7096 46212
rect 7112 46268 7176 46272
rect 7112 46212 7116 46268
rect 7116 46212 7172 46268
rect 7172 46212 7176 46268
rect 7112 46208 7176 46212
rect 7192 46268 7256 46272
rect 7192 46212 7196 46268
rect 7196 46212 7252 46268
rect 7252 46212 7256 46268
rect 7192 46208 7256 46212
rect 11952 46268 12016 46272
rect 11952 46212 11956 46268
rect 11956 46212 12012 46268
rect 12012 46212 12016 46268
rect 11952 46208 12016 46212
rect 12032 46268 12096 46272
rect 12032 46212 12036 46268
rect 12036 46212 12092 46268
rect 12092 46212 12096 46268
rect 12032 46208 12096 46212
rect 12112 46268 12176 46272
rect 12112 46212 12116 46268
rect 12116 46212 12172 46268
rect 12172 46212 12176 46268
rect 12112 46208 12176 46212
rect 12192 46268 12256 46272
rect 12192 46212 12196 46268
rect 12196 46212 12252 46268
rect 12252 46212 12256 46268
rect 12192 46208 12256 46212
rect 16952 46268 17016 46272
rect 16952 46212 16956 46268
rect 16956 46212 17012 46268
rect 17012 46212 17016 46268
rect 16952 46208 17016 46212
rect 17032 46268 17096 46272
rect 17032 46212 17036 46268
rect 17036 46212 17092 46268
rect 17092 46212 17096 46268
rect 17032 46208 17096 46212
rect 17112 46268 17176 46272
rect 17112 46212 17116 46268
rect 17116 46212 17172 46268
rect 17172 46212 17176 46268
rect 17112 46208 17176 46212
rect 17192 46268 17256 46272
rect 17192 46212 17196 46268
rect 17196 46212 17252 46268
rect 17252 46212 17256 46268
rect 17192 46208 17256 46212
rect 21952 46268 22016 46272
rect 21952 46212 21956 46268
rect 21956 46212 22012 46268
rect 22012 46212 22016 46268
rect 21952 46208 22016 46212
rect 22032 46268 22096 46272
rect 22032 46212 22036 46268
rect 22036 46212 22092 46268
rect 22092 46212 22096 46268
rect 22032 46208 22096 46212
rect 22112 46268 22176 46272
rect 22112 46212 22116 46268
rect 22116 46212 22172 46268
rect 22172 46212 22176 46268
rect 22112 46208 22176 46212
rect 22192 46268 22256 46272
rect 22192 46212 22196 46268
rect 22196 46212 22252 46268
rect 22252 46212 22256 46268
rect 22192 46208 22256 46212
rect 26952 46268 27016 46272
rect 26952 46212 26956 46268
rect 26956 46212 27012 46268
rect 27012 46212 27016 46268
rect 26952 46208 27016 46212
rect 27032 46268 27096 46272
rect 27032 46212 27036 46268
rect 27036 46212 27092 46268
rect 27092 46212 27096 46268
rect 27032 46208 27096 46212
rect 27112 46268 27176 46272
rect 27112 46212 27116 46268
rect 27116 46212 27172 46268
rect 27172 46212 27176 46268
rect 27112 46208 27176 46212
rect 27192 46268 27256 46272
rect 27192 46212 27196 46268
rect 27196 46212 27252 46268
rect 27252 46212 27256 46268
rect 27192 46208 27256 46212
rect 31952 46268 32016 46272
rect 31952 46212 31956 46268
rect 31956 46212 32012 46268
rect 32012 46212 32016 46268
rect 31952 46208 32016 46212
rect 32032 46268 32096 46272
rect 32032 46212 32036 46268
rect 32036 46212 32092 46268
rect 32092 46212 32096 46268
rect 32032 46208 32096 46212
rect 32112 46268 32176 46272
rect 32112 46212 32116 46268
rect 32116 46212 32172 46268
rect 32172 46212 32176 46268
rect 32112 46208 32176 46212
rect 32192 46268 32256 46272
rect 32192 46212 32196 46268
rect 32196 46212 32252 46268
rect 32252 46212 32256 46268
rect 32192 46208 32256 46212
rect 36952 46268 37016 46272
rect 36952 46212 36956 46268
rect 36956 46212 37012 46268
rect 37012 46212 37016 46268
rect 36952 46208 37016 46212
rect 37032 46268 37096 46272
rect 37032 46212 37036 46268
rect 37036 46212 37092 46268
rect 37092 46212 37096 46268
rect 37032 46208 37096 46212
rect 37112 46268 37176 46272
rect 37112 46212 37116 46268
rect 37116 46212 37172 46268
rect 37172 46212 37176 46268
rect 37112 46208 37176 46212
rect 37192 46268 37256 46272
rect 37192 46212 37196 46268
rect 37196 46212 37252 46268
rect 37252 46212 37256 46268
rect 37192 46208 37256 46212
rect 2612 45724 2676 45728
rect 2612 45668 2616 45724
rect 2616 45668 2672 45724
rect 2672 45668 2676 45724
rect 2612 45664 2676 45668
rect 2692 45724 2756 45728
rect 2692 45668 2696 45724
rect 2696 45668 2752 45724
rect 2752 45668 2756 45724
rect 2692 45664 2756 45668
rect 2772 45724 2836 45728
rect 2772 45668 2776 45724
rect 2776 45668 2832 45724
rect 2832 45668 2836 45724
rect 2772 45664 2836 45668
rect 2852 45724 2916 45728
rect 2852 45668 2856 45724
rect 2856 45668 2912 45724
rect 2912 45668 2916 45724
rect 2852 45664 2916 45668
rect 7612 45724 7676 45728
rect 7612 45668 7616 45724
rect 7616 45668 7672 45724
rect 7672 45668 7676 45724
rect 7612 45664 7676 45668
rect 7692 45724 7756 45728
rect 7692 45668 7696 45724
rect 7696 45668 7752 45724
rect 7752 45668 7756 45724
rect 7692 45664 7756 45668
rect 7772 45724 7836 45728
rect 7772 45668 7776 45724
rect 7776 45668 7832 45724
rect 7832 45668 7836 45724
rect 7772 45664 7836 45668
rect 7852 45724 7916 45728
rect 7852 45668 7856 45724
rect 7856 45668 7912 45724
rect 7912 45668 7916 45724
rect 7852 45664 7916 45668
rect 12612 45724 12676 45728
rect 12612 45668 12616 45724
rect 12616 45668 12672 45724
rect 12672 45668 12676 45724
rect 12612 45664 12676 45668
rect 12692 45724 12756 45728
rect 12692 45668 12696 45724
rect 12696 45668 12752 45724
rect 12752 45668 12756 45724
rect 12692 45664 12756 45668
rect 12772 45724 12836 45728
rect 12772 45668 12776 45724
rect 12776 45668 12832 45724
rect 12832 45668 12836 45724
rect 12772 45664 12836 45668
rect 12852 45724 12916 45728
rect 12852 45668 12856 45724
rect 12856 45668 12912 45724
rect 12912 45668 12916 45724
rect 12852 45664 12916 45668
rect 17612 45724 17676 45728
rect 17612 45668 17616 45724
rect 17616 45668 17672 45724
rect 17672 45668 17676 45724
rect 17612 45664 17676 45668
rect 17692 45724 17756 45728
rect 17692 45668 17696 45724
rect 17696 45668 17752 45724
rect 17752 45668 17756 45724
rect 17692 45664 17756 45668
rect 17772 45724 17836 45728
rect 17772 45668 17776 45724
rect 17776 45668 17832 45724
rect 17832 45668 17836 45724
rect 17772 45664 17836 45668
rect 17852 45724 17916 45728
rect 17852 45668 17856 45724
rect 17856 45668 17912 45724
rect 17912 45668 17916 45724
rect 17852 45664 17916 45668
rect 22612 45724 22676 45728
rect 22612 45668 22616 45724
rect 22616 45668 22672 45724
rect 22672 45668 22676 45724
rect 22612 45664 22676 45668
rect 22692 45724 22756 45728
rect 22692 45668 22696 45724
rect 22696 45668 22752 45724
rect 22752 45668 22756 45724
rect 22692 45664 22756 45668
rect 22772 45724 22836 45728
rect 22772 45668 22776 45724
rect 22776 45668 22832 45724
rect 22832 45668 22836 45724
rect 22772 45664 22836 45668
rect 22852 45724 22916 45728
rect 22852 45668 22856 45724
rect 22856 45668 22912 45724
rect 22912 45668 22916 45724
rect 22852 45664 22916 45668
rect 27612 45724 27676 45728
rect 27612 45668 27616 45724
rect 27616 45668 27672 45724
rect 27672 45668 27676 45724
rect 27612 45664 27676 45668
rect 27692 45724 27756 45728
rect 27692 45668 27696 45724
rect 27696 45668 27752 45724
rect 27752 45668 27756 45724
rect 27692 45664 27756 45668
rect 27772 45724 27836 45728
rect 27772 45668 27776 45724
rect 27776 45668 27832 45724
rect 27832 45668 27836 45724
rect 27772 45664 27836 45668
rect 27852 45724 27916 45728
rect 27852 45668 27856 45724
rect 27856 45668 27912 45724
rect 27912 45668 27916 45724
rect 27852 45664 27916 45668
rect 32612 45724 32676 45728
rect 32612 45668 32616 45724
rect 32616 45668 32672 45724
rect 32672 45668 32676 45724
rect 32612 45664 32676 45668
rect 32692 45724 32756 45728
rect 32692 45668 32696 45724
rect 32696 45668 32752 45724
rect 32752 45668 32756 45724
rect 32692 45664 32756 45668
rect 32772 45724 32836 45728
rect 32772 45668 32776 45724
rect 32776 45668 32832 45724
rect 32832 45668 32836 45724
rect 32772 45664 32836 45668
rect 32852 45724 32916 45728
rect 32852 45668 32856 45724
rect 32856 45668 32912 45724
rect 32912 45668 32916 45724
rect 32852 45664 32916 45668
rect 37612 45724 37676 45728
rect 37612 45668 37616 45724
rect 37616 45668 37672 45724
rect 37672 45668 37676 45724
rect 37612 45664 37676 45668
rect 37692 45724 37756 45728
rect 37692 45668 37696 45724
rect 37696 45668 37752 45724
rect 37752 45668 37756 45724
rect 37692 45664 37756 45668
rect 37772 45724 37836 45728
rect 37772 45668 37776 45724
rect 37776 45668 37832 45724
rect 37832 45668 37836 45724
rect 37772 45664 37836 45668
rect 37852 45724 37916 45728
rect 37852 45668 37856 45724
rect 37856 45668 37912 45724
rect 37912 45668 37916 45724
rect 37852 45664 37916 45668
rect 1952 45180 2016 45184
rect 1952 45124 1956 45180
rect 1956 45124 2012 45180
rect 2012 45124 2016 45180
rect 1952 45120 2016 45124
rect 2032 45180 2096 45184
rect 2032 45124 2036 45180
rect 2036 45124 2092 45180
rect 2092 45124 2096 45180
rect 2032 45120 2096 45124
rect 2112 45180 2176 45184
rect 2112 45124 2116 45180
rect 2116 45124 2172 45180
rect 2172 45124 2176 45180
rect 2112 45120 2176 45124
rect 2192 45180 2256 45184
rect 2192 45124 2196 45180
rect 2196 45124 2252 45180
rect 2252 45124 2256 45180
rect 2192 45120 2256 45124
rect 6952 45180 7016 45184
rect 6952 45124 6956 45180
rect 6956 45124 7012 45180
rect 7012 45124 7016 45180
rect 6952 45120 7016 45124
rect 7032 45180 7096 45184
rect 7032 45124 7036 45180
rect 7036 45124 7092 45180
rect 7092 45124 7096 45180
rect 7032 45120 7096 45124
rect 7112 45180 7176 45184
rect 7112 45124 7116 45180
rect 7116 45124 7172 45180
rect 7172 45124 7176 45180
rect 7112 45120 7176 45124
rect 7192 45180 7256 45184
rect 7192 45124 7196 45180
rect 7196 45124 7252 45180
rect 7252 45124 7256 45180
rect 7192 45120 7256 45124
rect 11952 45180 12016 45184
rect 11952 45124 11956 45180
rect 11956 45124 12012 45180
rect 12012 45124 12016 45180
rect 11952 45120 12016 45124
rect 12032 45180 12096 45184
rect 12032 45124 12036 45180
rect 12036 45124 12092 45180
rect 12092 45124 12096 45180
rect 12032 45120 12096 45124
rect 12112 45180 12176 45184
rect 12112 45124 12116 45180
rect 12116 45124 12172 45180
rect 12172 45124 12176 45180
rect 12112 45120 12176 45124
rect 12192 45180 12256 45184
rect 12192 45124 12196 45180
rect 12196 45124 12252 45180
rect 12252 45124 12256 45180
rect 12192 45120 12256 45124
rect 16952 45180 17016 45184
rect 16952 45124 16956 45180
rect 16956 45124 17012 45180
rect 17012 45124 17016 45180
rect 16952 45120 17016 45124
rect 17032 45180 17096 45184
rect 17032 45124 17036 45180
rect 17036 45124 17092 45180
rect 17092 45124 17096 45180
rect 17032 45120 17096 45124
rect 17112 45180 17176 45184
rect 17112 45124 17116 45180
rect 17116 45124 17172 45180
rect 17172 45124 17176 45180
rect 17112 45120 17176 45124
rect 17192 45180 17256 45184
rect 17192 45124 17196 45180
rect 17196 45124 17252 45180
rect 17252 45124 17256 45180
rect 17192 45120 17256 45124
rect 21952 45180 22016 45184
rect 21952 45124 21956 45180
rect 21956 45124 22012 45180
rect 22012 45124 22016 45180
rect 21952 45120 22016 45124
rect 22032 45180 22096 45184
rect 22032 45124 22036 45180
rect 22036 45124 22092 45180
rect 22092 45124 22096 45180
rect 22032 45120 22096 45124
rect 22112 45180 22176 45184
rect 22112 45124 22116 45180
rect 22116 45124 22172 45180
rect 22172 45124 22176 45180
rect 22112 45120 22176 45124
rect 22192 45180 22256 45184
rect 22192 45124 22196 45180
rect 22196 45124 22252 45180
rect 22252 45124 22256 45180
rect 22192 45120 22256 45124
rect 26952 45180 27016 45184
rect 26952 45124 26956 45180
rect 26956 45124 27012 45180
rect 27012 45124 27016 45180
rect 26952 45120 27016 45124
rect 27032 45180 27096 45184
rect 27032 45124 27036 45180
rect 27036 45124 27092 45180
rect 27092 45124 27096 45180
rect 27032 45120 27096 45124
rect 27112 45180 27176 45184
rect 27112 45124 27116 45180
rect 27116 45124 27172 45180
rect 27172 45124 27176 45180
rect 27112 45120 27176 45124
rect 27192 45180 27256 45184
rect 27192 45124 27196 45180
rect 27196 45124 27252 45180
rect 27252 45124 27256 45180
rect 27192 45120 27256 45124
rect 31952 45180 32016 45184
rect 31952 45124 31956 45180
rect 31956 45124 32012 45180
rect 32012 45124 32016 45180
rect 31952 45120 32016 45124
rect 32032 45180 32096 45184
rect 32032 45124 32036 45180
rect 32036 45124 32092 45180
rect 32092 45124 32096 45180
rect 32032 45120 32096 45124
rect 32112 45180 32176 45184
rect 32112 45124 32116 45180
rect 32116 45124 32172 45180
rect 32172 45124 32176 45180
rect 32112 45120 32176 45124
rect 32192 45180 32256 45184
rect 32192 45124 32196 45180
rect 32196 45124 32252 45180
rect 32252 45124 32256 45180
rect 32192 45120 32256 45124
rect 36952 45180 37016 45184
rect 36952 45124 36956 45180
rect 36956 45124 37012 45180
rect 37012 45124 37016 45180
rect 36952 45120 37016 45124
rect 37032 45180 37096 45184
rect 37032 45124 37036 45180
rect 37036 45124 37092 45180
rect 37092 45124 37096 45180
rect 37032 45120 37096 45124
rect 37112 45180 37176 45184
rect 37112 45124 37116 45180
rect 37116 45124 37172 45180
rect 37172 45124 37176 45180
rect 37112 45120 37176 45124
rect 37192 45180 37256 45184
rect 37192 45124 37196 45180
rect 37196 45124 37252 45180
rect 37252 45124 37256 45180
rect 37192 45120 37256 45124
rect 2612 44636 2676 44640
rect 2612 44580 2616 44636
rect 2616 44580 2672 44636
rect 2672 44580 2676 44636
rect 2612 44576 2676 44580
rect 2692 44636 2756 44640
rect 2692 44580 2696 44636
rect 2696 44580 2752 44636
rect 2752 44580 2756 44636
rect 2692 44576 2756 44580
rect 2772 44636 2836 44640
rect 2772 44580 2776 44636
rect 2776 44580 2832 44636
rect 2832 44580 2836 44636
rect 2772 44576 2836 44580
rect 2852 44636 2916 44640
rect 2852 44580 2856 44636
rect 2856 44580 2912 44636
rect 2912 44580 2916 44636
rect 2852 44576 2916 44580
rect 7612 44636 7676 44640
rect 7612 44580 7616 44636
rect 7616 44580 7672 44636
rect 7672 44580 7676 44636
rect 7612 44576 7676 44580
rect 7692 44636 7756 44640
rect 7692 44580 7696 44636
rect 7696 44580 7752 44636
rect 7752 44580 7756 44636
rect 7692 44576 7756 44580
rect 7772 44636 7836 44640
rect 7772 44580 7776 44636
rect 7776 44580 7832 44636
rect 7832 44580 7836 44636
rect 7772 44576 7836 44580
rect 7852 44636 7916 44640
rect 7852 44580 7856 44636
rect 7856 44580 7912 44636
rect 7912 44580 7916 44636
rect 7852 44576 7916 44580
rect 12612 44636 12676 44640
rect 12612 44580 12616 44636
rect 12616 44580 12672 44636
rect 12672 44580 12676 44636
rect 12612 44576 12676 44580
rect 12692 44636 12756 44640
rect 12692 44580 12696 44636
rect 12696 44580 12752 44636
rect 12752 44580 12756 44636
rect 12692 44576 12756 44580
rect 12772 44636 12836 44640
rect 12772 44580 12776 44636
rect 12776 44580 12832 44636
rect 12832 44580 12836 44636
rect 12772 44576 12836 44580
rect 12852 44636 12916 44640
rect 12852 44580 12856 44636
rect 12856 44580 12912 44636
rect 12912 44580 12916 44636
rect 12852 44576 12916 44580
rect 17612 44636 17676 44640
rect 17612 44580 17616 44636
rect 17616 44580 17672 44636
rect 17672 44580 17676 44636
rect 17612 44576 17676 44580
rect 17692 44636 17756 44640
rect 17692 44580 17696 44636
rect 17696 44580 17752 44636
rect 17752 44580 17756 44636
rect 17692 44576 17756 44580
rect 17772 44636 17836 44640
rect 17772 44580 17776 44636
rect 17776 44580 17832 44636
rect 17832 44580 17836 44636
rect 17772 44576 17836 44580
rect 17852 44636 17916 44640
rect 17852 44580 17856 44636
rect 17856 44580 17912 44636
rect 17912 44580 17916 44636
rect 17852 44576 17916 44580
rect 22612 44636 22676 44640
rect 22612 44580 22616 44636
rect 22616 44580 22672 44636
rect 22672 44580 22676 44636
rect 22612 44576 22676 44580
rect 22692 44636 22756 44640
rect 22692 44580 22696 44636
rect 22696 44580 22752 44636
rect 22752 44580 22756 44636
rect 22692 44576 22756 44580
rect 22772 44636 22836 44640
rect 22772 44580 22776 44636
rect 22776 44580 22832 44636
rect 22832 44580 22836 44636
rect 22772 44576 22836 44580
rect 22852 44636 22916 44640
rect 22852 44580 22856 44636
rect 22856 44580 22912 44636
rect 22912 44580 22916 44636
rect 22852 44576 22916 44580
rect 27612 44636 27676 44640
rect 27612 44580 27616 44636
rect 27616 44580 27672 44636
rect 27672 44580 27676 44636
rect 27612 44576 27676 44580
rect 27692 44636 27756 44640
rect 27692 44580 27696 44636
rect 27696 44580 27752 44636
rect 27752 44580 27756 44636
rect 27692 44576 27756 44580
rect 27772 44636 27836 44640
rect 27772 44580 27776 44636
rect 27776 44580 27832 44636
rect 27832 44580 27836 44636
rect 27772 44576 27836 44580
rect 27852 44636 27916 44640
rect 27852 44580 27856 44636
rect 27856 44580 27912 44636
rect 27912 44580 27916 44636
rect 27852 44576 27916 44580
rect 32612 44636 32676 44640
rect 32612 44580 32616 44636
rect 32616 44580 32672 44636
rect 32672 44580 32676 44636
rect 32612 44576 32676 44580
rect 32692 44636 32756 44640
rect 32692 44580 32696 44636
rect 32696 44580 32752 44636
rect 32752 44580 32756 44636
rect 32692 44576 32756 44580
rect 32772 44636 32836 44640
rect 32772 44580 32776 44636
rect 32776 44580 32832 44636
rect 32832 44580 32836 44636
rect 32772 44576 32836 44580
rect 32852 44636 32916 44640
rect 32852 44580 32856 44636
rect 32856 44580 32912 44636
rect 32912 44580 32916 44636
rect 32852 44576 32916 44580
rect 37612 44636 37676 44640
rect 37612 44580 37616 44636
rect 37616 44580 37672 44636
rect 37672 44580 37676 44636
rect 37612 44576 37676 44580
rect 37692 44636 37756 44640
rect 37692 44580 37696 44636
rect 37696 44580 37752 44636
rect 37752 44580 37756 44636
rect 37692 44576 37756 44580
rect 37772 44636 37836 44640
rect 37772 44580 37776 44636
rect 37776 44580 37832 44636
rect 37832 44580 37836 44636
rect 37772 44576 37836 44580
rect 37852 44636 37916 44640
rect 37852 44580 37856 44636
rect 37856 44580 37912 44636
rect 37912 44580 37916 44636
rect 37852 44576 37916 44580
rect 1952 44092 2016 44096
rect 1952 44036 1956 44092
rect 1956 44036 2012 44092
rect 2012 44036 2016 44092
rect 1952 44032 2016 44036
rect 2032 44092 2096 44096
rect 2032 44036 2036 44092
rect 2036 44036 2092 44092
rect 2092 44036 2096 44092
rect 2032 44032 2096 44036
rect 2112 44092 2176 44096
rect 2112 44036 2116 44092
rect 2116 44036 2172 44092
rect 2172 44036 2176 44092
rect 2112 44032 2176 44036
rect 2192 44092 2256 44096
rect 2192 44036 2196 44092
rect 2196 44036 2252 44092
rect 2252 44036 2256 44092
rect 2192 44032 2256 44036
rect 6952 44092 7016 44096
rect 6952 44036 6956 44092
rect 6956 44036 7012 44092
rect 7012 44036 7016 44092
rect 6952 44032 7016 44036
rect 7032 44092 7096 44096
rect 7032 44036 7036 44092
rect 7036 44036 7092 44092
rect 7092 44036 7096 44092
rect 7032 44032 7096 44036
rect 7112 44092 7176 44096
rect 7112 44036 7116 44092
rect 7116 44036 7172 44092
rect 7172 44036 7176 44092
rect 7112 44032 7176 44036
rect 7192 44092 7256 44096
rect 7192 44036 7196 44092
rect 7196 44036 7252 44092
rect 7252 44036 7256 44092
rect 7192 44032 7256 44036
rect 11952 44092 12016 44096
rect 11952 44036 11956 44092
rect 11956 44036 12012 44092
rect 12012 44036 12016 44092
rect 11952 44032 12016 44036
rect 12032 44092 12096 44096
rect 12032 44036 12036 44092
rect 12036 44036 12092 44092
rect 12092 44036 12096 44092
rect 12032 44032 12096 44036
rect 12112 44092 12176 44096
rect 12112 44036 12116 44092
rect 12116 44036 12172 44092
rect 12172 44036 12176 44092
rect 12112 44032 12176 44036
rect 12192 44092 12256 44096
rect 12192 44036 12196 44092
rect 12196 44036 12252 44092
rect 12252 44036 12256 44092
rect 12192 44032 12256 44036
rect 16952 44092 17016 44096
rect 16952 44036 16956 44092
rect 16956 44036 17012 44092
rect 17012 44036 17016 44092
rect 16952 44032 17016 44036
rect 17032 44092 17096 44096
rect 17032 44036 17036 44092
rect 17036 44036 17092 44092
rect 17092 44036 17096 44092
rect 17032 44032 17096 44036
rect 17112 44092 17176 44096
rect 17112 44036 17116 44092
rect 17116 44036 17172 44092
rect 17172 44036 17176 44092
rect 17112 44032 17176 44036
rect 17192 44092 17256 44096
rect 17192 44036 17196 44092
rect 17196 44036 17252 44092
rect 17252 44036 17256 44092
rect 17192 44032 17256 44036
rect 21952 44092 22016 44096
rect 21952 44036 21956 44092
rect 21956 44036 22012 44092
rect 22012 44036 22016 44092
rect 21952 44032 22016 44036
rect 22032 44092 22096 44096
rect 22032 44036 22036 44092
rect 22036 44036 22092 44092
rect 22092 44036 22096 44092
rect 22032 44032 22096 44036
rect 22112 44092 22176 44096
rect 22112 44036 22116 44092
rect 22116 44036 22172 44092
rect 22172 44036 22176 44092
rect 22112 44032 22176 44036
rect 22192 44092 22256 44096
rect 22192 44036 22196 44092
rect 22196 44036 22252 44092
rect 22252 44036 22256 44092
rect 22192 44032 22256 44036
rect 26952 44092 27016 44096
rect 26952 44036 26956 44092
rect 26956 44036 27012 44092
rect 27012 44036 27016 44092
rect 26952 44032 27016 44036
rect 27032 44092 27096 44096
rect 27032 44036 27036 44092
rect 27036 44036 27092 44092
rect 27092 44036 27096 44092
rect 27032 44032 27096 44036
rect 27112 44092 27176 44096
rect 27112 44036 27116 44092
rect 27116 44036 27172 44092
rect 27172 44036 27176 44092
rect 27112 44032 27176 44036
rect 27192 44092 27256 44096
rect 27192 44036 27196 44092
rect 27196 44036 27252 44092
rect 27252 44036 27256 44092
rect 27192 44032 27256 44036
rect 31952 44092 32016 44096
rect 31952 44036 31956 44092
rect 31956 44036 32012 44092
rect 32012 44036 32016 44092
rect 31952 44032 32016 44036
rect 32032 44092 32096 44096
rect 32032 44036 32036 44092
rect 32036 44036 32092 44092
rect 32092 44036 32096 44092
rect 32032 44032 32096 44036
rect 32112 44092 32176 44096
rect 32112 44036 32116 44092
rect 32116 44036 32172 44092
rect 32172 44036 32176 44092
rect 32112 44032 32176 44036
rect 32192 44092 32256 44096
rect 32192 44036 32196 44092
rect 32196 44036 32252 44092
rect 32252 44036 32256 44092
rect 32192 44032 32256 44036
rect 36952 44092 37016 44096
rect 36952 44036 36956 44092
rect 36956 44036 37012 44092
rect 37012 44036 37016 44092
rect 36952 44032 37016 44036
rect 37032 44092 37096 44096
rect 37032 44036 37036 44092
rect 37036 44036 37092 44092
rect 37092 44036 37096 44092
rect 37032 44032 37096 44036
rect 37112 44092 37176 44096
rect 37112 44036 37116 44092
rect 37116 44036 37172 44092
rect 37172 44036 37176 44092
rect 37112 44032 37176 44036
rect 37192 44092 37256 44096
rect 37192 44036 37196 44092
rect 37196 44036 37252 44092
rect 37252 44036 37256 44092
rect 37192 44032 37256 44036
rect 2612 43548 2676 43552
rect 2612 43492 2616 43548
rect 2616 43492 2672 43548
rect 2672 43492 2676 43548
rect 2612 43488 2676 43492
rect 2692 43548 2756 43552
rect 2692 43492 2696 43548
rect 2696 43492 2752 43548
rect 2752 43492 2756 43548
rect 2692 43488 2756 43492
rect 2772 43548 2836 43552
rect 2772 43492 2776 43548
rect 2776 43492 2832 43548
rect 2832 43492 2836 43548
rect 2772 43488 2836 43492
rect 2852 43548 2916 43552
rect 2852 43492 2856 43548
rect 2856 43492 2912 43548
rect 2912 43492 2916 43548
rect 2852 43488 2916 43492
rect 7612 43548 7676 43552
rect 7612 43492 7616 43548
rect 7616 43492 7672 43548
rect 7672 43492 7676 43548
rect 7612 43488 7676 43492
rect 7692 43548 7756 43552
rect 7692 43492 7696 43548
rect 7696 43492 7752 43548
rect 7752 43492 7756 43548
rect 7692 43488 7756 43492
rect 7772 43548 7836 43552
rect 7772 43492 7776 43548
rect 7776 43492 7832 43548
rect 7832 43492 7836 43548
rect 7772 43488 7836 43492
rect 7852 43548 7916 43552
rect 7852 43492 7856 43548
rect 7856 43492 7912 43548
rect 7912 43492 7916 43548
rect 7852 43488 7916 43492
rect 12612 43548 12676 43552
rect 12612 43492 12616 43548
rect 12616 43492 12672 43548
rect 12672 43492 12676 43548
rect 12612 43488 12676 43492
rect 12692 43548 12756 43552
rect 12692 43492 12696 43548
rect 12696 43492 12752 43548
rect 12752 43492 12756 43548
rect 12692 43488 12756 43492
rect 12772 43548 12836 43552
rect 12772 43492 12776 43548
rect 12776 43492 12832 43548
rect 12832 43492 12836 43548
rect 12772 43488 12836 43492
rect 12852 43548 12916 43552
rect 12852 43492 12856 43548
rect 12856 43492 12912 43548
rect 12912 43492 12916 43548
rect 12852 43488 12916 43492
rect 17612 43548 17676 43552
rect 17612 43492 17616 43548
rect 17616 43492 17672 43548
rect 17672 43492 17676 43548
rect 17612 43488 17676 43492
rect 17692 43548 17756 43552
rect 17692 43492 17696 43548
rect 17696 43492 17752 43548
rect 17752 43492 17756 43548
rect 17692 43488 17756 43492
rect 17772 43548 17836 43552
rect 17772 43492 17776 43548
rect 17776 43492 17832 43548
rect 17832 43492 17836 43548
rect 17772 43488 17836 43492
rect 17852 43548 17916 43552
rect 17852 43492 17856 43548
rect 17856 43492 17912 43548
rect 17912 43492 17916 43548
rect 17852 43488 17916 43492
rect 22612 43548 22676 43552
rect 22612 43492 22616 43548
rect 22616 43492 22672 43548
rect 22672 43492 22676 43548
rect 22612 43488 22676 43492
rect 22692 43548 22756 43552
rect 22692 43492 22696 43548
rect 22696 43492 22752 43548
rect 22752 43492 22756 43548
rect 22692 43488 22756 43492
rect 22772 43548 22836 43552
rect 22772 43492 22776 43548
rect 22776 43492 22832 43548
rect 22832 43492 22836 43548
rect 22772 43488 22836 43492
rect 22852 43548 22916 43552
rect 22852 43492 22856 43548
rect 22856 43492 22912 43548
rect 22912 43492 22916 43548
rect 22852 43488 22916 43492
rect 27612 43548 27676 43552
rect 27612 43492 27616 43548
rect 27616 43492 27672 43548
rect 27672 43492 27676 43548
rect 27612 43488 27676 43492
rect 27692 43548 27756 43552
rect 27692 43492 27696 43548
rect 27696 43492 27752 43548
rect 27752 43492 27756 43548
rect 27692 43488 27756 43492
rect 27772 43548 27836 43552
rect 27772 43492 27776 43548
rect 27776 43492 27832 43548
rect 27832 43492 27836 43548
rect 27772 43488 27836 43492
rect 27852 43548 27916 43552
rect 27852 43492 27856 43548
rect 27856 43492 27912 43548
rect 27912 43492 27916 43548
rect 27852 43488 27916 43492
rect 32612 43548 32676 43552
rect 32612 43492 32616 43548
rect 32616 43492 32672 43548
rect 32672 43492 32676 43548
rect 32612 43488 32676 43492
rect 32692 43548 32756 43552
rect 32692 43492 32696 43548
rect 32696 43492 32752 43548
rect 32752 43492 32756 43548
rect 32692 43488 32756 43492
rect 32772 43548 32836 43552
rect 32772 43492 32776 43548
rect 32776 43492 32832 43548
rect 32832 43492 32836 43548
rect 32772 43488 32836 43492
rect 32852 43548 32916 43552
rect 32852 43492 32856 43548
rect 32856 43492 32912 43548
rect 32912 43492 32916 43548
rect 32852 43488 32916 43492
rect 37612 43548 37676 43552
rect 37612 43492 37616 43548
rect 37616 43492 37672 43548
rect 37672 43492 37676 43548
rect 37612 43488 37676 43492
rect 37692 43548 37756 43552
rect 37692 43492 37696 43548
rect 37696 43492 37752 43548
rect 37752 43492 37756 43548
rect 37692 43488 37756 43492
rect 37772 43548 37836 43552
rect 37772 43492 37776 43548
rect 37776 43492 37832 43548
rect 37832 43492 37836 43548
rect 37772 43488 37836 43492
rect 37852 43548 37916 43552
rect 37852 43492 37856 43548
rect 37856 43492 37912 43548
rect 37912 43492 37916 43548
rect 37852 43488 37916 43492
rect 1952 43004 2016 43008
rect 1952 42948 1956 43004
rect 1956 42948 2012 43004
rect 2012 42948 2016 43004
rect 1952 42944 2016 42948
rect 2032 43004 2096 43008
rect 2032 42948 2036 43004
rect 2036 42948 2092 43004
rect 2092 42948 2096 43004
rect 2032 42944 2096 42948
rect 2112 43004 2176 43008
rect 2112 42948 2116 43004
rect 2116 42948 2172 43004
rect 2172 42948 2176 43004
rect 2112 42944 2176 42948
rect 2192 43004 2256 43008
rect 2192 42948 2196 43004
rect 2196 42948 2252 43004
rect 2252 42948 2256 43004
rect 2192 42944 2256 42948
rect 6952 43004 7016 43008
rect 6952 42948 6956 43004
rect 6956 42948 7012 43004
rect 7012 42948 7016 43004
rect 6952 42944 7016 42948
rect 7032 43004 7096 43008
rect 7032 42948 7036 43004
rect 7036 42948 7092 43004
rect 7092 42948 7096 43004
rect 7032 42944 7096 42948
rect 7112 43004 7176 43008
rect 7112 42948 7116 43004
rect 7116 42948 7172 43004
rect 7172 42948 7176 43004
rect 7112 42944 7176 42948
rect 7192 43004 7256 43008
rect 7192 42948 7196 43004
rect 7196 42948 7252 43004
rect 7252 42948 7256 43004
rect 7192 42944 7256 42948
rect 11952 43004 12016 43008
rect 11952 42948 11956 43004
rect 11956 42948 12012 43004
rect 12012 42948 12016 43004
rect 11952 42944 12016 42948
rect 12032 43004 12096 43008
rect 12032 42948 12036 43004
rect 12036 42948 12092 43004
rect 12092 42948 12096 43004
rect 12032 42944 12096 42948
rect 12112 43004 12176 43008
rect 12112 42948 12116 43004
rect 12116 42948 12172 43004
rect 12172 42948 12176 43004
rect 12112 42944 12176 42948
rect 12192 43004 12256 43008
rect 12192 42948 12196 43004
rect 12196 42948 12252 43004
rect 12252 42948 12256 43004
rect 12192 42944 12256 42948
rect 16952 43004 17016 43008
rect 16952 42948 16956 43004
rect 16956 42948 17012 43004
rect 17012 42948 17016 43004
rect 16952 42944 17016 42948
rect 17032 43004 17096 43008
rect 17032 42948 17036 43004
rect 17036 42948 17092 43004
rect 17092 42948 17096 43004
rect 17032 42944 17096 42948
rect 17112 43004 17176 43008
rect 17112 42948 17116 43004
rect 17116 42948 17172 43004
rect 17172 42948 17176 43004
rect 17112 42944 17176 42948
rect 17192 43004 17256 43008
rect 17192 42948 17196 43004
rect 17196 42948 17252 43004
rect 17252 42948 17256 43004
rect 17192 42944 17256 42948
rect 21952 43004 22016 43008
rect 21952 42948 21956 43004
rect 21956 42948 22012 43004
rect 22012 42948 22016 43004
rect 21952 42944 22016 42948
rect 22032 43004 22096 43008
rect 22032 42948 22036 43004
rect 22036 42948 22092 43004
rect 22092 42948 22096 43004
rect 22032 42944 22096 42948
rect 22112 43004 22176 43008
rect 22112 42948 22116 43004
rect 22116 42948 22172 43004
rect 22172 42948 22176 43004
rect 22112 42944 22176 42948
rect 22192 43004 22256 43008
rect 22192 42948 22196 43004
rect 22196 42948 22252 43004
rect 22252 42948 22256 43004
rect 22192 42944 22256 42948
rect 26952 43004 27016 43008
rect 26952 42948 26956 43004
rect 26956 42948 27012 43004
rect 27012 42948 27016 43004
rect 26952 42944 27016 42948
rect 27032 43004 27096 43008
rect 27032 42948 27036 43004
rect 27036 42948 27092 43004
rect 27092 42948 27096 43004
rect 27032 42944 27096 42948
rect 27112 43004 27176 43008
rect 27112 42948 27116 43004
rect 27116 42948 27172 43004
rect 27172 42948 27176 43004
rect 27112 42944 27176 42948
rect 27192 43004 27256 43008
rect 27192 42948 27196 43004
rect 27196 42948 27252 43004
rect 27252 42948 27256 43004
rect 27192 42944 27256 42948
rect 31952 43004 32016 43008
rect 31952 42948 31956 43004
rect 31956 42948 32012 43004
rect 32012 42948 32016 43004
rect 31952 42944 32016 42948
rect 32032 43004 32096 43008
rect 32032 42948 32036 43004
rect 32036 42948 32092 43004
rect 32092 42948 32096 43004
rect 32032 42944 32096 42948
rect 32112 43004 32176 43008
rect 32112 42948 32116 43004
rect 32116 42948 32172 43004
rect 32172 42948 32176 43004
rect 32112 42944 32176 42948
rect 32192 43004 32256 43008
rect 32192 42948 32196 43004
rect 32196 42948 32252 43004
rect 32252 42948 32256 43004
rect 32192 42944 32256 42948
rect 36952 43004 37016 43008
rect 36952 42948 36956 43004
rect 36956 42948 37012 43004
rect 37012 42948 37016 43004
rect 36952 42944 37016 42948
rect 37032 43004 37096 43008
rect 37032 42948 37036 43004
rect 37036 42948 37092 43004
rect 37092 42948 37096 43004
rect 37032 42944 37096 42948
rect 37112 43004 37176 43008
rect 37112 42948 37116 43004
rect 37116 42948 37172 43004
rect 37172 42948 37176 43004
rect 37112 42944 37176 42948
rect 37192 43004 37256 43008
rect 37192 42948 37196 43004
rect 37196 42948 37252 43004
rect 37252 42948 37256 43004
rect 37192 42944 37256 42948
rect 2612 42460 2676 42464
rect 2612 42404 2616 42460
rect 2616 42404 2672 42460
rect 2672 42404 2676 42460
rect 2612 42400 2676 42404
rect 2692 42460 2756 42464
rect 2692 42404 2696 42460
rect 2696 42404 2752 42460
rect 2752 42404 2756 42460
rect 2692 42400 2756 42404
rect 2772 42460 2836 42464
rect 2772 42404 2776 42460
rect 2776 42404 2832 42460
rect 2832 42404 2836 42460
rect 2772 42400 2836 42404
rect 2852 42460 2916 42464
rect 2852 42404 2856 42460
rect 2856 42404 2912 42460
rect 2912 42404 2916 42460
rect 2852 42400 2916 42404
rect 7612 42460 7676 42464
rect 7612 42404 7616 42460
rect 7616 42404 7672 42460
rect 7672 42404 7676 42460
rect 7612 42400 7676 42404
rect 7692 42460 7756 42464
rect 7692 42404 7696 42460
rect 7696 42404 7752 42460
rect 7752 42404 7756 42460
rect 7692 42400 7756 42404
rect 7772 42460 7836 42464
rect 7772 42404 7776 42460
rect 7776 42404 7832 42460
rect 7832 42404 7836 42460
rect 7772 42400 7836 42404
rect 7852 42460 7916 42464
rect 7852 42404 7856 42460
rect 7856 42404 7912 42460
rect 7912 42404 7916 42460
rect 7852 42400 7916 42404
rect 12612 42460 12676 42464
rect 12612 42404 12616 42460
rect 12616 42404 12672 42460
rect 12672 42404 12676 42460
rect 12612 42400 12676 42404
rect 12692 42460 12756 42464
rect 12692 42404 12696 42460
rect 12696 42404 12752 42460
rect 12752 42404 12756 42460
rect 12692 42400 12756 42404
rect 12772 42460 12836 42464
rect 12772 42404 12776 42460
rect 12776 42404 12832 42460
rect 12832 42404 12836 42460
rect 12772 42400 12836 42404
rect 12852 42460 12916 42464
rect 12852 42404 12856 42460
rect 12856 42404 12912 42460
rect 12912 42404 12916 42460
rect 12852 42400 12916 42404
rect 17612 42460 17676 42464
rect 17612 42404 17616 42460
rect 17616 42404 17672 42460
rect 17672 42404 17676 42460
rect 17612 42400 17676 42404
rect 17692 42460 17756 42464
rect 17692 42404 17696 42460
rect 17696 42404 17752 42460
rect 17752 42404 17756 42460
rect 17692 42400 17756 42404
rect 17772 42460 17836 42464
rect 17772 42404 17776 42460
rect 17776 42404 17832 42460
rect 17832 42404 17836 42460
rect 17772 42400 17836 42404
rect 17852 42460 17916 42464
rect 17852 42404 17856 42460
rect 17856 42404 17912 42460
rect 17912 42404 17916 42460
rect 17852 42400 17916 42404
rect 22612 42460 22676 42464
rect 22612 42404 22616 42460
rect 22616 42404 22672 42460
rect 22672 42404 22676 42460
rect 22612 42400 22676 42404
rect 22692 42460 22756 42464
rect 22692 42404 22696 42460
rect 22696 42404 22752 42460
rect 22752 42404 22756 42460
rect 22692 42400 22756 42404
rect 22772 42460 22836 42464
rect 22772 42404 22776 42460
rect 22776 42404 22832 42460
rect 22832 42404 22836 42460
rect 22772 42400 22836 42404
rect 22852 42460 22916 42464
rect 22852 42404 22856 42460
rect 22856 42404 22912 42460
rect 22912 42404 22916 42460
rect 22852 42400 22916 42404
rect 27612 42460 27676 42464
rect 27612 42404 27616 42460
rect 27616 42404 27672 42460
rect 27672 42404 27676 42460
rect 27612 42400 27676 42404
rect 27692 42460 27756 42464
rect 27692 42404 27696 42460
rect 27696 42404 27752 42460
rect 27752 42404 27756 42460
rect 27692 42400 27756 42404
rect 27772 42460 27836 42464
rect 27772 42404 27776 42460
rect 27776 42404 27832 42460
rect 27832 42404 27836 42460
rect 27772 42400 27836 42404
rect 27852 42460 27916 42464
rect 27852 42404 27856 42460
rect 27856 42404 27912 42460
rect 27912 42404 27916 42460
rect 27852 42400 27916 42404
rect 32612 42460 32676 42464
rect 32612 42404 32616 42460
rect 32616 42404 32672 42460
rect 32672 42404 32676 42460
rect 32612 42400 32676 42404
rect 32692 42460 32756 42464
rect 32692 42404 32696 42460
rect 32696 42404 32752 42460
rect 32752 42404 32756 42460
rect 32692 42400 32756 42404
rect 32772 42460 32836 42464
rect 32772 42404 32776 42460
rect 32776 42404 32832 42460
rect 32832 42404 32836 42460
rect 32772 42400 32836 42404
rect 32852 42460 32916 42464
rect 32852 42404 32856 42460
rect 32856 42404 32912 42460
rect 32912 42404 32916 42460
rect 32852 42400 32916 42404
rect 37612 42460 37676 42464
rect 37612 42404 37616 42460
rect 37616 42404 37672 42460
rect 37672 42404 37676 42460
rect 37612 42400 37676 42404
rect 37692 42460 37756 42464
rect 37692 42404 37696 42460
rect 37696 42404 37752 42460
rect 37752 42404 37756 42460
rect 37692 42400 37756 42404
rect 37772 42460 37836 42464
rect 37772 42404 37776 42460
rect 37776 42404 37832 42460
rect 37832 42404 37836 42460
rect 37772 42400 37836 42404
rect 37852 42460 37916 42464
rect 37852 42404 37856 42460
rect 37856 42404 37912 42460
rect 37912 42404 37916 42460
rect 37852 42400 37916 42404
rect 1952 41916 2016 41920
rect 1952 41860 1956 41916
rect 1956 41860 2012 41916
rect 2012 41860 2016 41916
rect 1952 41856 2016 41860
rect 2032 41916 2096 41920
rect 2032 41860 2036 41916
rect 2036 41860 2092 41916
rect 2092 41860 2096 41916
rect 2032 41856 2096 41860
rect 2112 41916 2176 41920
rect 2112 41860 2116 41916
rect 2116 41860 2172 41916
rect 2172 41860 2176 41916
rect 2112 41856 2176 41860
rect 2192 41916 2256 41920
rect 2192 41860 2196 41916
rect 2196 41860 2252 41916
rect 2252 41860 2256 41916
rect 2192 41856 2256 41860
rect 6952 41916 7016 41920
rect 6952 41860 6956 41916
rect 6956 41860 7012 41916
rect 7012 41860 7016 41916
rect 6952 41856 7016 41860
rect 7032 41916 7096 41920
rect 7032 41860 7036 41916
rect 7036 41860 7092 41916
rect 7092 41860 7096 41916
rect 7032 41856 7096 41860
rect 7112 41916 7176 41920
rect 7112 41860 7116 41916
rect 7116 41860 7172 41916
rect 7172 41860 7176 41916
rect 7112 41856 7176 41860
rect 7192 41916 7256 41920
rect 7192 41860 7196 41916
rect 7196 41860 7252 41916
rect 7252 41860 7256 41916
rect 7192 41856 7256 41860
rect 11952 41916 12016 41920
rect 11952 41860 11956 41916
rect 11956 41860 12012 41916
rect 12012 41860 12016 41916
rect 11952 41856 12016 41860
rect 12032 41916 12096 41920
rect 12032 41860 12036 41916
rect 12036 41860 12092 41916
rect 12092 41860 12096 41916
rect 12032 41856 12096 41860
rect 12112 41916 12176 41920
rect 12112 41860 12116 41916
rect 12116 41860 12172 41916
rect 12172 41860 12176 41916
rect 12112 41856 12176 41860
rect 12192 41916 12256 41920
rect 12192 41860 12196 41916
rect 12196 41860 12252 41916
rect 12252 41860 12256 41916
rect 12192 41856 12256 41860
rect 16952 41916 17016 41920
rect 16952 41860 16956 41916
rect 16956 41860 17012 41916
rect 17012 41860 17016 41916
rect 16952 41856 17016 41860
rect 17032 41916 17096 41920
rect 17032 41860 17036 41916
rect 17036 41860 17092 41916
rect 17092 41860 17096 41916
rect 17032 41856 17096 41860
rect 17112 41916 17176 41920
rect 17112 41860 17116 41916
rect 17116 41860 17172 41916
rect 17172 41860 17176 41916
rect 17112 41856 17176 41860
rect 17192 41916 17256 41920
rect 17192 41860 17196 41916
rect 17196 41860 17252 41916
rect 17252 41860 17256 41916
rect 17192 41856 17256 41860
rect 21952 41916 22016 41920
rect 21952 41860 21956 41916
rect 21956 41860 22012 41916
rect 22012 41860 22016 41916
rect 21952 41856 22016 41860
rect 22032 41916 22096 41920
rect 22032 41860 22036 41916
rect 22036 41860 22092 41916
rect 22092 41860 22096 41916
rect 22032 41856 22096 41860
rect 22112 41916 22176 41920
rect 22112 41860 22116 41916
rect 22116 41860 22172 41916
rect 22172 41860 22176 41916
rect 22112 41856 22176 41860
rect 22192 41916 22256 41920
rect 22192 41860 22196 41916
rect 22196 41860 22252 41916
rect 22252 41860 22256 41916
rect 22192 41856 22256 41860
rect 26952 41916 27016 41920
rect 26952 41860 26956 41916
rect 26956 41860 27012 41916
rect 27012 41860 27016 41916
rect 26952 41856 27016 41860
rect 27032 41916 27096 41920
rect 27032 41860 27036 41916
rect 27036 41860 27092 41916
rect 27092 41860 27096 41916
rect 27032 41856 27096 41860
rect 27112 41916 27176 41920
rect 27112 41860 27116 41916
rect 27116 41860 27172 41916
rect 27172 41860 27176 41916
rect 27112 41856 27176 41860
rect 27192 41916 27256 41920
rect 27192 41860 27196 41916
rect 27196 41860 27252 41916
rect 27252 41860 27256 41916
rect 27192 41856 27256 41860
rect 31952 41916 32016 41920
rect 31952 41860 31956 41916
rect 31956 41860 32012 41916
rect 32012 41860 32016 41916
rect 31952 41856 32016 41860
rect 32032 41916 32096 41920
rect 32032 41860 32036 41916
rect 32036 41860 32092 41916
rect 32092 41860 32096 41916
rect 32032 41856 32096 41860
rect 32112 41916 32176 41920
rect 32112 41860 32116 41916
rect 32116 41860 32172 41916
rect 32172 41860 32176 41916
rect 32112 41856 32176 41860
rect 32192 41916 32256 41920
rect 32192 41860 32196 41916
rect 32196 41860 32252 41916
rect 32252 41860 32256 41916
rect 32192 41856 32256 41860
rect 36952 41916 37016 41920
rect 36952 41860 36956 41916
rect 36956 41860 37012 41916
rect 37012 41860 37016 41916
rect 36952 41856 37016 41860
rect 37032 41916 37096 41920
rect 37032 41860 37036 41916
rect 37036 41860 37092 41916
rect 37092 41860 37096 41916
rect 37032 41856 37096 41860
rect 37112 41916 37176 41920
rect 37112 41860 37116 41916
rect 37116 41860 37172 41916
rect 37172 41860 37176 41916
rect 37112 41856 37176 41860
rect 37192 41916 37256 41920
rect 37192 41860 37196 41916
rect 37196 41860 37252 41916
rect 37252 41860 37256 41916
rect 37192 41856 37256 41860
rect 2612 41372 2676 41376
rect 2612 41316 2616 41372
rect 2616 41316 2672 41372
rect 2672 41316 2676 41372
rect 2612 41312 2676 41316
rect 2692 41372 2756 41376
rect 2692 41316 2696 41372
rect 2696 41316 2752 41372
rect 2752 41316 2756 41372
rect 2692 41312 2756 41316
rect 2772 41372 2836 41376
rect 2772 41316 2776 41372
rect 2776 41316 2832 41372
rect 2832 41316 2836 41372
rect 2772 41312 2836 41316
rect 2852 41372 2916 41376
rect 2852 41316 2856 41372
rect 2856 41316 2912 41372
rect 2912 41316 2916 41372
rect 2852 41312 2916 41316
rect 7612 41372 7676 41376
rect 7612 41316 7616 41372
rect 7616 41316 7672 41372
rect 7672 41316 7676 41372
rect 7612 41312 7676 41316
rect 7692 41372 7756 41376
rect 7692 41316 7696 41372
rect 7696 41316 7752 41372
rect 7752 41316 7756 41372
rect 7692 41312 7756 41316
rect 7772 41372 7836 41376
rect 7772 41316 7776 41372
rect 7776 41316 7832 41372
rect 7832 41316 7836 41372
rect 7772 41312 7836 41316
rect 7852 41372 7916 41376
rect 7852 41316 7856 41372
rect 7856 41316 7912 41372
rect 7912 41316 7916 41372
rect 7852 41312 7916 41316
rect 12612 41372 12676 41376
rect 12612 41316 12616 41372
rect 12616 41316 12672 41372
rect 12672 41316 12676 41372
rect 12612 41312 12676 41316
rect 12692 41372 12756 41376
rect 12692 41316 12696 41372
rect 12696 41316 12752 41372
rect 12752 41316 12756 41372
rect 12692 41312 12756 41316
rect 12772 41372 12836 41376
rect 12772 41316 12776 41372
rect 12776 41316 12832 41372
rect 12832 41316 12836 41372
rect 12772 41312 12836 41316
rect 12852 41372 12916 41376
rect 12852 41316 12856 41372
rect 12856 41316 12912 41372
rect 12912 41316 12916 41372
rect 12852 41312 12916 41316
rect 17612 41372 17676 41376
rect 17612 41316 17616 41372
rect 17616 41316 17672 41372
rect 17672 41316 17676 41372
rect 17612 41312 17676 41316
rect 17692 41372 17756 41376
rect 17692 41316 17696 41372
rect 17696 41316 17752 41372
rect 17752 41316 17756 41372
rect 17692 41312 17756 41316
rect 17772 41372 17836 41376
rect 17772 41316 17776 41372
rect 17776 41316 17832 41372
rect 17832 41316 17836 41372
rect 17772 41312 17836 41316
rect 17852 41372 17916 41376
rect 17852 41316 17856 41372
rect 17856 41316 17912 41372
rect 17912 41316 17916 41372
rect 17852 41312 17916 41316
rect 22612 41372 22676 41376
rect 22612 41316 22616 41372
rect 22616 41316 22672 41372
rect 22672 41316 22676 41372
rect 22612 41312 22676 41316
rect 22692 41372 22756 41376
rect 22692 41316 22696 41372
rect 22696 41316 22752 41372
rect 22752 41316 22756 41372
rect 22692 41312 22756 41316
rect 22772 41372 22836 41376
rect 22772 41316 22776 41372
rect 22776 41316 22832 41372
rect 22832 41316 22836 41372
rect 22772 41312 22836 41316
rect 22852 41372 22916 41376
rect 22852 41316 22856 41372
rect 22856 41316 22912 41372
rect 22912 41316 22916 41372
rect 22852 41312 22916 41316
rect 27612 41372 27676 41376
rect 27612 41316 27616 41372
rect 27616 41316 27672 41372
rect 27672 41316 27676 41372
rect 27612 41312 27676 41316
rect 27692 41372 27756 41376
rect 27692 41316 27696 41372
rect 27696 41316 27752 41372
rect 27752 41316 27756 41372
rect 27692 41312 27756 41316
rect 27772 41372 27836 41376
rect 27772 41316 27776 41372
rect 27776 41316 27832 41372
rect 27832 41316 27836 41372
rect 27772 41312 27836 41316
rect 27852 41372 27916 41376
rect 27852 41316 27856 41372
rect 27856 41316 27912 41372
rect 27912 41316 27916 41372
rect 27852 41312 27916 41316
rect 32612 41372 32676 41376
rect 32612 41316 32616 41372
rect 32616 41316 32672 41372
rect 32672 41316 32676 41372
rect 32612 41312 32676 41316
rect 32692 41372 32756 41376
rect 32692 41316 32696 41372
rect 32696 41316 32752 41372
rect 32752 41316 32756 41372
rect 32692 41312 32756 41316
rect 32772 41372 32836 41376
rect 32772 41316 32776 41372
rect 32776 41316 32832 41372
rect 32832 41316 32836 41372
rect 32772 41312 32836 41316
rect 32852 41372 32916 41376
rect 32852 41316 32856 41372
rect 32856 41316 32912 41372
rect 32912 41316 32916 41372
rect 32852 41312 32916 41316
rect 37612 41372 37676 41376
rect 37612 41316 37616 41372
rect 37616 41316 37672 41372
rect 37672 41316 37676 41372
rect 37612 41312 37676 41316
rect 37692 41372 37756 41376
rect 37692 41316 37696 41372
rect 37696 41316 37752 41372
rect 37752 41316 37756 41372
rect 37692 41312 37756 41316
rect 37772 41372 37836 41376
rect 37772 41316 37776 41372
rect 37776 41316 37832 41372
rect 37832 41316 37836 41372
rect 37772 41312 37836 41316
rect 37852 41372 37916 41376
rect 37852 41316 37856 41372
rect 37856 41316 37912 41372
rect 37912 41316 37916 41372
rect 37852 41312 37916 41316
rect 1952 40828 2016 40832
rect 1952 40772 1956 40828
rect 1956 40772 2012 40828
rect 2012 40772 2016 40828
rect 1952 40768 2016 40772
rect 2032 40828 2096 40832
rect 2032 40772 2036 40828
rect 2036 40772 2092 40828
rect 2092 40772 2096 40828
rect 2032 40768 2096 40772
rect 2112 40828 2176 40832
rect 2112 40772 2116 40828
rect 2116 40772 2172 40828
rect 2172 40772 2176 40828
rect 2112 40768 2176 40772
rect 2192 40828 2256 40832
rect 2192 40772 2196 40828
rect 2196 40772 2252 40828
rect 2252 40772 2256 40828
rect 2192 40768 2256 40772
rect 6952 40828 7016 40832
rect 6952 40772 6956 40828
rect 6956 40772 7012 40828
rect 7012 40772 7016 40828
rect 6952 40768 7016 40772
rect 7032 40828 7096 40832
rect 7032 40772 7036 40828
rect 7036 40772 7092 40828
rect 7092 40772 7096 40828
rect 7032 40768 7096 40772
rect 7112 40828 7176 40832
rect 7112 40772 7116 40828
rect 7116 40772 7172 40828
rect 7172 40772 7176 40828
rect 7112 40768 7176 40772
rect 7192 40828 7256 40832
rect 7192 40772 7196 40828
rect 7196 40772 7252 40828
rect 7252 40772 7256 40828
rect 7192 40768 7256 40772
rect 11952 40828 12016 40832
rect 11952 40772 11956 40828
rect 11956 40772 12012 40828
rect 12012 40772 12016 40828
rect 11952 40768 12016 40772
rect 12032 40828 12096 40832
rect 12032 40772 12036 40828
rect 12036 40772 12092 40828
rect 12092 40772 12096 40828
rect 12032 40768 12096 40772
rect 12112 40828 12176 40832
rect 12112 40772 12116 40828
rect 12116 40772 12172 40828
rect 12172 40772 12176 40828
rect 12112 40768 12176 40772
rect 12192 40828 12256 40832
rect 12192 40772 12196 40828
rect 12196 40772 12252 40828
rect 12252 40772 12256 40828
rect 12192 40768 12256 40772
rect 16952 40828 17016 40832
rect 16952 40772 16956 40828
rect 16956 40772 17012 40828
rect 17012 40772 17016 40828
rect 16952 40768 17016 40772
rect 17032 40828 17096 40832
rect 17032 40772 17036 40828
rect 17036 40772 17092 40828
rect 17092 40772 17096 40828
rect 17032 40768 17096 40772
rect 17112 40828 17176 40832
rect 17112 40772 17116 40828
rect 17116 40772 17172 40828
rect 17172 40772 17176 40828
rect 17112 40768 17176 40772
rect 17192 40828 17256 40832
rect 17192 40772 17196 40828
rect 17196 40772 17252 40828
rect 17252 40772 17256 40828
rect 17192 40768 17256 40772
rect 21952 40828 22016 40832
rect 21952 40772 21956 40828
rect 21956 40772 22012 40828
rect 22012 40772 22016 40828
rect 21952 40768 22016 40772
rect 22032 40828 22096 40832
rect 22032 40772 22036 40828
rect 22036 40772 22092 40828
rect 22092 40772 22096 40828
rect 22032 40768 22096 40772
rect 22112 40828 22176 40832
rect 22112 40772 22116 40828
rect 22116 40772 22172 40828
rect 22172 40772 22176 40828
rect 22112 40768 22176 40772
rect 22192 40828 22256 40832
rect 22192 40772 22196 40828
rect 22196 40772 22252 40828
rect 22252 40772 22256 40828
rect 22192 40768 22256 40772
rect 26952 40828 27016 40832
rect 26952 40772 26956 40828
rect 26956 40772 27012 40828
rect 27012 40772 27016 40828
rect 26952 40768 27016 40772
rect 27032 40828 27096 40832
rect 27032 40772 27036 40828
rect 27036 40772 27092 40828
rect 27092 40772 27096 40828
rect 27032 40768 27096 40772
rect 27112 40828 27176 40832
rect 27112 40772 27116 40828
rect 27116 40772 27172 40828
rect 27172 40772 27176 40828
rect 27112 40768 27176 40772
rect 27192 40828 27256 40832
rect 27192 40772 27196 40828
rect 27196 40772 27252 40828
rect 27252 40772 27256 40828
rect 27192 40768 27256 40772
rect 31952 40828 32016 40832
rect 31952 40772 31956 40828
rect 31956 40772 32012 40828
rect 32012 40772 32016 40828
rect 31952 40768 32016 40772
rect 32032 40828 32096 40832
rect 32032 40772 32036 40828
rect 32036 40772 32092 40828
rect 32092 40772 32096 40828
rect 32032 40768 32096 40772
rect 32112 40828 32176 40832
rect 32112 40772 32116 40828
rect 32116 40772 32172 40828
rect 32172 40772 32176 40828
rect 32112 40768 32176 40772
rect 32192 40828 32256 40832
rect 32192 40772 32196 40828
rect 32196 40772 32252 40828
rect 32252 40772 32256 40828
rect 32192 40768 32256 40772
rect 36952 40828 37016 40832
rect 36952 40772 36956 40828
rect 36956 40772 37012 40828
rect 37012 40772 37016 40828
rect 36952 40768 37016 40772
rect 37032 40828 37096 40832
rect 37032 40772 37036 40828
rect 37036 40772 37092 40828
rect 37092 40772 37096 40828
rect 37032 40768 37096 40772
rect 37112 40828 37176 40832
rect 37112 40772 37116 40828
rect 37116 40772 37172 40828
rect 37172 40772 37176 40828
rect 37112 40768 37176 40772
rect 37192 40828 37256 40832
rect 37192 40772 37196 40828
rect 37196 40772 37252 40828
rect 37252 40772 37256 40828
rect 37192 40768 37256 40772
rect 23612 40624 23676 40628
rect 23612 40568 23626 40624
rect 23626 40568 23676 40624
rect 23612 40564 23676 40568
rect 2612 40284 2676 40288
rect 2612 40228 2616 40284
rect 2616 40228 2672 40284
rect 2672 40228 2676 40284
rect 2612 40224 2676 40228
rect 2692 40284 2756 40288
rect 2692 40228 2696 40284
rect 2696 40228 2752 40284
rect 2752 40228 2756 40284
rect 2692 40224 2756 40228
rect 2772 40284 2836 40288
rect 2772 40228 2776 40284
rect 2776 40228 2832 40284
rect 2832 40228 2836 40284
rect 2772 40224 2836 40228
rect 2852 40284 2916 40288
rect 2852 40228 2856 40284
rect 2856 40228 2912 40284
rect 2912 40228 2916 40284
rect 2852 40224 2916 40228
rect 7612 40284 7676 40288
rect 7612 40228 7616 40284
rect 7616 40228 7672 40284
rect 7672 40228 7676 40284
rect 7612 40224 7676 40228
rect 7692 40284 7756 40288
rect 7692 40228 7696 40284
rect 7696 40228 7752 40284
rect 7752 40228 7756 40284
rect 7692 40224 7756 40228
rect 7772 40284 7836 40288
rect 7772 40228 7776 40284
rect 7776 40228 7832 40284
rect 7832 40228 7836 40284
rect 7772 40224 7836 40228
rect 7852 40284 7916 40288
rect 7852 40228 7856 40284
rect 7856 40228 7912 40284
rect 7912 40228 7916 40284
rect 7852 40224 7916 40228
rect 12612 40284 12676 40288
rect 12612 40228 12616 40284
rect 12616 40228 12672 40284
rect 12672 40228 12676 40284
rect 12612 40224 12676 40228
rect 12692 40284 12756 40288
rect 12692 40228 12696 40284
rect 12696 40228 12752 40284
rect 12752 40228 12756 40284
rect 12692 40224 12756 40228
rect 12772 40284 12836 40288
rect 12772 40228 12776 40284
rect 12776 40228 12832 40284
rect 12832 40228 12836 40284
rect 12772 40224 12836 40228
rect 12852 40284 12916 40288
rect 12852 40228 12856 40284
rect 12856 40228 12912 40284
rect 12912 40228 12916 40284
rect 12852 40224 12916 40228
rect 17612 40284 17676 40288
rect 17612 40228 17616 40284
rect 17616 40228 17672 40284
rect 17672 40228 17676 40284
rect 17612 40224 17676 40228
rect 17692 40284 17756 40288
rect 17692 40228 17696 40284
rect 17696 40228 17752 40284
rect 17752 40228 17756 40284
rect 17692 40224 17756 40228
rect 17772 40284 17836 40288
rect 17772 40228 17776 40284
rect 17776 40228 17832 40284
rect 17832 40228 17836 40284
rect 17772 40224 17836 40228
rect 17852 40284 17916 40288
rect 17852 40228 17856 40284
rect 17856 40228 17912 40284
rect 17912 40228 17916 40284
rect 17852 40224 17916 40228
rect 22612 40284 22676 40288
rect 22612 40228 22616 40284
rect 22616 40228 22672 40284
rect 22672 40228 22676 40284
rect 22612 40224 22676 40228
rect 22692 40284 22756 40288
rect 22692 40228 22696 40284
rect 22696 40228 22752 40284
rect 22752 40228 22756 40284
rect 22692 40224 22756 40228
rect 22772 40284 22836 40288
rect 22772 40228 22776 40284
rect 22776 40228 22832 40284
rect 22832 40228 22836 40284
rect 22772 40224 22836 40228
rect 22852 40284 22916 40288
rect 22852 40228 22856 40284
rect 22856 40228 22912 40284
rect 22912 40228 22916 40284
rect 22852 40224 22916 40228
rect 27612 40284 27676 40288
rect 27612 40228 27616 40284
rect 27616 40228 27672 40284
rect 27672 40228 27676 40284
rect 27612 40224 27676 40228
rect 27692 40284 27756 40288
rect 27692 40228 27696 40284
rect 27696 40228 27752 40284
rect 27752 40228 27756 40284
rect 27692 40224 27756 40228
rect 27772 40284 27836 40288
rect 27772 40228 27776 40284
rect 27776 40228 27832 40284
rect 27832 40228 27836 40284
rect 27772 40224 27836 40228
rect 27852 40284 27916 40288
rect 27852 40228 27856 40284
rect 27856 40228 27912 40284
rect 27912 40228 27916 40284
rect 27852 40224 27916 40228
rect 32612 40284 32676 40288
rect 32612 40228 32616 40284
rect 32616 40228 32672 40284
rect 32672 40228 32676 40284
rect 32612 40224 32676 40228
rect 32692 40284 32756 40288
rect 32692 40228 32696 40284
rect 32696 40228 32752 40284
rect 32752 40228 32756 40284
rect 32692 40224 32756 40228
rect 32772 40284 32836 40288
rect 32772 40228 32776 40284
rect 32776 40228 32832 40284
rect 32832 40228 32836 40284
rect 32772 40224 32836 40228
rect 32852 40284 32916 40288
rect 32852 40228 32856 40284
rect 32856 40228 32912 40284
rect 32912 40228 32916 40284
rect 32852 40224 32916 40228
rect 37612 40284 37676 40288
rect 37612 40228 37616 40284
rect 37616 40228 37672 40284
rect 37672 40228 37676 40284
rect 37612 40224 37676 40228
rect 37692 40284 37756 40288
rect 37692 40228 37696 40284
rect 37696 40228 37752 40284
rect 37752 40228 37756 40284
rect 37692 40224 37756 40228
rect 37772 40284 37836 40288
rect 37772 40228 37776 40284
rect 37776 40228 37832 40284
rect 37832 40228 37836 40284
rect 37772 40224 37836 40228
rect 37852 40284 37916 40288
rect 37852 40228 37856 40284
rect 37856 40228 37912 40284
rect 37912 40228 37916 40284
rect 37852 40224 37916 40228
rect 30604 40080 30668 40084
rect 30604 40024 30618 40080
rect 30618 40024 30668 40080
rect 30604 40020 30668 40024
rect 1952 39740 2016 39744
rect 1952 39684 1956 39740
rect 1956 39684 2012 39740
rect 2012 39684 2016 39740
rect 1952 39680 2016 39684
rect 2032 39740 2096 39744
rect 2032 39684 2036 39740
rect 2036 39684 2092 39740
rect 2092 39684 2096 39740
rect 2032 39680 2096 39684
rect 2112 39740 2176 39744
rect 2112 39684 2116 39740
rect 2116 39684 2172 39740
rect 2172 39684 2176 39740
rect 2112 39680 2176 39684
rect 2192 39740 2256 39744
rect 2192 39684 2196 39740
rect 2196 39684 2252 39740
rect 2252 39684 2256 39740
rect 2192 39680 2256 39684
rect 6952 39740 7016 39744
rect 6952 39684 6956 39740
rect 6956 39684 7012 39740
rect 7012 39684 7016 39740
rect 6952 39680 7016 39684
rect 7032 39740 7096 39744
rect 7032 39684 7036 39740
rect 7036 39684 7092 39740
rect 7092 39684 7096 39740
rect 7032 39680 7096 39684
rect 7112 39740 7176 39744
rect 7112 39684 7116 39740
rect 7116 39684 7172 39740
rect 7172 39684 7176 39740
rect 7112 39680 7176 39684
rect 7192 39740 7256 39744
rect 7192 39684 7196 39740
rect 7196 39684 7252 39740
rect 7252 39684 7256 39740
rect 7192 39680 7256 39684
rect 11952 39740 12016 39744
rect 11952 39684 11956 39740
rect 11956 39684 12012 39740
rect 12012 39684 12016 39740
rect 11952 39680 12016 39684
rect 12032 39740 12096 39744
rect 12032 39684 12036 39740
rect 12036 39684 12092 39740
rect 12092 39684 12096 39740
rect 12032 39680 12096 39684
rect 12112 39740 12176 39744
rect 12112 39684 12116 39740
rect 12116 39684 12172 39740
rect 12172 39684 12176 39740
rect 12112 39680 12176 39684
rect 12192 39740 12256 39744
rect 12192 39684 12196 39740
rect 12196 39684 12252 39740
rect 12252 39684 12256 39740
rect 12192 39680 12256 39684
rect 16952 39740 17016 39744
rect 16952 39684 16956 39740
rect 16956 39684 17012 39740
rect 17012 39684 17016 39740
rect 16952 39680 17016 39684
rect 17032 39740 17096 39744
rect 17032 39684 17036 39740
rect 17036 39684 17092 39740
rect 17092 39684 17096 39740
rect 17032 39680 17096 39684
rect 17112 39740 17176 39744
rect 17112 39684 17116 39740
rect 17116 39684 17172 39740
rect 17172 39684 17176 39740
rect 17112 39680 17176 39684
rect 17192 39740 17256 39744
rect 17192 39684 17196 39740
rect 17196 39684 17252 39740
rect 17252 39684 17256 39740
rect 17192 39680 17256 39684
rect 21952 39740 22016 39744
rect 21952 39684 21956 39740
rect 21956 39684 22012 39740
rect 22012 39684 22016 39740
rect 21952 39680 22016 39684
rect 22032 39740 22096 39744
rect 22032 39684 22036 39740
rect 22036 39684 22092 39740
rect 22092 39684 22096 39740
rect 22032 39680 22096 39684
rect 22112 39740 22176 39744
rect 22112 39684 22116 39740
rect 22116 39684 22172 39740
rect 22172 39684 22176 39740
rect 22112 39680 22176 39684
rect 22192 39740 22256 39744
rect 22192 39684 22196 39740
rect 22196 39684 22252 39740
rect 22252 39684 22256 39740
rect 22192 39680 22256 39684
rect 26952 39740 27016 39744
rect 26952 39684 26956 39740
rect 26956 39684 27012 39740
rect 27012 39684 27016 39740
rect 26952 39680 27016 39684
rect 27032 39740 27096 39744
rect 27032 39684 27036 39740
rect 27036 39684 27092 39740
rect 27092 39684 27096 39740
rect 27032 39680 27096 39684
rect 27112 39740 27176 39744
rect 27112 39684 27116 39740
rect 27116 39684 27172 39740
rect 27172 39684 27176 39740
rect 27112 39680 27176 39684
rect 27192 39740 27256 39744
rect 27192 39684 27196 39740
rect 27196 39684 27252 39740
rect 27252 39684 27256 39740
rect 27192 39680 27256 39684
rect 31952 39740 32016 39744
rect 31952 39684 31956 39740
rect 31956 39684 32012 39740
rect 32012 39684 32016 39740
rect 31952 39680 32016 39684
rect 32032 39740 32096 39744
rect 32032 39684 32036 39740
rect 32036 39684 32092 39740
rect 32092 39684 32096 39740
rect 32032 39680 32096 39684
rect 32112 39740 32176 39744
rect 32112 39684 32116 39740
rect 32116 39684 32172 39740
rect 32172 39684 32176 39740
rect 32112 39680 32176 39684
rect 32192 39740 32256 39744
rect 32192 39684 32196 39740
rect 32196 39684 32252 39740
rect 32252 39684 32256 39740
rect 32192 39680 32256 39684
rect 36952 39740 37016 39744
rect 36952 39684 36956 39740
rect 36956 39684 37012 39740
rect 37012 39684 37016 39740
rect 36952 39680 37016 39684
rect 37032 39740 37096 39744
rect 37032 39684 37036 39740
rect 37036 39684 37092 39740
rect 37092 39684 37096 39740
rect 37032 39680 37096 39684
rect 37112 39740 37176 39744
rect 37112 39684 37116 39740
rect 37116 39684 37172 39740
rect 37172 39684 37176 39740
rect 37112 39680 37176 39684
rect 37192 39740 37256 39744
rect 37192 39684 37196 39740
rect 37196 39684 37252 39740
rect 37252 39684 37256 39740
rect 37192 39680 37256 39684
rect 2612 39196 2676 39200
rect 2612 39140 2616 39196
rect 2616 39140 2672 39196
rect 2672 39140 2676 39196
rect 2612 39136 2676 39140
rect 2692 39196 2756 39200
rect 2692 39140 2696 39196
rect 2696 39140 2752 39196
rect 2752 39140 2756 39196
rect 2692 39136 2756 39140
rect 2772 39196 2836 39200
rect 2772 39140 2776 39196
rect 2776 39140 2832 39196
rect 2832 39140 2836 39196
rect 2772 39136 2836 39140
rect 2852 39196 2916 39200
rect 2852 39140 2856 39196
rect 2856 39140 2912 39196
rect 2912 39140 2916 39196
rect 2852 39136 2916 39140
rect 7612 39196 7676 39200
rect 7612 39140 7616 39196
rect 7616 39140 7672 39196
rect 7672 39140 7676 39196
rect 7612 39136 7676 39140
rect 7692 39196 7756 39200
rect 7692 39140 7696 39196
rect 7696 39140 7752 39196
rect 7752 39140 7756 39196
rect 7692 39136 7756 39140
rect 7772 39196 7836 39200
rect 7772 39140 7776 39196
rect 7776 39140 7832 39196
rect 7832 39140 7836 39196
rect 7772 39136 7836 39140
rect 7852 39196 7916 39200
rect 7852 39140 7856 39196
rect 7856 39140 7912 39196
rect 7912 39140 7916 39196
rect 7852 39136 7916 39140
rect 12612 39196 12676 39200
rect 12612 39140 12616 39196
rect 12616 39140 12672 39196
rect 12672 39140 12676 39196
rect 12612 39136 12676 39140
rect 12692 39196 12756 39200
rect 12692 39140 12696 39196
rect 12696 39140 12752 39196
rect 12752 39140 12756 39196
rect 12692 39136 12756 39140
rect 12772 39196 12836 39200
rect 12772 39140 12776 39196
rect 12776 39140 12832 39196
rect 12832 39140 12836 39196
rect 12772 39136 12836 39140
rect 12852 39196 12916 39200
rect 12852 39140 12856 39196
rect 12856 39140 12912 39196
rect 12912 39140 12916 39196
rect 12852 39136 12916 39140
rect 17612 39196 17676 39200
rect 17612 39140 17616 39196
rect 17616 39140 17672 39196
rect 17672 39140 17676 39196
rect 17612 39136 17676 39140
rect 17692 39196 17756 39200
rect 17692 39140 17696 39196
rect 17696 39140 17752 39196
rect 17752 39140 17756 39196
rect 17692 39136 17756 39140
rect 17772 39196 17836 39200
rect 17772 39140 17776 39196
rect 17776 39140 17832 39196
rect 17832 39140 17836 39196
rect 17772 39136 17836 39140
rect 17852 39196 17916 39200
rect 17852 39140 17856 39196
rect 17856 39140 17912 39196
rect 17912 39140 17916 39196
rect 17852 39136 17916 39140
rect 22612 39196 22676 39200
rect 22612 39140 22616 39196
rect 22616 39140 22672 39196
rect 22672 39140 22676 39196
rect 22612 39136 22676 39140
rect 22692 39196 22756 39200
rect 22692 39140 22696 39196
rect 22696 39140 22752 39196
rect 22752 39140 22756 39196
rect 22692 39136 22756 39140
rect 22772 39196 22836 39200
rect 22772 39140 22776 39196
rect 22776 39140 22832 39196
rect 22832 39140 22836 39196
rect 22772 39136 22836 39140
rect 22852 39196 22916 39200
rect 22852 39140 22856 39196
rect 22856 39140 22912 39196
rect 22912 39140 22916 39196
rect 22852 39136 22916 39140
rect 27612 39196 27676 39200
rect 27612 39140 27616 39196
rect 27616 39140 27672 39196
rect 27672 39140 27676 39196
rect 27612 39136 27676 39140
rect 27692 39196 27756 39200
rect 27692 39140 27696 39196
rect 27696 39140 27752 39196
rect 27752 39140 27756 39196
rect 27692 39136 27756 39140
rect 27772 39196 27836 39200
rect 27772 39140 27776 39196
rect 27776 39140 27832 39196
rect 27832 39140 27836 39196
rect 27772 39136 27836 39140
rect 27852 39196 27916 39200
rect 27852 39140 27856 39196
rect 27856 39140 27912 39196
rect 27912 39140 27916 39196
rect 27852 39136 27916 39140
rect 32612 39196 32676 39200
rect 32612 39140 32616 39196
rect 32616 39140 32672 39196
rect 32672 39140 32676 39196
rect 32612 39136 32676 39140
rect 32692 39196 32756 39200
rect 32692 39140 32696 39196
rect 32696 39140 32752 39196
rect 32752 39140 32756 39196
rect 32692 39136 32756 39140
rect 32772 39196 32836 39200
rect 32772 39140 32776 39196
rect 32776 39140 32832 39196
rect 32832 39140 32836 39196
rect 32772 39136 32836 39140
rect 32852 39196 32916 39200
rect 32852 39140 32856 39196
rect 32856 39140 32912 39196
rect 32912 39140 32916 39196
rect 32852 39136 32916 39140
rect 37612 39196 37676 39200
rect 37612 39140 37616 39196
rect 37616 39140 37672 39196
rect 37672 39140 37676 39196
rect 37612 39136 37676 39140
rect 37692 39196 37756 39200
rect 37692 39140 37696 39196
rect 37696 39140 37752 39196
rect 37752 39140 37756 39196
rect 37692 39136 37756 39140
rect 37772 39196 37836 39200
rect 37772 39140 37776 39196
rect 37776 39140 37832 39196
rect 37832 39140 37836 39196
rect 37772 39136 37836 39140
rect 37852 39196 37916 39200
rect 37852 39140 37856 39196
rect 37856 39140 37912 39196
rect 37912 39140 37916 39196
rect 37852 39136 37916 39140
rect 23244 38660 23308 38724
rect 1952 38652 2016 38656
rect 1952 38596 1956 38652
rect 1956 38596 2012 38652
rect 2012 38596 2016 38652
rect 1952 38592 2016 38596
rect 2032 38652 2096 38656
rect 2032 38596 2036 38652
rect 2036 38596 2092 38652
rect 2092 38596 2096 38652
rect 2032 38592 2096 38596
rect 2112 38652 2176 38656
rect 2112 38596 2116 38652
rect 2116 38596 2172 38652
rect 2172 38596 2176 38652
rect 2112 38592 2176 38596
rect 2192 38652 2256 38656
rect 2192 38596 2196 38652
rect 2196 38596 2252 38652
rect 2252 38596 2256 38652
rect 2192 38592 2256 38596
rect 6952 38652 7016 38656
rect 6952 38596 6956 38652
rect 6956 38596 7012 38652
rect 7012 38596 7016 38652
rect 6952 38592 7016 38596
rect 7032 38652 7096 38656
rect 7032 38596 7036 38652
rect 7036 38596 7092 38652
rect 7092 38596 7096 38652
rect 7032 38592 7096 38596
rect 7112 38652 7176 38656
rect 7112 38596 7116 38652
rect 7116 38596 7172 38652
rect 7172 38596 7176 38652
rect 7112 38592 7176 38596
rect 7192 38652 7256 38656
rect 7192 38596 7196 38652
rect 7196 38596 7252 38652
rect 7252 38596 7256 38652
rect 7192 38592 7256 38596
rect 11952 38652 12016 38656
rect 11952 38596 11956 38652
rect 11956 38596 12012 38652
rect 12012 38596 12016 38652
rect 11952 38592 12016 38596
rect 12032 38652 12096 38656
rect 12032 38596 12036 38652
rect 12036 38596 12092 38652
rect 12092 38596 12096 38652
rect 12032 38592 12096 38596
rect 12112 38652 12176 38656
rect 12112 38596 12116 38652
rect 12116 38596 12172 38652
rect 12172 38596 12176 38652
rect 12112 38592 12176 38596
rect 12192 38652 12256 38656
rect 12192 38596 12196 38652
rect 12196 38596 12252 38652
rect 12252 38596 12256 38652
rect 12192 38592 12256 38596
rect 16952 38652 17016 38656
rect 16952 38596 16956 38652
rect 16956 38596 17012 38652
rect 17012 38596 17016 38652
rect 16952 38592 17016 38596
rect 17032 38652 17096 38656
rect 17032 38596 17036 38652
rect 17036 38596 17092 38652
rect 17092 38596 17096 38652
rect 17032 38592 17096 38596
rect 17112 38652 17176 38656
rect 17112 38596 17116 38652
rect 17116 38596 17172 38652
rect 17172 38596 17176 38652
rect 17112 38592 17176 38596
rect 17192 38652 17256 38656
rect 17192 38596 17196 38652
rect 17196 38596 17252 38652
rect 17252 38596 17256 38652
rect 17192 38592 17256 38596
rect 21952 38652 22016 38656
rect 21952 38596 21956 38652
rect 21956 38596 22012 38652
rect 22012 38596 22016 38652
rect 21952 38592 22016 38596
rect 22032 38652 22096 38656
rect 22032 38596 22036 38652
rect 22036 38596 22092 38652
rect 22092 38596 22096 38652
rect 22032 38592 22096 38596
rect 22112 38652 22176 38656
rect 22112 38596 22116 38652
rect 22116 38596 22172 38652
rect 22172 38596 22176 38652
rect 22112 38592 22176 38596
rect 22192 38652 22256 38656
rect 22192 38596 22196 38652
rect 22196 38596 22252 38652
rect 22252 38596 22256 38652
rect 22192 38592 22256 38596
rect 26952 38652 27016 38656
rect 26952 38596 26956 38652
rect 26956 38596 27012 38652
rect 27012 38596 27016 38652
rect 26952 38592 27016 38596
rect 27032 38652 27096 38656
rect 27032 38596 27036 38652
rect 27036 38596 27092 38652
rect 27092 38596 27096 38652
rect 27032 38592 27096 38596
rect 27112 38652 27176 38656
rect 27112 38596 27116 38652
rect 27116 38596 27172 38652
rect 27172 38596 27176 38652
rect 27112 38592 27176 38596
rect 27192 38652 27256 38656
rect 27192 38596 27196 38652
rect 27196 38596 27252 38652
rect 27252 38596 27256 38652
rect 27192 38592 27256 38596
rect 31952 38652 32016 38656
rect 31952 38596 31956 38652
rect 31956 38596 32012 38652
rect 32012 38596 32016 38652
rect 31952 38592 32016 38596
rect 32032 38652 32096 38656
rect 32032 38596 32036 38652
rect 32036 38596 32092 38652
rect 32092 38596 32096 38652
rect 32032 38592 32096 38596
rect 32112 38652 32176 38656
rect 32112 38596 32116 38652
rect 32116 38596 32172 38652
rect 32172 38596 32176 38652
rect 32112 38592 32176 38596
rect 32192 38652 32256 38656
rect 32192 38596 32196 38652
rect 32196 38596 32252 38652
rect 32252 38596 32256 38652
rect 32192 38592 32256 38596
rect 36952 38652 37016 38656
rect 36952 38596 36956 38652
rect 36956 38596 37012 38652
rect 37012 38596 37016 38652
rect 36952 38592 37016 38596
rect 37032 38652 37096 38656
rect 37032 38596 37036 38652
rect 37036 38596 37092 38652
rect 37092 38596 37096 38652
rect 37032 38592 37096 38596
rect 37112 38652 37176 38656
rect 37112 38596 37116 38652
rect 37116 38596 37172 38652
rect 37172 38596 37176 38652
rect 37112 38592 37176 38596
rect 37192 38652 37256 38656
rect 37192 38596 37196 38652
rect 37196 38596 37252 38652
rect 37252 38596 37256 38652
rect 37192 38592 37256 38596
rect 24716 38448 24780 38452
rect 24716 38392 24766 38448
rect 24766 38392 24780 38448
rect 24716 38388 24780 38392
rect 2612 38108 2676 38112
rect 2612 38052 2616 38108
rect 2616 38052 2672 38108
rect 2672 38052 2676 38108
rect 2612 38048 2676 38052
rect 2692 38108 2756 38112
rect 2692 38052 2696 38108
rect 2696 38052 2752 38108
rect 2752 38052 2756 38108
rect 2692 38048 2756 38052
rect 2772 38108 2836 38112
rect 2772 38052 2776 38108
rect 2776 38052 2832 38108
rect 2832 38052 2836 38108
rect 2772 38048 2836 38052
rect 2852 38108 2916 38112
rect 2852 38052 2856 38108
rect 2856 38052 2912 38108
rect 2912 38052 2916 38108
rect 2852 38048 2916 38052
rect 7612 38108 7676 38112
rect 7612 38052 7616 38108
rect 7616 38052 7672 38108
rect 7672 38052 7676 38108
rect 7612 38048 7676 38052
rect 7692 38108 7756 38112
rect 7692 38052 7696 38108
rect 7696 38052 7752 38108
rect 7752 38052 7756 38108
rect 7692 38048 7756 38052
rect 7772 38108 7836 38112
rect 7772 38052 7776 38108
rect 7776 38052 7832 38108
rect 7832 38052 7836 38108
rect 7772 38048 7836 38052
rect 7852 38108 7916 38112
rect 7852 38052 7856 38108
rect 7856 38052 7912 38108
rect 7912 38052 7916 38108
rect 7852 38048 7916 38052
rect 12612 38108 12676 38112
rect 12612 38052 12616 38108
rect 12616 38052 12672 38108
rect 12672 38052 12676 38108
rect 12612 38048 12676 38052
rect 12692 38108 12756 38112
rect 12692 38052 12696 38108
rect 12696 38052 12752 38108
rect 12752 38052 12756 38108
rect 12692 38048 12756 38052
rect 12772 38108 12836 38112
rect 12772 38052 12776 38108
rect 12776 38052 12832 38108
rect 12832 38052 12836 38108
rect 12772 38048 12836 38052
rect 12852 38108 12916 38112
rect 12852 38052 12856 38108
rect 12856 38052 12912 38108
rect 12912 38052 12916 38108
rect 12852 38048 12916 38052
rect 17612 38108 17676 38112
rect 17612 38052 17616 38108
rect 17616 38052 17672 38108
rect 17672 38052 17676 38108
rect 17612 38048 17676 38052
rect 17692 38108 17756 38112
rect 17692 38052 17696 38108
rect 17696 38052 17752 38108
rect 17752 38052 17756 38108
rect 17692 38048 17756 38052
rect 17772 38108 17836 38112
rect 17772 38052 17776 38108
rect 17776 38052 17832 38108
rect 17832 38052 17836 38108
rect 17772 38048 17836 38052
rect 17852 38108 17916 38112
rect 17852 38052 17856 38108
rect 17856 38052 17912 38108
rect 17912 38052 17916 38108
rect 17852 38048 17916 38052
rect 22612 38108 22676 38112
rect 22612 38052 22616 38108
rect 22616 38052 22672 38108
rect 22672 38052 22676 38108
rect 22612 38048 22676 38052
rect 22692 38108 22756 38112
rect 22692 38052 22696 38108
rect 22696 38052 22752 38108
rect 22752 38052 22756 38108
rect 22692 38048 22756 38052
rect 22772 38108 22836 38112
rect 22772 38052 22776 38108
rect 22776 38052 22832 38108
rect 22832 38052 22836 38108
rect 22772 38048 22836 38052
rect 22852 38108 22916 38112
rect 22852 38052 22856 38108
rect 22856 38052 22912 38108
rect 22912 38052 22916 38108
rect 22852 38048 22916 38052
rect 27612 38108 27676 38112
rect 27612 38052 27616 38108
rect 27616 38052 27672 38108
rect 27672 38052 27676 38108
rect 27612 38048 27676 38052
rect 27692 38108 27756 38112
rect 27692 38052 27696 38108
rect 27696 38052 27752 38108
rect 27752 38052 27756 38108
rect 27692 38048 27756 38052
rect 27772 38108 27836 38112
rect 27772 38052 27776 38108
rect 27776 38052 27832 38108
rect 27832 38052 27836 38108
rect 27772 38048 27836 38052
rect 27852 38108 27916 38112
rect 27852 38052 27856 38108
rect 27856 38052 27912 38108
rect 27912 38052 27916 38108
rect 27852 38048 27916 38052
rect 32612 38108 32676 38112
rect 32612 38052 32616 38108
rect 32616 38052 32672 38108
rect 32672 38052 32676 38108
rect 32612 38048 32676 38052
rect 32692 38108 32756 38112
rect 32692 38052 32696 38108
rect 32696 38052 32752 38108
rect 32752 38052 32756 38108
rect 32692 38048 32756 38052
rect 32772 38108 32836 38112
rect 32772 38052 32776 38108
rect 32776 38052 32832 38108
rect 32832 38052 32836 38108
rect 32772 38048 32836 38052
rect 32852 38108 32916 38112
rect 32852 38052 32856 38108
rect 32856 38052 32912 38108
rect 32912 38052 32916 38108
rect 32852 38048 32916 38052
rect 37612 38108 37676 38112
rect 37612 38052 37616 38108
rect 37616 38052 37672 38108
rect 37672 38052 37676 38108
rect 37612 38048 37676 38052
rect 37692 38108 37756 38112
rect 37692 38052 37696 38108
rect 37696 38052 37752 38108
rect 37752 38052 37756 38108
rect 37692 38048 37756 38052
rect 37772 38108 37836 38112
rect 37772 38052 37776 38108
rect 37776 38052 37832 38108
rect 37832 38052 37836 38108
rect 37772 38048 37836 38052
rect 37852 38108 37916 38112
rect 37852 38052 37856 38108
rect 37856 38052 37912 38108
rect 37912 38052 37916 38108
rect 37852 38048 37916 38052
rect 25268 38040 25332 38044
rect 25268 37984 25282 38040
rect 25282 37984 25332 38040
rect 25268 37980 25332 37984
rect 1952 37564 2016 37568
rect 1952 37508 1956 37564
rect 1956 37508 2012 37564
rect 2012 37508 2016 37564
rect 1952 37504 2016 37508
rect 2032 37564 2096 37568
rect 2032 37508 2036 37564
rect 2036 37508 2092 37564
rect 2092 37508 2096 37564
rect 2032 37504 2096 37508
rect 2112 37564 2176 37568
rect 2112 37508 2116 37564
rect 2116 37508 2172 37564
rect 2172 37508 2176 37564
rect 2112 37504 2176 37508
rect 2192 37564 2256 37568
rect 2192 37508 2196 37564
rect 2196 37508 2252 37564
rect 2252 37508 2256 37564
rect 2192 37504 2256 37508
rect 6952 37564 7016 37568
rect 6952 37508 6956 37564
rect 6956 37508 7012 37564
rect 7012 37508 7016 37564
rect 6952 37504 7016 37508
rect 7032 37564 7096 37568
rect 7032 37508 7036 37564
rect 7036 37508 7092 37564
rect 7092 37508 7096 37564
rect 7032 37504 7096 37508
rect 7112 37564 7176 37568
rect 7112 37508 7116 37564
rect 7116 37508 7172 37564
rect 7172 37508 7176 37564
rect 7112 37504 7176 37508
rect 7192 37564 7256 37568
rect 7192 37508 7196 37564
rect 7196 37508 7252 37564
rect 7252 37508 7256 37564
rect 7192 37504 7256 37508
rect 11952 37564 12016 37568
rect 11952 37508 11956 37564
rect 11956 37508 12012 37564
rect 12012 37508 12016 37564
rect 11952 37504 12016 37508
rect 12032 37564 12096 37568
rect 12032 37508 12036 37564
rect 12036 37508 12092 37564
rect 12092 37508 12096 37564
rect 12032 37504 12096 37508
rect 12112 37564 12176 37568
rect 12112 37508 12116 37564
rect 12116 37508 12172 37564
rect 12172 37508 12176 37564
rect 12112 37504 12176 37508
rect 12192 37564 12256 37568
rect 12192 37508 12196 37564
rect 12196 37508 12252 37564
rect 12252 37508 12256 37564
rect 12192 37504 12256 37508
rect 16952 37564 17016 37568
rect 16952 37508 16956 37564
rect 16956 37508 17012 37564
rect 17012 37508 17016 37564
rect 16952 37504 17016 37508
rect 17032 37564 17096 37568
rect 17032 37508 17036 37564
rect 17036 37508 17092 37564
rect 17092 37508 17096 37564
rect 17032 37504 17096 37508
rect 17112 37564 17176 37568
rect 17112 37508 17116 37564
rect 17116 37508 17172 37564
rect 17172 37508 17176 37564
rect 17112 37504 17176 37508
rect 17192 37564 17256 37568
rect 17192 37508 17196 37564
rect 17196 37508 17252 37564
rect 17252 37508 17256 37564
rect 17192 37504 17256 37508
rect 21952 37564 22016 37568
rect 21952 37508 21956 37564
rect 21956 37508 22012 37564
rect 22012 37508 22016 37564
rect 21952 37504 22016 37508
rect 22032 37564 22096 37568
rect 22032 37508 22036 37564
rect 22036 37508 22092 37564
rect 22092 37508 22096 37564
rect 22032 37504 22096 37508
rect 22112 37564 22176 37568
rect 22112 37508 22116 37564
rect 22116 37508 22172 37564
rect 22172 37508 22176 37564
rect 22112 37504 22176 37508
rect 22192 37564 22256 37568
rect 22192 37508 22196 37564
rect 22196 37508 22252 37564
rect 22252 37508 22256 37564
rect 22192 37504 22256 37508
rect 26952 37564 27016 37568
rect 26952 37508 26956 37564
rect 26956 37508 27012 37564
rect 27012 37508 27016 37564
rect 26952 37504 27016 37508
rect 27032 37564 27096 37568
rect 27032 37508 27036 37564
rect 27036 37508 27092 37564
rect 27092 37508 27096 37564
rect 27032 37504 27096 37508
rect 27112 37564 27176 37568
rect 27112 37508 27116 37564
rect 27116 37508 27172 37564
rect 27172 37508 27176 37564
rect 27112 37504 27176 37508
rect 27192 37564 27256 37568
rect 27192 37508 27196 37564
rect 27196 37508 27252 37564
rect 27252 37508 27256 37564
rect 27192 37504 27256 37508
rect 31952 37564 32016 37568
rect 31952 37508 31956 37564
rect 31956 37508 32012 37564
rect 32012 37508 32016 37564
rect 31952 37504 32016 37508
rect 32032 37564 32096 37568
rect 32032 37508 32036 37564
rect 32036 37508 32092 37564
rect 32092 37508 32096 37564
rect 32032 37504 32096 37508
rect 32112 37564 32176 37568
rect 32112 37508 32116 37564
rect 32116 37508 32172 37564
rect 32172 37508 32176 37564
rect 32112 37504 32176 37508
rect 32192 37564 32256 37568
rect 32192 37508 32196 37564
rect 32196 37508 32252 37564
rect 32252 37508 32256 37564
rect 32192 37504 32256 37508
rect 36952 37564 37016 37568
rect 36952 37508 36956 37564
rect 36956 37508 37012 37564
rect 37012 37508 37016 37564
rect 36952 37504 37016 37508
rect 37032 37564 37096 37568
rect 37032 37508 37036 37564
rect 37036 37508 37092 37564
rect 37092 37508 37096 37564
rect 37032 37504 37096 37508
rect 37112 37564 37176 37568
rect 37112 37508 37116 37564
rect 37116 37508 37172 37564
rect 37172 37508 37176 37564
rect 37112 37504 37176 37508
rect 37192 37564 37256 37568
rect 37192 37508 37196 37564
rect 37196 37508 37252 37564
rect 37252 37508 37256 37564
rect 37192 37504 37256 37508
rect 2612 37020 2676 37024
rect 2612 36964 2616 37020
rect 2616 36964 2672 37020
rect 2672 36964 2676 37020
rect 2612 36960 2676 36964
rect 2692 37020 2756 37024
rect 2692 36964 2696 37020
rect 2696 36964 2752 37020
rect 2752 36964 2756 37020
rect 2692 36960 2756 36964
rect 2772 37020 2836 37024
rect 2772 36964 2776 37020
rect 2776 36964 2832 37020
rect 2832 36964 2836 37020
rect 2772 36960 2836 36964
rect 2852 37020 2916 37024
rect 2852 36964 2856 37020
rect 2856 36964 2912 37020
rect 2912 36964 2916 37020
rect 2852 36960 2916 36964
rect 7612 37020 7676 37024
rect 7612 36964 7616 37020
rect 7616 36964 7672 37020
rect 7672 36964 7676 37020
rect 7612 36960 7676 36964
rect 7692 37020 7756 37024
rect 7692 36964 7696 37020
rect 7696 36964 7752 37020
rect 7752 36964 7756 37020
rect 7692 36960 7756 36964
rect 7772 37020 7836 37024
rect 7772 36964 7776 37020
rect 7776 36964 7832 37020
rect 7832 36964 7836 37020
rect 7772 36960 7836 36964
rect 7852 37020 7916 37024
rect 7852 36964 7856 37020
rect 7856 36964 7912 37020
rect 7912 36964 7916 37020
rect 7852 36960 7916 36964
rect 12612 37020 12676 37024
rect 12612 36964 12616 37020
rect 12616 36964 12672 37020
rect 12672 36964 12676 37020
rect 12612 36960 12676 36964
rect 12692 37020 12756 37024
rect 12692 36964 12696 37020
rect 12696 36964 12752 37020
rect 12752 36964 12756 37020
rect 12692 36960 12756 36964
rect 12772 37020 12836 37024
rect 12772 36964 12776 37020
rect 12776 36964 12832 37020
rect 12832 36964 12836 37020
rect 12772 36960 12836 36964
rect 12852 37020 12916 37024
rect 12852 36964 12856 37020
rect 12856 36964 12912 37020
rect 12912 36964 12916 37020
rect 12852 36960 12916 36964
rect 17612 37020 17676 37024
rect 17612 36964 17616 37020
rect 17616 36964 17672 37020
rect 17672 36964 17676 37020
rect 17612 36960 17676 36964
rect 17692 37020 17756 37024
rect 17692 36964 17696 37020
rect 17696 36964 17752 37020
rect 17752 36964 17756 37020
rect 17692 36960 17756 36964
rect 17772 37020 17836 37024
rect 17772 36964 17776 37020
rect 17776 36964 17832 37020
rect 17832 36964 17836 37020
rect 17772 36960 17836 36964
rect 17852 37020 17916 37024
rect 17852 36964 17856 37020
rect 17856 36964 17912 37020
rect 17912 36964 17916 37020
rect 17852 36960 17916 36964
rect 22612 37020 22676 37024
rect 22612 36964 22616 37020
rect 22616 36964 22672 37020
rect 22672 36964 22676 37020
rect 22612 36960 22676 36964
rect 22692 37020 22756 37024
rect 22692 36964 22696 37020
rect 22696 36964 22752 37020
rect 22752 36964 22756 37020
rect 22692 36960 22756 36964
rect 22772 37020 22836 37024
rect 22772 36964 22776 37020
rect 22776 36964 22832 37020
rect 22832 36964 22836 37020
rect 22772 36960 22836 36964
rect 22852 37020 22916 37024
rect 22852 36964 22856 37020
rect 22856 36964 22912 37020
rect 22912 36964 22916 37020
rect 22852 36960 22916 36964
rect 27612 37020 27676 37024
rect 27612 36964 27616 37020
rect 27616 36964 27672 37020
rect 27672 36964 27676 37020
rect 27612 36960 27676 36964
rect 27692 37020 27756 37024
rect 27692 36964 27696 37020
rect 27696 36964 27752 37020
rect 27752 36964 27756 37020
rect 27692 36960 27756 36964
rect 27772 37020 27836 37024
rect 27772 36964 27776 37020
rect 27776 36964 27832 37020
rect 27832 36964 27836 37020
rect 27772 36960 27836 36964
rect 27852 37020 27916 37024
rect 27852 36964 27856 37020
rect 27856 36964 27912 37020
rect 27912 36964 27916 37020
rect 27852 36960 27916 36964
rect 32612 37020 32676 37024
rect 32612 36964 32616 37020
rect 32616 36964 32672 37020
rect 32672 36964 32676 37020
rect 32612 36960 32676 36964
rect 32692 37020 32756 37024
rect 32692 36964 32696 37020
rect 32696 36964 32752 37020
rect 32752 36964 32756 37020
rect 32692 36960 32756 36964
rect 32772 37020 32836 37024
rect 32772 36964 32776 37020
rect 32776 36964 32832 37020
rect 32832 36964 32836 37020
rect 32772 36960 32836 36964
rect 32852 37020 32916 37024
rect 32852 36964 32856 37020
rect 32856 36964 32912 37020
rect 32912 36964 32916 37020
rect 32852 36960 32916 36964
rect 37612 37020 37676 37024
rect 37612 36964 37616 37020
rect 37616 36964 37672 37020
rect 37672 36964 37676 37020
rect 37612 36960 37676 36964
rect 37692 37020 37756 37024
rect 37692 36964 37696 37020
rect 37696 36964 37752 37020
rect 37752 36964 37756 37020
rect 37692 36960 37756 36964
rect 37772 37020 37836 37024
rect 37772 36964 37776 37020
rect 37776 36964 37832 37020
rect 37832 36964 37836 37020
rect 37772 36960 37836 36964
rect 37852 37020 37916 37024
rect 37852 36964 37856 37020
rect 37856 36964 37912 37020
rect 37912 36964 37916 37020
rect 37852 36960 37916 36964
rect 1952 36476 2016 36480
rect 1952 36420 1956 36476
rect 1956 36420 2012 36476
rect 2012 36420 2016 36476
rect 1952 36416 2016 36420
rect 2032 36476 2096 36480
rect 2032 36420 2036 36476
rect 2036 36420 2092 36476
rect 2092 36420 2096 36476
rect 2032 36416 2096 36420
rect 2112 36476 2176 36480
rect 2112 36420 2116 36476
rect 2116 36420 2172 36476
rect 2172 36420 2176 36476
rect 2112 36416 2176 36420
rect 2192 36476 2256 36480
rect 2192 36420 2196 36476
rect 2196 36420 2252 36476
rect 2252 36420 2256 36476
rect 2192 36416 2256 36420
rect 6952 36476 7016 36480
rect 6952 36420 6956 36476
rect 6956 36420 7012 36476
rect 7012 36420 7016 36476
rect 6952 36416 7016 36420
rect 7032 36476 7096 36480
rect 7032 36420 7036 36476
rect 7036 36420 7092 36476
rect 7092 36420 7096 36476
rect 7032 36416 7096 36420
rect 7112 36476 7176 36480
rect 7112 36420 7116 36476
rect 7116 36420 7172 36476
rect 7172 36420 7176 36476
rect 7112 36416 7176 36420
rect 7192 36476 7256 36480
rect 7192 36420 7196 36476
rect 7196 36420 7252 36476
rect 7252 36420 7256 36476
rect 7192 36416 7256 36420
rect 11952 36476 12016 36480
rect 11952 36420 11956 36476
rect 11956 36420 12012 36476
rect 12012 36420 12016 36476
rect 11952 36416 12016 36420
rect 12032 36476 12096 36480
rect 12032 36420 12036 36476
rect 12036 36420 12092 36476
rect 12092 36420 12096 36476
rect 12032 36416 12096 36420
rect 12112 36476 12176 36480
rect 12112 36420 12116 36476
rect 12116 36420 12172 36476
rect 12172 36420 12176 36476
rect 12112 36416 12176 36420
rect 12192 36476 12256 36480
rect 12192 36420 12196 36476
rect 12196 36420 12252 36476
rect 12252 36420 12256 36476
rect 12192 36416 12256 36420
rect 16952 36476 17016 36480
rect 16952 36420 16956 36476
rect 16956 36420 17012 36476
rect 17012 36420 17016 36476
rect 16952 36416 17016 36420
rect 17032 36476 17096 36480
rect 17032 36420 17036 36476
rect 17036 36420 17092 36476
rect 17092 36420 17096 36476
rect 17032 36416 17096 36420
rect 17112 36476 17176 36480
rect 17112 36420 17116 36476
rect 17116 36420 17172 36476
rect 17172 36420 17176 36476
rect 17112 36416 17176 36420
rect 17192 36476 17256 36480
rect 17192 36420 17196 36476
rect 17196 36420 17252 36476
rect 17252 36420 17256 36476
rect 17192 36416 17256 36420
rect 21952 36476 22016 36480
rect 21952 36420 21956 36476
rect 21956 36420 22012 36476
rect 22012 36420 22016 36476
rect 21952 36416 22016 36420
rect 22032 36476 22096 36480
rect 22032 36420 22036 36476
rect 22036 36420 22092 36476
rect 22092 36420 22096 36476
rect 22032 36416 22096 36420
rect 22112 36476 22176 36480
rect 22112 36420 22116 36476
rect 22116 36420 22172 36476
rect 22172 36420 22176 36476
rect 22112 36416 22176 36420
rect 22192 36476 22256 36480
rect 22192 36420 22196 36476
rect 22196 36420 22252 36476
rect 22252 36420 22256 36476
rect 22192 36416 22256 36420
rect 26952 36476 27016 36480
rect 26952 36420 26956 36476
rect 26956 36420 27012 36476
rect 27012 36420 27016 36476
rect 26952 36416 27016 36420
rect 27032 36476 27096 36480
rect 27032 36420 27036 36476
rect 27036 36420 27092 36476
rect 27092 36420 27096 36476
rect 27032 36416 27096 36420
rect 27112 36476 27176 36480
rect 27112 36420 27116 36476
rect 27116 36420 27172 36476
rect 27172 36420 27176 36476
rect 27112 36416 27176 36420
rect 27192 36476 27256 36480
rect 27192 36420 27196 36476
rect 27196 36420 27252 36476
rect 27252 36420 27256 36476
rect 27192 36416 27256 36420
rect 31952 36476 32016 36480
rect 31952 36420 31956 36476
rect 31956 36420 32012 36476
rect 32012 36420 32016 36476
rect 31952 36416 32016 36420
rect 32032 36476 32096 36480
rect 32032 36420 32036 36476
rect 32036 36420 32092 36476
rect 32092 36420 32096 36476
rect 32032 36416 32096 36420
rect 32112 36476 32176 36480
rect 32112 36420 32116 36476
rect 32116 36420 32172 36476
rect 32172 36420 32176 36476
rect 32112 36416 32176 36420
rect 32192 36476 32256 36480
rect 32192 36420 32196 36476
rect 32196 36420 32252 36476
rect 32252 36420 32256 36476
rect 32192 36416 32256 36420
rect 36952 36476 37016 36480
rect 36952 36420 36956 36476
rect 36956 36420 37012 36476
rect 37012 36420 37016 36476
rect 36952 36416 37016 36420
rect 37032 36476 37096 36480
rect 37032 36420 37036 36476
rect 37036 36420 37092 36476
rect 37092 36420 37096 36476
rect 37032 36416 37096 36420
rect 37112 36476 37176 36480
rect 37112 36420 37116 36476
rect 37116 36420 37172 36476
rect 37172 36420 37176 36476
rect 37112 36416 37176 36420
rect 37192 36476 37256 36480
rect 37192 36420 37196 36476
rect 37196 36420 37252 36476
rect 37252 36420 37256 36476
rect 37192 36416 37256 36420
rect 2612 35932 2676 35936
rect 2612 35876 2616 35932
rect 2616 35876 2672 35932
rect 2672 35876 2676 35932
rect 2612 35872 2676 35876
rect 2692 35932 2756 35936
rect 2692 35876 2696 35932
rect 2696 35876 2752 35932
rect 2752 35876 2756 35932
rect 2692 35872 2756 35876
rect 2772 35932 2836 35936
rect 2772 35876 2776 35932
rect 2776 35876 2832 35932
rect 2832 35876 2836 35932
rect 2772 35872 2836 35876
rect 2852 35932 2916 35936
rect 2852 35876 2856 35932
rect 2856 35876 2912 35932
rect 2912 35876 2916 35932
rect 2852 35872 2916 35876
rect 7612 35932 7676 35936
rect 7612 35876 7616 35932
rect 7616 35876 7672 35932
rect 7672 35876 7676 35932
rect 7612 35872 7676 35876
rect 7692 35932 7756 35936
rect 7692 35876 7696 35932
rect 7696 35876 7752 35932
rect 7752 35876 7756 35932
rect 7692 35872 7756 35876
rect 7772 35932 7836 35936
rect 7772 35876 7776 35932
rect 7776 35876 7832 35932
rect 7832 35876 7836 35932
rect 7772 35872 7836 35876
rect 7852 35932 7916 35936
rect 7852 35876 7856 35932
rect 7856 35876 7912 35932
rect 7912 35876 7916 35932
rect 7852 35872 7916 35876
rect 12612 35932 12676 35936
rect 12612 35876 12616 35932
rect 12616 35876 12672 35932
rect 12672 35876 12676 35932
rect 12612 35872 12676 35876
rect 12692 35932 12756 35936
rect 12692 35876 12696 35932
rect 12696 35876 12752 35932
rect 12752 35876 12756 35932
rect 12692 35872 12756 35876
rect 12772 35932 12836 35936
rect 12772 35876 12776 35932
rect 12776 35876 12832 35932
rect 12832 35876 12836 35932
rect 12772 35872 12836 35876
rect 12852 35932 12916 35936
rect 12852 35876 12856 35932
rect 12856 35876 12912 35932
rect 12912 35876 12916 35932
rect 12852 35872 12916 35876
rect 17612 35932 17676 35936
rect 17612 35876 17616 35932
rect 17616 35876 17672 35932
rect 17672 35876 17676 35932
rect 17612 35872 17676 35876
rect 17692 35932 17756 35936
rect 17692 35876 17696 35932
rect 17696 35876 17752 35932
rect 17752 35876 17756 35932
rect 17692 35872 17756 35876
rect 17772 35932 17836 35936
rect 17772 35876 17776 35932
rect 17776 35876 17832 35932
rect 17832 35876 17836 35932
rect 17772 35872 17836 35876
rect 17852 35932 17916 35936
rect 17852 35876 17856 35932
rect 17856 35876 17912 35932
rect 17912 35876 17916 35932
rect 17852 35872 17916 35876
rect 22612 35932 22676 35936
rect 22612 35876 22616 35932
rect 22616 35876 22672 35932
rect 22672 35876 22676 35932
rect 22612 35872 22676 35876
rect 22692 35932 22756 35936
rect 22692 35876 22696 35932
rect 22696 35876 22752 35932
rect 22752 35876 22756 35932
rect 22692 35872 22756 35876
rect 22772 35932 22836 35936
rect 22772 35876 22776 35932
rect 22776 35876 22832 35932
rect 22832 35876 22836 35932
rect 22772 35872 22836 35876
rect 22852 35932 22916 35936
rect 22852 35876 22856 35932
rect 22856 35876 22912 35932
rect 22912 35876 22916 35932
rect 22852 35872 22916 35876
rect 27612 35932 27676 35936
rect 27612 35876 27616 35932
rect 27616 35876 27672 35932
rect 27672 35876 27676 35932
rect 27612 35872 27676 35876
rect 27692 35932 27756 35936
rect 27692 35876 27696 35932
rect 27696 35876 27752 35932
rect 27752 35876 27756 35932
rect 27692 35872 27756 35876
rect 27772 35932 27836 35936
rect 27772 35876 27776 35932
rect 27776 35876 27832 35932
rect 27832 35876 27836 35932
rect 27772 35872 27836 35876
rect 27852 35932 27916 35936
rect 27852 35876 27856 35932
rect 27856 35876 27912 35932
rect 27912 35876 27916 35932
rect 27852 35872 27916 35876
rect 32612 35932 32676 35936
rect 32612 35876 32616 35932
rect 32616 35876 32672 35932
rect 32672 35876 32676 35932
rect 32612 35872 32676 35876
rect 32692 35932 32756 35936
rect 32692 35876 32696 35932
rect 32696 35876 32752 35932
rect 32752 35876 32756 35932
rect 32692 35872 32756 35876
rect 32772 35932 32836 35936
rect 32772 35876 32776 35932
rect 32776 35876 32832 35932
rect 32832 35876 32836 35932
rect 32772 35872 32836 35876
rect 32852 35932 32916 35936
rect 32852 35876 32856 35932
rect 32856 35876 32912 35932
rect 32912 35876 32916 35932
rect 32852 35872 32916 35876
rect 37612 35932 37676 35936
rect 37612 35876 37616 35932
rect 37616 35876 37672 35932
rect 37672 35876 37676 35932
rect 37612 35872 37676 35876
rect 37692 35932 37756 35936
rect 37692 35876 37696 35932
rect 37696 35876 37752 35932
rect 37752 35876 37756 35932
rect 37692 35872 37756 35876
rect 37772 35932 37836 35936
rect 37772 35876 37776 35932
rect 37776 35876 37832 35932
rect 37832 35876 37836 35932
rect 37772 35872 37836 35876
rect 37852 35932 37916 35936
rect 37852 35876 37856 35932
rect 37856 35876 37912 35932
rect 37912 35876 37916 35932
rect 37852 35872 37916 35876
rect 1952 35388 2016 35392
rect 1952 35332 1956 35388
rect 1956 35332 2012 35388
rect 2012 35332 2016 35388
rect 1952 35328 2016 35332
rect 2032 35388 2096 35392
rect 2032 35332 2036 35388
rect 2036 35332 2092 35388
rect 2092 35332 2096 35388
rect 2032 35328 2096 35332
rect 2112 35388 2176 35392
rect 2112 35332 2116 35388
rect 2116 35332 2172 35388
rect 2172 35332 2176 35388
rect 2112 35328 2176 35332
rect 2192 35388 2256 35392
rect 2192 35332 2196 35388
rect 2196 35332 2252 35388
rect 2252 35332 2256 35388
rect 2192 35328 2256 35332
rect 6952 35388 7016 35392
rect 6952 35332 6956 35388
rect 6956 35332 7012 35388
rect 7012 35332 7016 35388
rect 6952 35328 7016 35332
rect 7032 35388 7096 35392
rect 7032 35332 7036 35388
rect 7036 35332 7092 35388
rect 7092 35332 7096 35388
rect 7032 35328 7096 35332
rect 7112 35388 7176 35392
rect 7112 35332 7116 35388
rect 7116 35332 7172 35388
rect 7172 35332 7176 35388
rect 7112 35328 7176 35332
rect 7192 35388 7256 35392
rect 7192 35332 7196 35388
rect 7196 35332 7252 35388
rect 7252 35332 7256 35388
rect 7192 35328 7256 35332
rect 11952 35388 12016 35392
rect 11952 35332 11956 35388
rect 11956 35332 12012 35388
rect 12012 35332 12016 35388
rect 11952 35328 12016 35332
rect 12032 35388 12096 35392
rect 12032 35332 12036 35388
rect 12036 35332 12092 35388
rect 12092 35332 12096 35388
rect 12032 35328 12096 35332
rect 12112 35388 12176 35392
rect 12112 35332 12116 35388
rect 12116 35332 12172 35388
rect 12172 35332 12176 35388
rect 12112 35328 12176 35332
rect 12192 35388 12256 35392
rect 12192 35332 12196 35388
rect 12196 35332 12252 35388
rect 12252 35332 12256 35388
rect 12192 35328 12256 35332
rect 16952 35388 17016 35392
rect 16952 35332 16956 35388
rect 16956 35332 17012 35388
rect 17012 35332 17016 35388
rect 16952 35328 17016 35332
rect 17032 35388 17096 35392
rect 17032 35332 17036 35388
rect 17036 35332 17092 35388
rect 17092 35332 17096 35388
rect 17032 35328 17096 35332
rect 17112 35388 17176 35392
rect 17112 35332 17116 35388
rect 17116 35332 17172 35388
rect 17172 35332 17176 35388
rect 17112 35328 17176 35332
rect 17192 35388 17256 35392
rect 17192 35332 17196 35388
rect 17196 35332 17252 35388
rect 17252 35332 17256 35388
rect 17192 35328 17256 35332
rect 21952 35388 22016 35392
rect 21952 35332 21956 35388
rect 21956 35332 22012 35388
rect 22012 35332 22016 35388
rect 21952 35328 22016 35332
rect 22032 35388 22096 35392
rect 22032 35332 22036 35388
rect 22036 35332 22092 35388
rect 22092 35332 22096 35388
rect 22032 35328 22096 35332
rect 22112 35388 22176 35392
rect 22112 35332 22116 35388
rect 22116 35332 22172 35388
rect 22172 35332 22176 35388
rect 22112 35328 22176 35332
rect 22192 35388 22256 35392
rect 22192 35332 22196 35388
rect 22196 35332 22252 35388
rect 22252 35332 22256 35388
rect 22192 35328 22256 35332
rect 26952 35388 27016 35392
rect 26952 35332 26956 35388
rect 26956 35332 27012 35388
rect 27012 35332 27016 35388
rect 26952 35328 27016 35332
rect 27032 35388 27096 35392
rect 27032 35332 27036 35388
rect 27036 35332 27092 35388
rect 27092 35332 27096 35388
rect 27032 35328 27096 35332
rect 27112 35388 27176 35392
rect 27112 35332 27116 35388
rect 27116 35332 27172 35388
rect 27172 35332 27176 35388
rect 27112 35328 27176 35332
rect 27192 35388 27256 35392
rect 27192 35332 27196 35388
rect 27196 35332 27252 35388
rect 27252 35332 27256 35388
rect 27192 35328 27256 35332
rect 31952 35388 32016 35392
rect 31952 35332 31956 35388
rect 31956 35332 32012 35388
rect 32012 35332 32016 35388
rect 31952 35328 32016 35332
rect 32032 35388 32096 35392
rect 32032 35332 32036 35388
rect 32036 35332 32092 35388
rect 32092 35332 32096 35388
rect 32032 35328 32096 35332
rect 32112 35388 32176 35392
rect 32112 35332 32116 35388
rect 32116 35332 32172 35388
rect 32172 35332 32176 35388
rect 32112 35328 32176 35332
rect 32192 35388 32256 35392
rect 32192 35332 32196 35388
rect 32196 35332 32252 35388
rect 32252 35332 32256 35388
rect 32192 35328 32256 35332
rect 36952 35388 37016 35392
rect 36952 35332 36956 35388
rect 36956 35332 37012 35388
rect 37012 35332 37016 35388
rect 36952 35328 37016 35332
rect 37032 35388 37096 35392
rect 37032 35332 37036 35388
rect 37036 35332 37092 35388
rect 37092 35332 37096 35388
rect 37032 35328 37096 35332
rect 37112 35388 37176 35392
rect 37112 35332 37116 35388
rect 37116 35332 37172 35388
rect 37172 35332 37176 35388
rect 37112 35328 37176 35332
rect 37192 35388 37256 35392
rect 37192 35332 37196 35388
rect 37196 35332 37252 35388
rect 37252 35332 37256 35388
rect 37192 35328 37256 35332
rect 2612 34844 2676 34848
rect 2612 34788 2616 34844
rect 2616 34788 2672 34844
rect 2672 34788 2676 34844
rect 2612 34784 2676 34788
rect 2692 34844 2756 34848
rect 2692 34788 2696 34844
rect 2696 34788 2752 34844
rect 2752 34788 2756 34844
rect 2692 34784 2756 34788
rect 2772 34844 2836 34848
rect 2772 34788 2776 34844
rect 2776 34788 2832 34844
rect 2832 34788 2836 34844
rect 2772 34784 2836 34788
rect 2852 34844 2916 34848
rect 2852 34788 2856 34844
rect 2856 34788 2912 34844
rect 2912 34788 2916 34844
rect 2852 34784 2916 34788
rect 7612 34844 7676 34848
rect 7612 34788 7616 34844
rect 7616 34788 7672 34844
rect 7672 34788 7676 34844
rect 7612 34784 7676 34788
rect 7692 34844 7756 34848
rect 7692 34788 7696 34844
rect 7696 34788 7752 34844
rect 7752 34788 7756 34844
rect 7692 34784 7756 34788
rect 7772 34844 7836 34848
rect 7772 34788 7776 34844
rect 7776 34788 7832 34844
rect 7832 34788 7836 34844
rect 7772 34784 7836 34788
rect 7852 34844 7916 34848
rect 7852 34788 7856 34844
rect 7856 34788 7912 34844
rect 7912 34788 7916 34844
rect 7852 34784 7916 34788
rect 12612 34844 12676 34848
rect 12612 34788 12616 34844
rect 12616 34788 12672 34844
rect 12672 34788 12676 34844
rect 12612 34784 12676 34788
rect 12692 34844 12756 34848
rect 12692 34788 12696 34844
rect 12696 34788 12752 34844
rect 12752 34788 12756 34844
rect 12692 34784 12756 34788
rect 12772 34844 12836 34848
rect 12772 34788 12776 34844
rect 12776 34788 12832 34844
rect 12832 34788 12836 34844
rect 12772 34784 12836 34788
rect 12852 34844 12916 34848
rect 12852 34788 12856 34844
rect 12856 34788 12912 34844
rect 12912 34788 12916 34844
rect 12852 34784 12916 34788
rect 17612 34844 17676 34848
rect 17612 34788 17616 34844
rect 17616 34788 17672 34844
rect 17672 34788 17676 34844
rect 17612 34784 17676 34788
rect 17692 34844 17756 34848
rect 17692 34788 17696 34844
rect 17696 34788 17752 34844
rect 17752 34788 17756 34844
rect 17692 34784 17756 34788
rect 17772 34844 17836 34848
rect 17772 34788 17776 34844
rect 17776 34788 17832 34844
rect 17832 34788 17836 34844
rect 17772 34784 17836 34788
rect 17852 34844 17916 34848
rect 17852 34788 17856 34844
rect 17856 34788 17912 34844
rect 17912 34788 17916 34844
rect 17852 34784 17916 34788
rect 22612 34844 22676 34848
rect 22612 34788 22616 34844
rect 22616 34788 22672 34844
rect 22672 34788 22676 34844
rect 22612 34784 22676 34788
rect 22692 34844 22756 34848
rect 22692 34788 22696 34844
rect 22696 34788 22752 34844
rect 22752 34788 22756 34844
rect 22692 34784 22756 34788
rect 22772 34844 22836 34848
rect 22772 34788 22776 34844
rect 22776 34788 22832 34844
rect 22832 34788 22836 34844
rect 22772 34784 22836 34788
rect 22852 34844 22916 34848
rect 22852 34788 22856 34844
rect 22856 34788 22912 34844
rect 22912 34788 22916 34844
rect 22852 34784 22916 34788
rect 27612 34844 27676 34848
rect 27612 34788 27616 34844
rect 27616 34788 27672 34844
rect 27672 34788 27676 34844
rect 27612 34784 27676 34788
rect 27692 34844 27756 34848
rect 27692 34788 27696 34844
rect 27696 34788 27752 34844
rect 27752 34788 27756 34844
rect 27692 34784 27756 34788
rect 27772 34844 27836 34848
rect 27772 34788 27776 34844
rect 27776 34788 27832 34844
rect 27832 34788 27836 34844
rect 27772 34784 27836 34788
rect 27852 34844 27916 34848
rect 27852 34788 27856 34844
rect 27856 34788 27912 34844
rect 27912 34788 27916 34844
rect 27852 34784 27916 34788
rect 32612 34844 32676 34848
rect 32612 34788 32616 34844
rect 32616 34788 32672 34844
rect 32672 34788 32676 34844
rect 32612 34784 32676 34788
rect 32692 34844 32756 34848
rect 32692 34788 32696 34844
rect 32696 34788 32752 34844
rect 32752 34788 32756 34844
rect 32692 34784 32756 34788
rect 32772 34844 32836 34848
rect 32772 34788 32776 34844
rect 32776 34788 32832 34844
rect 32832 34788 32836 34844
rect 32772 34784 32836 34788
rect 32852 34844 32916 34848
rect 32852 34788 32856 34844
rect 32856 34788 32912 34844
rect 32912 34788 32916 34844
rect 32852 34784 32916 34788
rect 37612 34844 37676 34848
rect 37612 34788 37616 34844
rect 37616 34788 37672 34844
rect 37672 34788 37676 34844
rect 37612 34784 37676 34788
rect 37692 34844 37756 34848
rect 37692 34788 37696 34844
rect 37696 34788 37752 34844
rect 37752 34788 37756 34844
rect 37692 34784 37756 34788
rect 37772 34844 37836 34848
rect 37772 34788 37776 34844
rect 37776 34788 37832 34844
rect 37832 34788 37836 34844
rect 37772 34784 37836 34788
rect 37852 34844 37916 34848
rect 37852 34788 37856 34844
rect 37856 34788 37912 34844
rect 37912 34788 37916 34844
rect 37852 34784 37916 34788
rect 1952 34300 2016 34304
rect 1952 34244 1956 34300
rect 1956 34244 2012 34300
rect 2012 34244 2016 34300
rect 1952 34240 2016 34244
rect 2032 34300 2096 34304
rect 2032 34244 2036 34300
rect 2036 34244 2092 34300
rect 2092 34244 2096 34300
rect 2032 34240 2096 34244
rect 2112 34300 2176 34304
rect 2112 34244 2116 34300
rect 2116 34244 2172 34300
rect 2172 34244 2176 34300
rect 2112 34240 2176 34244
rect 2192 34300 2256 34304
rect 2192 34244 2196 34300
rect 2196 34244 2252 34300
rect 2252 34244 2256 34300
rect 2192 34240 2256 34244
rect 6952 34300 7016 34304
rect 6952 34244 6956 34300
rect 6956 34244 7012 34300
rect 7012 34244 7016 34300
rect 6952 34240 7016 34244
rect 7032 34300 7096 34304
rect 7032 34244 7036 34300
rect 7036 34244 7092 34300
rect 7092 34244 7096 34300
rect 7032 34240 7096 34244
rect 7112 34300 7176 34304
rect 7112 34244 7116 34300
rect 7116 34244 7172 34300
rect 7172 34244 7176 34300
rect 7112 34240 7176 34244
rect 7192 34300 7256 34304
rect 7192 34244 7196 34300
rect 7196 34244 7252 34300
rect 7252 34244 7256 34300
rect 7192 34240 7256 34244
rect 11952 34300 12016 34304
rect 11952 34244 11956 34300
rect 11956 34244 12012 34300
rect 12012 34244 12016 34300
rect 11952 34240 12016 34244
rect 12032 34300 12096 34304
rect 12032 34244 12036 34300
rect 12036 34244 12092 34300
rect 12092 34244 12096 34300
rect 12032 34240 12096 34244
rect 12112 34300 12176 34304
rect 12112 34244 12116 34300
rect 12116 34244 12172 34300
rect 12172 34244 12176 34300
rect 12112 34240 12176 34244
rect 12192 34300 12256 34304
rect 12192 34244 12196 34300
rect 12196 34244 12252 34300
rect 12252 34244 12256 34300
rect 12192 34240 12256 34244
rect 16952 34300 17016 34304
rect 16952 34244 16956 34300
rect 16956 34244 17012 34300
rect 17012 34244 17016 34300
rect 16952 34240 17016 34244
rect 17032 34300 17096 34304
rect 17032 34244 17036 34300
rect 17036 34244 17092 34300
rect 17092 34244 17096 34300
rect 17032 34240 17096 34244
rect 17112 34300 17176 34304
rect 17112 34244 17116 34300
rect 17116 34244 17172 34300
rect 17172 34244 17176 34300
rect 17112 34240 17176 34244
rect 17192 34300 17256 34304
rect 17192 34244 17196 34300
rect 17196 34244 17252 34300
rect 17252 34244 17256 34300
rect 17192 34240 17256 34244
rect 21952 34300 22016 34304
rect 21952 34244 21956 34300
rect 21956 34244 22012 34300
rect 22012 34244 22016 34300
rect 21952 34240 22016 34244
rect 22032 34300 22096 34304
rect 22032 34244 22036 34300
rect 22036 34244 22092 34300
rect 22092 34244 22096 34300
rect 22032 34240 22096 34244
rect 22112 34300 22176 34304
rect 22112 34244 22116 34300
rect 22116 34244 22172 34300
rect 22172 34244 22176 34300
rect 22112 34240 22176 34244
rect 22192 34300 22256 34304
rect 22192 34244 22196 34300
rect 22196 34244 22252 34300
rect 22252 34244 22256 34300
rect 22192 34240 22256 34244
rect 26952 34300 27016 34304
rect 26952 34244 26956 34300
rect 26956 34244 27012 34300
rect 27012 34244 27016 34300
rect 26952 34240 27016 34244
rect 27032 34300 27096 34304
rect 27032 34244 27036 34300
rect 27036 34244 27092 34300
rect 27092 34244 27096 34300
rect 27032 34240 27096 34244
rect 27112 34300 27176 34304
rect 27112 34244 27116 34300
rect 27116 34244 27172 34300
rect 27172 34244 27176 34300
rect 27112 34240 27176 34244
rect 27192 34300 27256 34304
rect 27192 34244 27196 34300
rect 27196 34244 27252 34300
rect 27252 34244 27256 34300
rect 27192 34240 27256 34244
rect 31952 34300 32016 34304
rect 31952 34244 31956 34300
rect 31956 34244 32012 34300
rect 32012 34244 32016 34300
rect 31952 34240 32016 34244
rect 32032 34300 32096 34304
rect 32032 34244 32036 34300
rect 32036 34244 32092 34300
rect 32092 34244 32096 34300
rect 32032 34240 32096 34244
rect 32112 34300 32176 34304
rect 32112 34244 32116 34300
rect 32116 34244 32172 34300
rect 32172 34244 32176 34300
rect 32112 34240 32176 34244
rect 32192 34300 32256 34304
rect 32192 34244 32196 34300
rect 32196 34244 32252 34300
rect 32252 34244 32256 34300
rect 32192 34240 32256 34244
rect 36952 34300 37016 34304
rect 36952 34244 36956 34300
rect 36956 34244 37012 34300
rect 37012 34244 37016 34300
rect 36952 34240 37016 34244
rect 37032 34300 37096 34304
rect 37032 34244 37036 34300
rect 37036 34244 37092 34300
rect 37092 34244 37096 34300
rect 37032 34240 37096 34244
rect 37112 34300 37176 34304
rect 37112 34244 37116 34300
rect 37116 34244 37172 34300
rect 37172 34244 37176 34300
rect 37112 34240 37176 34244
rect 37192 34300 37256 34304
rect 37192 34244 37196 34300
rect 37196 34244 37252 34300
rect 37252 34244 37256 34300
rect 37192 34240 37256 34244
rect 2612 33756 2676 33760
rect 2612 33700 2616 33756
rect 2616 33700 2672 33756
rect 2672 33700 2676 33756
rect 2612 33696 2676 33700
rect 2692 33756 2756 33760
rect 2692 33700 2696 33756
rect 2696 33700 2752 33756
rect 2752 33700 2756 33756
rect 2692 33696 2756 33700
rect 2772 33756 2836 33760
rect 2772 33700 2776 33756
rect 2776 33700 2832 33756
rect 2832 33700 2836 33756
rect 2772 33696 2836 33700
rect 2852 33756 2916 33760
rect 2852 33700 2856 33756
rect 2856 33700 2912 33756
rect 2912 33700 2916 33756
rect 2852 33696 2916 33700
rect 7612 33756 7676 33760
rect 7612 33700 7616 33756
rect 7616 33700 7672 33756
rect 7672 33700 7676 33756
rect 7612 33696 7676 33700
rect 7692 33756 7756 33760
rect 7692 33700 7696 33756
rect 7696 33700 7752 33756
rect 7752 33700 7756 33756
rect 7692 33696 7756 33700
rect 7772 33756 7836 33760
rect 7772 33700 7776 33756
rect 7776 33700 7832 33756
rect 7832 33700 7836 33756
rect 7772 33696 7836 33700
rect 7852 33756 7916 33760
rect 7852 33700 7856 33756
rect 7856 33700 7912 33756
rect 7912 33700 7916 33756
rect 7852 33696 7916 33700
rect 12612 33756 12676 33760
rect 12612 33700 12616 33756
rect 12616 33700 12672 33756
rect 12672 33700 12676 33756
rect 12612 33696 12676 33700
rect 12692 33756 12756 33760
rect 12692 33700 12696 33756
rect 12696 33700 12752 33756
rect 12752 33700 12756 33756
rect 12692 33696 12756 33700
rect 12772 33756 12836 33760
rect 12772 33700 12776 33756
rect 12776 33700 12832 33756
rect 12832 33700 12836 33756
rect 12772 33696 12836 33700
rect 12852 33756 12916 33760
rect 12852 33700 12856 33756
rect 12856 33700 12912 33756
rect 12912 33700 12916 33756
rect 12852 33696 12916 33700
rect 17612 33756 17676 33760
rect 17612 33700 17616 33756
rect 17616 33700 17672 33756
rect 17672 33700 17676 33756
rect 17612 33696 17676 33700
rect 17692 33756 17756 33760
rect 17692 33700 17696 33756
rect 17696 33700 17752 33756
rect 17752 33700 17756 33756
rect 17692 33696 17756 33700
rect 17772 33756 17836 33760
rect 17772 33700 17776 33756
rect 17776 33700 17832 33756
rect 17832 33700 17836 33756
rect 17772 33696 17836 33700
rect 17852 33756 17916 33760
rect 17852 33700 17856 33756
rect 17856 33700 17912 33756
rect 17912 33700 17916 33756
rect 17852 33696 17916 33700
rect 22612 33756 22676 33760
rect 22612 33700 22616 33756
rect 22616 33700 22672 33756
rect 22672 33700 22676 33756
rect 22612 33696 22676 33700
rect 22692 33756 22756 33760
rect 22692 33700 22696 33756
rect 22696 33700 22752 33756
rect 22752 33700 22756 33756
rect 22692 33696 22756 33700
rect 22772 33756 22836 33760
rect 22772 33700 22776 33756
rect 22776 33700 22832 33756
rect 22832 33700 22836 33756
rect 22772 33696 22836 33700
rect 22852 33756 22916 33760
rect 22852 33700 22856 33756
rect 22856 33700 22912 33756
rect 22912 33700 22916 33756
rect 22852 33696 22916 33700
rect 27612 33756 27676 33760
rect 27612 33700 27616 33756
rect 27616 33700 27672 33756
rect 27672 33700 27676 33756
rect 27612 33696 27676 33700
rect 27692 33756 27756 33760
rect 27692 33700 27696 33756
rect 27696 33700 27752 33756
rect 27752 33700 27756 33756
rect 27692 33696 27756 33700
rect 27772 33756 27836 33760
rect 27772 33700 27776 33756
rect 27776 33700 27832 33756
rect 27832 33700 27836 33756
rect 27772 33696 27836 33700
rect 27852 33756 27916 33760
rect 27852 33700 27856 33756
rect 27856 33700 27912 33756
rect 27912 33700 27916 33756
rect 27852 33696 27916 33700
rect 32612 33756 32676 33760
rect 32612 33700 32616 33756
rect 32616 33700 32672 33756
rect 32672 33700 32676 33756
rect 32612 33696 32676 33700
rect 32692 33756 32756 33760
rect 32692 33700 32696 33756
rect 32696 33700 32752 33756
rect 32752 33700 32756 33756
rect 32692 33696 32756 33700
rect 32772 33756 32836 33760
rect 32772 33700 32776 33756
rect 32776 33700 32832 33756
rect 32832 33700 32836 33756
rect 32772 33696 32836 33700
rect 32852 33756 32916 33760
rect 32852 33700 32856 33756
rect 32856 33700 32912 33756
rect 32912 33700 32916 33756
rect 32852 33696 32916 33700
rect 37612 33756 37676 33760
rect 37612 33700 37616 33756
rect 37616 33700 37672 33756
rect 37672 33700 37676 33756
rect 37612 33696 37676 33700
rect 37692 33756 37756 33760
rect 37692 33700 37696 33756
rect 37696 33700 37752 33756
rect 37752 33700 37756 33756
rect 37692 33696 37756 33700
rect 37772 33756 37836 33760
rect 37772 33700 37776 33756
rect 37776 33700 37832 33756
rect 37832 33700 37836 33756
rect 37772 33696 37836 33700
rect 37852 33756 37916 33760
rect 37852 33700 37856 33756
rect 37856 33700 37912 33756
rect 37912 33700 37916 33756
rect 37852 33696 37916 33700
rect 1952 33212 2016 33216
rect 1952 33156 1956 33212
rect 1956 33156 2012 33212
rect 2012 33156 2016 33212
rect 1952 33152 2016 33156
rect 2032 33212 2096 33216
rect 2032 33156 2036 33212
rect 2036 33156 2092 33212
rect 2092 33156 2096 33212
rect 2032 33152 2096 33156
rect 2112 33212 2176 33216
rect 2112 33156 2116 33212
rect 2116 33156 2172 33212
rect 2172 33156 2176 33212
rect 2112 33152 2176 33156
rect 2192 33212 2256 33216
rect 2192 33156 2196 33212
rect 2196 33156 2252 33212
rect 2252 33156 2256 33212
rect 2192 33152 2256 33156
rect 6952 33212 7016 33216
rect 6952 33156 6956 33212
rect 6956 33156 7012 33212
rect 7012 33156 7016 33212
rect 6952 33152 7016 33156
rect 7032 33212 7096 33216
rect 7032 33156 7036 33212
rect 7036 33156 7092 33212
rect 7092 33156 7096 33212
rect 7032 33152 7096 33156
rect 7112 33212 7176 33216
rect 7112 33156 7116 33212
rect 7116 33156 7172 33212
rect 7172 33156 7176 33212
rect 7112 33152 7176 33156
rect 7192 33212 7256 33216
rect 7192 33156 7196 33212
rect 7196 33156 7252 33212
rect 7252 33156 7256 33212
rect 7192 33152 7256 33156
rect 11952 33212 12016 33216
rect 11952 33156 11956 33212
rect 11956 33156 12012 33212
rect 12012 33156 12016 33212
rect 11952 33152 12016 33156
rect 12032 33212 12096 33216
rect 12032 33156 12036 33212
rect 12036 33156 12092 33212
rect 12092 33156 12096 33212
rect 12032 33152 12096 33156
rect 12112 33212 12176 33216
rect 12112 33156 12116 33212
rect 12116 33156 12172 33212
rect 12172 33156 12176 33212
rect 12112 33152 12176 33156
rect 12192 33212 12256 33216
rect 12192 33156 12196 33212
rect 12196 33156 12252 33212
rect 12252 33156 12256 33212
rect 12192 33152 12256 33156
rect 16952 33212 17016 33216
rect 16952 33156 16956 33212
rect 16956 33156 17012 33212
rect 17012 33156 17016 33212
rect 16952 33152 17016 33156
rect 17032 33212 17096 33216
rect 17032 33156 17036 33212
rect 17036 33156 17092 33212
rect 17092 33156 17096 33212
rect 17032 33152 17096 33156
rect 17112 33212 17176 33216
rect 17112 33156 17116 33212
rect 17116 33156 17172 33212
rect 17172 33156 17176 33212
rect 17112 33152 17176 33156
rect 17192 33212 17256 33216
rect 17192 33156 17196 33212
rect 17196 33156 17252 33212
rect 17252 33156 17256 33212
rect 17192 33152 17256 33156
rect 21952 33212 22016 33216
rect 21952 33156 21956 33212
rect 21956 33156 22012 33212
rect 22012 33156 22016 33212
rect 21952 33152 22016 33156
rect 22032 33212 22096 33216
rect 22032 33156 22036 33212
rect 22036 33156 22092 33212
rect 22092 33156 22096 33212
rect 22032 33152 22096 33156
rect 22112 33212 22176 33216
rect 22112 33156 22116 33212
rect 22116 33156 22172 33212
rect 22172 33156 22176 33212
rect 22112 33152 22176 33156
rect 22192 33212 22256 33216
rect 22192 33156 22196 33212
rect 22196 33156 22252 33212
rect 22252 33156 22256 33212
rect 22192 33152 22256 33156
rect 26952 33212 27016 33216
rect 26952 33156 26956 33212
rect 26956 33156 27012 33212
rect 27012 33156 27016 33212
rect 26952 33152 27016 33156
rect 27032 33212 27096 33216
rect 27032 33156 27036 33212
rect 27036 33156 27092 33212
rect 27092 33156 27096 33212
rect 27032 33152 27096 33156
rect 27112 33212 27176 33216
rect 27112 33156 27116 33212
rect 27116 33156 27172 33212
rect 27172 33156 27176 33212
rect 27112 33152 27176 33156
rect 27192 33212 27256 33216
rect 27192 33156 27196 33212
rect 27196 33156 27252 33212
rect 27252 33156 27256 33212
rect 27192 33152 27256 33156
rect 31952 33212 32016 33216
rect 31952 33156 31956 33212
rect 31956 33156 32012 33212
rect 32012 33156 32016 33212
rect 31952 33152 32016 33156
rect 32032 33212 32096 33216
rect 32032 33156 32036 33212
rect 32036 33156 32092 33212
rect 32092 33156 32096 33212
rect 32032 33152 32096 33156
rect 32112 33212 32176 33216
rect 32112 33156 32116 33212
rect 32116 33156 32172 33212
rect 32172 33156 32176 33212
rect 32112 33152 32176 33156
rect 32192 33212 32256 33216
rect 32192 33156 32196 33212
rect 32196 33156 32252 33212
rect 32252 33156 32256 33212
rect 32192 33152 32256 33156
rect 36952 33212 37016 33216
rect 36952 33156 36956 33212
rect 36956 33156 37012 33212
rect 37012 33156 37016 33212
rect 36952 33152 37016 33156
rect 37032 33212 37096 33216
rect 37032 33156 37036 33212
rect 37036 33156 37092 33212
rect 37092 33156 37096 33212
rect 37032 33152 37096 33156
rect 37112 33212 37176 33216
rect 37112 33156 37116 33212
rect 37116 33156 37172 33212
rect 37172 33156 37176 33212
rect 37112 33152 37176 33156
rect 37192 33212 37256 33216
rect 37192 33156 37196 33212
rect 37196 33156 37252 33212
rect 37252 33156 37256 33212
rect 37192 33152 37256 33156
rect 2612 32668 2676 32672
rect 2612 32612 2616 32668
rect 2616 32612 2672 32668
rect 2672 32612 2676 32668
rect 2612 32608 2676 32612
rect 2692 32668 2756 32672
rect 2692 32612 2696 32668
rect 2696 32612 2752 32668
rect 2752 32612 2756 32668
rect 2692 32608 2756 32612
rect 2772 32668 2836 32672
rect 2772 32612 2776 32668
rect 2776 32612 2832 32668
rect 2832 32612 2836 32668
rect 2772 32608 2836 32612
rect 2852 32668 2916 32672
rect 2852 32612 2856 32668
rect 2856 32612 2912 32668
rect 2912 32612 2916 32668
rect 2852 32608 2916 32612
rect 7612 32668 7676 32672
rect 7612 32612 7616 32668
rect 7616 32612 7672 32668
rect 7672 32612 7676 32668
rect 7612 32608 7676 32612
rect 7692 32668 7756 32672
rect 7692 32612 7696 32668
rect 7696 32612 7752 32668
rect 7752 32612 7756 32668
rect 7692 32608 7756 32612
rect 7772 32668 7836 32672
rect 7772 32612 7776 32668
rect 7776 32612 7832 32668
rect 7832 32612 7836 32668
rect 7772 32608 7836 32612
rect 7852 32668 7916 32672
rect 7852 32612 7856 32668
rect 7856 32612 7912 32668
rect 7912 32612 7916 32668
rect 7852 32608 7916 32612
rect 12612 32668 12676 32672
rect 12612 32612 12616 32668
rect 12616 32612 12672 32668
rect 12672 32612 12676 32668
rect 12612 32608 12676 32612
rect 12692 32668 12756 32672
rect 12692 32612 12696 32668
rect 12696 32612 12752 32668
rect 12752 32612 12756 32668
rect 12692 32608 12756 32612
rect 12772 32668 12836 32672
rect 12772 32612 12776 32668
rect 12776 32612 12832 32668
rect 12832 32612 12836 32668
rect 12772 32608 12836 32612
rect 12852 32668 12916 32672
rect 12852 32612 12856 32668
rect 12856 32612 12912 32668
rect 12912 32612 12916 32668
rect 12852 32608 12916 32612
rect 17612 32668 17676 32672
rect 17612 32612 17616 32668
rect 17616 32612 17672 32668
rect 17672 32612 17676 32668
rect 17612 32608 17676 32612
rect 17692 32668 17756 32672
rect 17692 32612 17696 32668
rect 17696 32612 17752 32668
rect 17752 32612 17756 32668
rect 17692 32608 17756 32612
rect 17772 32668 17836 32672
rect 17772 32612 17776 32668
rect 17776 32612 17832 32668
rect 17832 32612 17836 32668
rect 17772 32608 17836 32612
rect 17852 32668 17916 32672
rect 17852 32612 17856 32668
rect 17856 32612 17912 32668
rect 17912 32612 17916 32668
rect 17852 32608 17916 32612
rect 22612 32668 22676 32672
rect 22612 32612 22616 32668
rect 22616 32612 22672 32668
rect 22672 32612 22676 32668
rect 22612 32608 22676 32612
rect 22692 32668 22756 32672
rect 22692 32612 22696 32668
rect 22696 32612 22752 32668
rect 22752 32612 22756 32668
rect 22692 32608 22756 32612
rect 22772 32668 22836 32672
rect 22772 32612 22776 32668
rect 22776 32612 22832 32668
rect 22832 32612 22836 32668
rect 22772 32608 22836 32612
rect 22852 32668 22916 32672
rect 22852 32612 22856 32668
rect 22856 32612 22912 32668
rect 22912 32612 22916 32668
rect 22852 32608 22916 32612
rect 27612 32668 27676 32672
rect 27612 32612 27616 32668
rect 27616 32612 27672 32668
rect 27672 32612 27676 32668
rect 27612 32608 27676 32612
rect 27692 32668 27756 32672
rect 27692 32612 27696 32668
rect 27696 32612 27752 32668
rect 27752 32612 27756 32668
rect 27692 32608 27756 32612
rect 27772 32668 27836 32672
rect 27772 32612 27776 32668
rect 27776 32612 27832 32668
rect 27832 32612 27836 32668
rect 27772 32608 27836 32612
rect 27852 32668 27916 32672
rect 27852 32612 27856 32668
rect 27856 32612 27912 32668
rect 27912 32612 27916 32668
rect 27852 32608 27916 32612
rect 32612 32668 32676 32672
rect 32612 32612 32616 32668
rect 32616 32612 32672 32668
rect 32672 32612 32676 32668
rect 32612 32608 32676 32612
rect 32692 32668 32756 32672
rect 32692 32612 32696 32668
rect 32696 32612 32752 32668
rect 32752 32612 32756 32668
rect 32692 32608 32756 32612
rect 32772 32668 32836 32672
rect 32772 32612 32776 32668
rect 32776 32612 32832 32668
rect 32832 32612 32836 32668
rect 32772 32608 32836 32612
rect 32852 32668 32916 32672
rect 32852 32612 32856 32668
rect 32856 32612 32912 32668
rect 32912 32612 32916 32668
rect 32852 32608 32916 32612
rect 37612 32668 37676 32672
rect 37612 32612 37616 32668
rect 37616 32612 37672 32668
rect 37672 32612 37676 32668
rect 37612 32608 37676 32612
rect 37692 32668 37756 32672
rect 37692 32612 37696 32668
rect 37696 32612 37752 32668
rect 37752 32612 37756 32668
rect 37692 32608 37756 32612
rect 37772 32668 37836 32672
rect 37772 32612 37776 32668
rect 37776 32612 37832 32668
rect 37832 32612 37836 32668
rect 37772 32608 37836 32612
rect 37852 32668 37916 32672
rect 37852 32612 37856 32668
rect 37856 32612 37912 32668
rect 37912 32612 37916 32668
rect 37852 32608 37916 32612
rect 1952 32124 2016 32128
rect 1952 32068 1956 32124
rect 1956 32068 2012 32124
rect 2012 32068 2016 32124
rect 1952 32064 2016 32068
rect 2032 32124 2096 32128
rect 2032 32068 2036 32124
rect 2036 32068 2092 32124
rect 2092 32068 2096 32124
rect 2032 32064 2096 32068
rect 2112 32124 2176 32128
rect 2112 32068 2116 32124
rect 2116 32068 2172 32124
rect 2172 32068 2176 32124
rect 2112 32064 2176 32068
rect 2192 32124 2256 32128
rect 2192 32068 2196 32124
rect 2196 32068 2252 32124
rect 2252 32068 2256 32124
rect 2192 32064 2256 32068
rect 6952 32124 7016 32128
rect 6952 32068 6956 32124
rect 6956 32068 7012 32124
rect 7012 32068 7016 32124
rect 6952 32064 7016 32068
rect 7032 32124 7096 32128
rect 7032 32068 7036 32124
rect 7036 32068 7092 32124
rect 7092 32068 7096 32124
rect 7032 32064 7096 32068
rect 7112 32124 7176 32128
rect 7112 32068 7116 32124
rect 7116 32068 7172 32124
rect 7172 32068 7176 32124
rect 7112 32064 7176 32068
rect 7192 32124 7256 32128
rect 7192 32068 7196 32124
rect 7196 32068 7252 32124
rect 7252 32068 7256 32124
rect 7192 32064 7256 32068
rect 11952 32124 12016 32128
rect 11952 32068 11956 32124
rect 11956 32068 12012 32124
rect 12012 32068 12016 32124
rect 11952 32064 12016 32068
rect 12032 32124 12096 32128
rect 12032 32068 12036 32124
rect 12036 32068 12092 32124
rect 12092 32068 12096 32124
rect 12032 32064 12096 32068
rect 12112 32124 12176 32128
rect 12112 32068 12116 32124
rect 12116 32068 12172 32124
rect 12172 32068 12176 32124
rect 12112 32064 12176 32068
rect 12192 32124 12256 32128
rect 12192 32068 12196 32124
rect 12196 32068 12252 32124
rect 12252 32068 12256 32124
rect 12192 32064 12256 32068
rect 16952 32124 17016 32128
rect 16952 32068 16956 32124
rect 16956 32068 17012 32124
rect 17012 32068 17016 32124
rect 16952 32064 17016 32068
rect 17032 32124 17096 32128
rect 17032 32068 17036 32124
rect 17036 32068 17092 32124
rect 17092 32068 17096 32124
rect 17032 32064 17096 32068
rect 17112 32124 17176 32128
rect 17112 32068 17116 32124
rect 17116 32068 17172 32124
rect 17172 32068 17176 32124
rect 17112 32064 17176 32068
rect 17192 32124 17256 32128
rect 17192 32068 17196 32124
rect 17196 32068 17252 32124
rect 17252 32068 17256 32124
rect 17192 32064 17256 32068
rect 21952 32124 22016 32128
rect 21952 32068 21956 32124
rect 21956 32068 22012 32124
rect 22012 32068 22016 32124
rect 21952 32064 22016 32068
rect 22032 32124 22096 32128
rect 22032 32068 22036 32124
rect 22036 32068 22092 32124
rect 22092 32068 22096 32124
rect 22032 32064 22096 32068
rect 22112 32124 22176 32128
rect 22112 32068 22116 32124
rect 22116 32068 22172 32124
rect 22172 32068 22176 32124
rect 22112 32064 22176 32068
rect 22192 32124 22256 32128
rect 22192 32068 22196 32124
rect 22196 32068 22252 32124
rect 22252 32068 22256 32124
rect 22192 32064 22256 32068
rect 26952 32124 27016 32128
rect 26952 32068 26956 32124
rect 26956 32068 27012 32124
rect 27012 32068 27016 32124
rect 26952 32064 27016 32068
rect 27032 32124 27096 32128
rect 27032 32068 27036 32124
rect 27036 32068 27092 32124
rect 27092 32068 27096 32124
rect 27032 32064 27096 32068
rect 27112 32124 27176 32128
rect 27112 32068 27116 32124
rect 27116 32068 27172 32124
rect 27172 32068 27176 32124
rect 27112 32064 27176 32068
rect 27192 32124 27256 32128
rect 27192 32068 27196 32124
rect 27196 32068 27252 32124
rect 27252 32068 27256 32124
rect 27192 32064 27256 32068
rect 31952 32124 32016 32128
rect 31952 32068 31956 32124
rect 31956 32068 32012 32124
rect 32012 32068 32016 32124
rect 31952 32064 32016 32068
rect 32032 32124 32096 32128
rect 32032 32068 32036 32124
rect 32036 32068 32092 32124
rect 32092 32068 32096 32124
rect 32032 32064 32096 32068
rect 32112 32124 32176 32128
rect 32112 32068 32116 32124
rect 32116 32068 32172 32124
rect 32172 32068 32176 32124
rect 32112 32064 32176 32068
rect 32192 32124 32256 32128
rect 32192 32068 32196 32124
rect 32196 32068 32252 32124
rect 32252 32068 32256 32124
rect 32192 32064 32256 32068
rect 36952 32124 37016 32128
rect 36952 32068 36956 32124
rect 36956 32068 37012 32124
rect 37012 32068 37016 32124
rect 36952 32064 37016 32068
rect 37032 32124 37096 32128
rect 37032 32068 37036 32124
rect 37036 32068 37092 32124
rect 37092 32068 37096 32124
rect 37032 32064 37096 32068
rect 37112 32124 37176 32128
rect 37112 32068 37116 32124
rect 37116 32068 37172 32124
rect 37172 32068 37176 32124
rect 37112 32064 37176 32068
rect 37192 32124 37256 32128
rect 37192 32068 37196 32124
rect 37196 32068 37252 32124
rect 37252 32068 37256 32124
rect 37192 32064 37256 32068
rect 2612 31580 2676 31584
rect 2612 31524 2616 31580
rect 2616 31524 2672 31580
rect 2672 31524 2676 31580
rect 2612 31520 2676 31524
rect 2692 31580 2756 31584
rect 2692 31524 2696 31580
rect 2696 31524 2752 31580
rect 2752 31524 2756 31580
rect 2692 31520 2756 31524
rect 2772 31580 2836 31584
rect 2772 31524 2776 31580
rect 2776 31524 2832 31580
rect 2832 31524 2836 31580
rect 2772 31520 2836 31524
rect 2852 31580 2916 31584
rect 2852 31524 2856 31580
rect 2856 31524 2912 31580
rect 2912 31524 2916 31580
rect 2852 31520 2916 31524
rect 7612 31580 7676 31584
rect 7612 31524 7616 31580
rect 7616 31524 7672 31580
rect 7672 31524 7676 31580
rect 7612 31520 7676 31524
rect 7692 31580 7756 31584
rect 7692 31524 7696 31580
rect 7696 31524 7752 31580
rect 7752 31524 7756 31580
rect 7692 31520 7756 31524
rect 7772 31580 7836 31584
rect 7772 31524 7776 31580
rect 7776 31524 7832 31580
rect 7832 31524 7836 31580
rect 7772 31520 7836 31524
rect 7852 31580 7916 31584
rect 7852 31524 7856 31580
rect 7856 31524 7912 31580
rect 7912 31524 7916 31580
rect 7852 31520 7916 31524
rect 12612 31580 12676 31584
rect 12612 31524 12616 31580
rect 12616 31524 12672 31580
rect 12672 31524 12676 31580
rect 12612 31520 12676 31524
rect 12692 31580 12756 31584
rect 12692 31524 12696 31580
rect 12696 31524 12752 31580
rect 12752 31524 12756 31580
rect 12692 31520 12756 31524
rect 12772 31580 12836 31584
rect 12772 31524 12776 31580
rect 12776 31524 12832 31580
rect 12832 31524 12836 31580
rect 12772 31520 12836 31524
rect 12852 31580 12916 31584
rect 12852 31524 12856 31580
rect 12856 31524 12912 31580
rect 12912 31524 12916 31580
rect 12852 31520 12916 31524
rect 17612 31580 17676 31584
rect 17612 31524 17616 31580
rect 17616 31524 17672 31580
rect 17672 31524 17676 31580
rect 17612 31520 17676 31524
rect 17692 31580 17756 31584
rect 17692 31524 17696 31580
rect 17696 31524 17752 31580
rect 17752 31524 17756 31580
rect 17692 31520 17756 31524
rect 17772 31580 17836 31584
rect 17772 31524 17776 31580
rect 17776 31524 17832 31580
rect 17832 31524 17836 31580
rect 17772 31520 17836 31524
rect 17852 31580 17916 31584
rect 17852 31524 17856 31580
rect 17856 31524 17912 31580
rect 17912 31524 17916 31580
rect 17852 31520 17916 31524
rect 22612 31580 22676 31584
rect 22612 31524 22616 31580
rect 22616 31524 22672 31580
rect 22672 31524 22676 31580
rect 22612 31520 22676 31524
rect 22692 31580 22756 31584
rect 22692 31524 22696 31580
rect 22696 31524 22752 31580
rect 22752 31524 22756 31580
rect 22692 31520 22756 31524
rect 22772 31580 22836 31584
rect 22772 31524 22776 31580
rect 22776 31524 22832 31580
rect 22832 31524 22836 31580
rect 22772 31520 22836 31524
rect 22852 31580 22916 31584
rect 22852 31524 22856 31580
rect 22856 31524 22912 31580
rect 22912 31524 22916 31580
rect 22852 31520 22916 31524
rect 27612 31580 27676 31584
rect 27612 31524 27616 31580
rect 27616 31524 27672 31580
rect 27672 31524 27676 31580
rect 27612 31520 27676 31524
rect 27692 31580 27756 31584
rect 27692 31524 27696 31580
rect 27696 31524 27752 31580
rect 27752 31524 27756 31580
rect 27692 31520 27756 31524
rect 27772 31580 27836 31584
rect 27772 31524 27776 31580
rect 27776 31524 27832 31580
rect 27832 31524 27836 31580
rect 27772 31520 27836 31524
rect 27852 31580 27916 31584
rect 27852 31524 27856 31580
rect 27856 31524 27912 31580
rect 27912 31524 27916 31580
rect 27852 31520 27916 31524
rect 32612 31580 32676 31584
rect 32612 31524 32616 31580
rect 32616 31524 32672 31580
rect 32672 31524 32676 31580
rect 32612 31520 32676 31524
rect 32692 31580 32756 31584
rect 32692 31524 32696 31580
rect 32696 31524 32752 31580
rect 32752 31524 32756 31580
rect 32692 31520 32756 31524
rect 32772 31580 32836 31584
rect 32772 31524 32776 31580
rect 32776 31524 32832 31580
rect 32832 31524 32836 31580
rect 32772 31520 32836 31524
rect 32852 31580 32916 31584
rect 32852 31524 32856 31580
rect 32856 31524 32912 31580
rect 32912 31524 32916 31580
rect 32852 31520 32916 31524
rect 37612 31580 37676 31584
rect 37612 31524 37616 31580
rect 37616 31524 37672 31580
rect 37672 31524 37676 31580
rect 37612 31520 37676 31524
rect 37692 31580 37756 31584
rect 37692 31524 37696 31580
rect 37696 31524 37752 31580
rect 37752 31524 37756 31580
rect 37692 31520 37756 31524
rect 37772 31580 37836 31584
rect 37772 31524 37776 31580
rect 37776 31524 37832 31580
rect 37832 31524 37836 31580
rect 37772 31520 37836 31524
rect 37852 31580 37916 31584
rect 37852 31524 37856 31580
rect 37856 31524 37912 31580
rect 37912 31524 37916 31580
rect 37852 31520 37916 31524
rect 30604 31180 30668 31244
rect 23244 31044 23308 31108
rect 1952 31036 2016 31040
rect 1952 30980 1956 31036
rect 1956 30980 2012 31036
rect 2012 30980 2016 31036
rect 1952 30976 2016 30980
rect 2032 31036 2096 31040
rect 2032 30980 2036 31036
rect 2036 30980 2092 31036
rect 2092 30980 2096 31036
rect 2032 30976 2096 30980
rect 2112 31036 2176 31040
rect 2112 30980 2116 31036
rect 2116 30980 2172 31036
rect 2172 30980 2176 31036
rect 2112 30976 2176 30980
rect 2192 31036 2256 31040
rect 2192 30980 2196 31036
rect 2196 30980 2252 31036
rect 2252 30980 2256 31036
rect 2192 30976 2256 30980
rect 6952 31036 7016 31040
rect 6952 30980 6956 31036
rect 6956 30980 7012 31036
rect 7012 30980 7016 31036
rect 6952 30976 7016 30980
rect 7032 31036 7096 31040
rect 7032 30980 7036 31036
rect 7036 30980 7092 31036
rect 7092 30980 7096 31036
rect 7032 30976 7096 30980
rect 7112 31036 7176 31040
rect 7112 30980 7116 31036
rect 7116 30980 7172 31036
rect 7172 30980 7176 31036
rect 7112 30976 7176 30980
rect 7192 31036 7256 31040
rect 7192 30980 7196 31036
rect 7196 30980 7252 31036
rect 7252 30980 7256 31036
rect 7192 30976 7256 30980
rect 11952 31036 12016 31040
rect 11952 30980 11956 31036
rect 11956 30980 12012 31036
rect 12012 30980 12016 31036
rect 11952 30976 12016 30980
rect 12032 31036 12096 31040
rect 12032 30980 12036 31036
rect 12036 30980 12092 31036
rect 12092 30980 12096 31036
rect 12032 30976 12096 30980
rect 12112 31036 12176 31040
rect 12112 30980 12116 31036
rect 12116 30980 12172 31036
rect 12172 30980 12176 31036
rect 12112 30976 12176 30980
rect 12192 31036 12256 31040
rect 12192 30980 12196 31036
rect 12196 30980 12252 31036
rect 12252 30980 12256 31036
rect 12192 30976 12256 30980
rect 16952 31036 17016 31040
rect 16952 30980 16956 31036
rect 16956 30980 17012 31036
rect 17012 30980 17016 31036
rect 16952 30976 17016 30980
rect 17032 31036 17096 31040
rect 17032 30980 17036 31036
rect 17036 30980 17092 31036
rect 17092 30980 17096 31036
rect 17032 30976 17096 30980
rect 17112 31036 17176 31040
rect 17112 30980 17116 31036
rect 17116 30980 17172 31036
rect 17172 30980 17176 31036
rect 17112 30976 17176 30980
rect 17192 31036 17256 31040
rect 17192 30980 17196 31036
rect 17196 30980 17252 31036
rect 17252 30980 17256 31036
rect 17192 30976 17256 30980
rect 21952 31036 22016 31040
rect 21952 30980 21956 31036
rect 21956 30980 22012 31036
rect 22012 30980 22016 31036
rect 21952 30976 22016 30980
rect 22032 31036 22096 31040
rect 22032 30980 22036 31036
rect 22036 30980 22092 31036
rect 22092 30980 22096 31036
rect 22032 30976 22096 30980
rect 22112 31036 22176 31040
rect 22112 30980 22116 31036
rect 22116 30980 22172 31036
rect 22172 30980 22176 31036
rect 22112 30976 22176 30980
rect 22192 31036 22256 31040
rect 22192 30980 22196 31036
rect 22196 30980 22252 31036
rect 22252 30980 22256 31036
rect 22192 30976 22256 30980
rect 26952 31036 27016 31040
rect 26952 30980 26956 31036
rect 26956 30980 27012 31036
rect 27012 30980 27016 31036
rect 26952 30976 27016 30980
rect 27032 31036 27096 31040
rect 27032 30980 27036 31036
rect 27036 30980 27092 31036
rect 27092 30980 27096 31036
rect 27032 30976 27096 30980
rect 27112 31036 27176 31040
rect 27112 30980 27116 31036
rect 27116 30980 27172 31036
rect 27172 30980 27176 31036
rect 27112 30976 27176 30980
rect 27192 31036 27256 31040
rect 27192 30980 27196 31036
rect 27196 30980 27252 31036
rect 27252 30980 27256 31036
rect 27192 30976 27256 30980
rect 31952 31036 32016 31040
rect 31952 30980 31956 31036
rect 31956 30980 32012 31036
rect 32012 30980 32016 31036
rect 31952 30976 32016 30980
rect 32032 31036 32096 31040
rect 32032 30980 32036 31036
rect 32036 30980 32092 31036
rect 32092 30980 32096 31036
rect 32032 30976 32096 30980
rect 32112 31036 32176 31040
rect 32112 30980 32116 31036
rect 32116 30980 32172 31036
rect 32172 30980 32176 31036
rect 32112 30976 32176 30980
rect 32192 31036 32256 31040
rect 32192 30980 32196 31036
rect 32196 30980 32252 31036
rect 32252 30980 32256 31036
rect 32192 30976 32256 30980
rect 36952 31036 37016 31040
rect 36952 30980 36956 31036
rect 36956 30980 37012 31036
rect 37012 30980 37016 31036
rect 36952 30976 37016 30980
rect 37032 31036 37096 31040
rect 37032 30980 37036 31036
rect 37036 30980 37092 31036
rect 37092 30980 37096 31036
rect 37032 30976 37096 30980
rect 37112 31036 37176 31040
rect 37112 30980 37116 31036
rect 37116 30980 37172 31036
rect 37172 30980 37176 31036
rect 37112 30976 37176 30980
rect 37192 31036 37256 31040
rect 37192 30980 37196 31036
rect 37196 30980 37252 31036
rect 37252 30980 37256 31036
rect 37192 30976 37256 30980
rect 2612 30492 2676 30496
rect 2612 30436 2616 30492
rect 2616 30436 2672 30492
rect 2672 30436 2676 30492
rect 2612 30432 2676 30436
rect 2692 30492 2756 30496
rect 2692 30436 2696 30492
rect 2696 30436 2752 30492
rect 2752 30436 2756 30492
rect 2692 30432 2756 30436
rect 2772 30492 2836 30496
rect 2772 30436 2776 30492
rect 2776 30436 2832 30492
rect 2832 30436 2836 30492
rect 2772 30432 2836 30436
rect 2852 30492 2916 30496
rect 2852 30436 2856 30492
rect 2856 30436 2912 30492
rect 2912 30436 2916 30492
rect 2852 30432 2916 30436
rect 7612 30492 7676 30496
rect 7612 30436 7616 30492
rect 7616 30436 7672 30492
rect 7672 30436 7676 30492
rect 7612 30432 7676 30436
rect 7692 30492 7756 30496
rect 7692 30436 7696 30492
rect 7696 30436 7752 30492
rect 7752 30436 7756 30492
rect 7692 30432 7756 30436
rect 7772 30492 7836 30496
rect 7772 30436 7776 30492
rect 7776 30436 7832 30492
rect 7832 30436 7836 30492
rect 7772 30432 7836 30436
rect 7852 30492 7916 30496
rect 7852 30436 7856 30492
rect 7856 30436 7912 30492
rect 7912 30436 7916 30492
rect 7852 30432 7916 30436
rect 12612 30492 12676 30496
rect 12612 30436 12616 30492
rect 12616 30436 12672 30492
rect 12672 30436 12676 30492
rect 12612 30432 12676 30436
rect 12692 30492 12756 30496
rect 12692 30436 12696 30492
rect 12696 30436 12752 30492
rect 12752 30436 12756 30492
rect 12692 30432 12756 30436
rect 12772 30492 12836 30496
rect 12772 30436 12776 30492
rect 12776 30436 12832 30492
rect 12832 30436 12836 30492
rect 12772 30432 12836 30436
rect 12852 30492 12916 30496
rect 12852 30436 12856 30492
rect 12856 30436 12912 30492
rect 12912 30436 12916 30492
rect 12852 30432 12916 30436
rect 17612 30492 17676 30496
rect 17612 30436 17616 30492
rect 17616 30436 17672 30492
rect 17672 30436 17676 30492
rect 17612 30432 17676 30436
rect 17692 30492 17756 30496
rect 17692 30436 17696 30492
rect 17696 30436 17752 30492
rect 17752 30436 17756 30492
rect 17692 30432 17756 30436
rect 17772 30492 17836 30496
rect 17772 30436 17776 30492
rect 17776 30436 17832 30492
rect 17832 30436 17836 30492
rect 17772 30432 17836 30436
rect 17852 30492 17916 30496
rect 17852 30436 17856 30492
rect 17856 30436 17912 30492
rect 17912 30436 17916 30492
rect 17852 30432 17916 30436
rect 22612 30492 22676 30496
rect 22612 30436 22616 30492
rect 22616 30436 22672 30492
rect 22672 30436 22676 30492
rect 22612 30432 22676 30436
rect 22692 30492 22756 30496
rect 22692 30436 22696 30492
rect 22696 30436 22752 30492
rect 22752 30436 22756 30492
rect 22692 30432 22756 30436
rect 22772 30492 22836 30496
rect 22772 30436 22776 30492
rect 22776 30436 22832 30492
rect 22832 30436 22836 30492
rect 22772 30432 22836 30436
rect 22852 30492 22916 30496
rect 22852 30436 22856 30492
rect 22856 30436 22912 30492
rect 22912 30436 22916 30492
rect 22852 30432 22916 30436
rect 27612 30492 27676 30496
rect 27612 30436 27616 30492
rect 27616 30436 27672 30492
rect 27672 30436 27676 30492
rect 27612 30432 27676 30436
rect 27692 30492 27756 30496
rect 27692 30436 27696 30492
rect 27696 30436 27752 30492
rect 27752 30436 27756 30492
rect 27692 30432 27756 30436
rect 27772 30492 27836 30496
rect 27772 30436 27776 30492
rect 27776 30436 27832 30492
rect 27832 30436 27836 30492
rect 27772 30432 27836 30436
rect 27852 30492 27916 30496
rect 27852 30436 27856 30492
rect 27856 30436 27912 30492
rect 27912 30436 27916 30492
rect 27852 30432 27916 30436
rect 32612 30492 32676 30496
rect 32612 30436 32616 30492
rect 32616 30436 32672 30492
rect 32672 30436 32676 30492
rect 32612 30432 32676 30436
rect 32692 30492 32756 30496
rect 32692 30436 32696 30492
rect 32696 30436 32752 30492
rect 32752 30436 32756 30492
rect 32692 30432 32756 30436
rect 32772 30492 32836 30496
rect 32772 30436 32776 30492
rect 32776 30436 32832 30492
rect 32832 30436 32836 30492
rect 32772 30432 32836 30436
rect 32852 30492 32916 30496
rect 32852 30436 32856 30492
rect 32856 30436 32912 30492
rect 32912 30436 32916 30492
rect 32852 30432 32916 30436
rect 37612 30492 37676 30496
rect 37612 30436 37616 30492
rect 37616 30436 37672 30492
rect 37672 30436 37676 30492
rect 37612 30432 37676 30436
rect 37692 30492 37756 30496
rect 37692 30436 37696 30492
rect 37696 30436 37752 30492
rect 37752 30436 37756 30492
rect 37692 30432 37756 30436
rect 37772 30492 37836 30496
rect 37772 30436 37776 30492
rect 37776 30436 37832 30492
rect 37832 30436 37836 30492
rect 37772 30432 37836 30436
rect 37852 30492 37916 30496
rect 37852 30436 37856 30492
rect 37856 30436 37912 30492
rect 37912 30436 37916 30492
rect 37852 30432 37916 30436
rect 1952 29948 2016 29952
rect 1952 29892 1956 29948
rect 1956 29892 2012 29948
rect 2012 29892 2016 29948
rect 1952 29888 2016 29892
rect 2032 29948 2096 29952
rect 2032 29892 2036 29948
rect 2036 29892 2092 29948
rect 2092 29892 2096 29948
rect 2032 29888 2096 29892
rect 2112 29948 2176 29952
rect 2112 29892 2116 29948
rect 2116 29892 2172 29948
rect 2172 29892 2176 29948
rect 2112 29888 2176 29892
rect 2192 29948 2256 29952
rect 2192 29892 2196 29948
rect 2196 29892 2252 29948
rect 2252 29892 2256 29948
rect 2192 29888 2256 29892
rect 6952 29948 7016 29952
rect 6952 29892 6956 29948
rect 6956 29892 7012 29948
rect 7012 29892 7016 29948
rect 6952 29888 7016 29892
rect 7032 29948 7096 29952
rect 7032 29892 7036 29948
rect 7036 29892 7092 29948
rect 7092 29892 7096 29948
rect 7032 29888 7096 29892
rect 7112 29948 7176 29952
rect 7112 29892 7116 29948
rect 7116 29892 7172 29948
rect 7172 29892 7176 29948
rect 7112 29888 7176 29892
rect 7192 29948 7256 29952
rect 7192 29892 7196 29948
rect 7196 29892 7252 29948
rect 7252 29892 7256 29948
rect 7192 29888 7256 29892
rect 11952 29948 12016 29952
rect 11952 29892 11956 29948
rect 11956 29892 12012 29948
rect 12012 29892 12016 29948
rect 11952 29888 12016 29892
rect 12032 29948 12096 29952
rect 12032 29892 12036 29948
rect 12036 29892 12092 29948
rect 12092 29892 12096 29948
rect 12032 29888 12096 29892
rect 12112 29948 12176 29952
rect 12112 29892 12116 29948
rect 12116 29892 12172 29948
rect 12172 29892 12176 29948
rect 12112 29888 12176 29892
rect 12192 29948 12256 29952
rect 12192 29892 12196 29948
rect 12196 29892 12252 29948
rect 12252 29892 12256 29948
rect 12192 29888 12256 29892
rect 16952 29948 17016 29952
rect 16952 29892 16956 29948
rect 16956 29892 17012 29948
rect 17012 29892 17016 29948
rect 16952 29888 17016 29892
rect 17032 29948 17096 29952
rect 17032 29892 17036 29948
rect 17036 29892 17092 29948
rect 17092 29892 17096 29948
rect 17032 29888 17096 29892
rect 17112 29948 17176 29952
rect 17112 29892 17116 29948
rect 17116 29892 17172 29948
rect 17172 29892 17176 29948
rect 17112 29888 17176 29892
rect 17192 29948 17256 29952
rect 17192 29892 17196 29948
rect 17196 29892 17252 29948
rect 17252 29892 17256 29948
rect 17192 29888 17256 29892
rect 21952 29948 22016 29952
rect 21952 29892 21956 29948
rect 21956 29892 22012 29948
rect 22012 29892 22016 29948
rect 21952 29888 22016 29892
rect 22032 29948 22096 29952
rect 22032 29892 22036 29948
rect 22036 29892 22092 29948
rect 22092 29892 22096 29948
rect 22032 29888 22096 29892
rect 22112 29948 22176 29952
rect 22112 29892 22116 29948
rect 22116 29892 22172 29948
rect 22172 29892 22176 29948
rect 22112 29888 22176 29892
rect 22192 29948 22256 29952
rect 22192 29892 22196 29948
rect 22196 29892 22252 29948
rect 22252 29892 22256 29948
rect 22192 29888 22256 29892
rect 26952 29948 27016 29952
rect 26952 29892 26956 29948
rect 26956 29892 27012 29948
rect 27012 29892 27016 29948
rect 26952 29888 27016 29892
rect 27032 29948 27096 29952
rect 27032 29892 27036 29948
rect 27036 29892 27092 29948
rect 27092 29892 27096 29948
rect 27032 29888 27096 29892
rect 27112 29948 27176 29952
rect 27112 29892 27116 29948
rect 27116 29892 27172 29948
rect 27172 29892 27176 29948
rect 27112 29888 27176 29892
rect 27192 29948 27256 29952
rect 27192 29892 27196 29948
rect 27196 29892 27252 29948
rect 27252 29892 27256 29948
rect 27192 29888 27256 29892
rect 31952 29948 32016 29952
rect 31952 29892 31956 29948
rect 31956 29892 32012 29948
rect 32012 29892 32016 29948
rect 31952 29888 32016 29892
rect 32032 29948 32096 29952
rect 32032 29892 32036 29948
rect 32036 29892 32092 29948
rect 32092 29892 32096 29948
rect 32032 29888 32096 29892
rect 32112 29948 32176 29952
rect 32112 29892 32116 29948
rect 32116 29892 32172 29948
rect 32172 29892 32176 29948
rect 32112 29888 32176 29892
rect 32192 29948 32256 29952
rect 32192 29892 32196 29948
rect 32196 29892 32252 29948
rect 32252 29892 32256 29948
rect 32192 29888 32256 29892
rect 36952 29948 37016 29952
rect 36952 29892 36956 29948
rect 36956 29892 37012 29948
rect 37012 29892 37016 29948
rect 36952 29888 37016 29892
rect 37032 29948 37096 29952
rect 37032 29892 37036 29948
rect 37036 29892 37092 29948
rect 37092 29892 37096 29948
rect 37032 29888 37096 29892
rect 37112 29948 37176 29952
rect 37112 29892 37116 29948
rect 37116 29892 37172 29948
rect 37172 29892 37176 29948
rect 37112 29888 37176 29892
rect 37192 29948 37256 29952
rect 37192 29892 37196 29948
rect 37196 29892 37252 29948
rect 37252 29892 37256 29948
rect 37192 29888 37256 29892
rect 2612 29404 2676 29408
rect 2612 29348 2616 29404
rect 2616 29348 2672 29404
rect 2672 29348 2676 29404
rect 2612 29344 2676 29348
rect 2692 29404 2756 29408
rect 2692 29348 2696 29404
rect 2696 29348 2752 29404
rect 2752 29348 2756 29404
rect 2692 29344 2756 29348
rect 2772 29404 2836 29408
rect 2772 29348 2776 29404
rect 2776 29348 2832 29404
rect 2832 29348 2836 29404
rect 2772 29344 2836 29348
rect 2852 29404 2916 29408
rect 2852 29348 2856 29404
rect 2856 29348 2912 29404
rect 2912 29348 2916 29404
rect 2852 29344 2916 29348
rect 7612 29404 7676 29408
rect 7612 29348 7616 29404
rect 7616 29348 7672 29404
rect 7672 29348 7676 29404
rect 7612 29344 7676 29348
rect 7692 29404 7756 29408
rect 7692 29348 7696 29404
rect 7696 29348 7752 29404
rect 7752 29348 7756 29404
rect 7692 29344 7756 29348
rect 7772 29404 7836 29408
rect 7772 29348 7776 29404
rect 7776 29348 7832 29404
rect 7832 29348 7836 29404
rect 7772 29344 7836 29348
rect 7852 29404 7916 29408
rect 7852 29348 7856 29404
rect 7856 29348 7912 29404
rect 7912 29348 7916 29404
rect 7852 29344 7916 29348
rect 12612 29404 12676 29408
rect 12612 29348 12616 29404
rect 12616 29348 12672 29404
rect 12672 29348 12676 29404
rect 12612 29344 12676 29348
rect 12692 29404 12756 29408
rect 12692 29348 12696 29404
rect 12696 29348 12752 29404
rect 12752 29348 12756 29404
rect 12692 29344 12756 29348
rect 12772 29404 12836 29408
rect 12772 29348 12776 29404
rect 12776 29348 12832 29404
rect 12832 29348 12836 29404
rect 12772 29344 12836 29348
rect 12852 29404 12916 29408
rect 12852 29348 12856 29404
rect 12856 29348 12912 29404
rect 12912 29348 12916 29404
rect 12852 29344 12916 29348
rect 17612 29404 17676 29408
rect 17612 29348 17616 29404
rect 17616 29348 17672 29404
rect 17672 29348 17676 29404
rect 17612 29344 17676 29348
rect 17692 29404 17756 29408
rect 17692 29348 17696 29404
rect 17696 29348 17752 29404
rect 17752 29348 17756 29404
rect 17692 29344 17756 29348
rect 17772 29404 17836 29408
rect 17772 29348 17776 29404
rect 17776 29348 17832 29404
rect 17832 29348 17836 29404
rect 17772 29344 17836 29348
rect 17852 29404 17916 29408
rect 17852 29348 17856 29404
rect 17856 29348 17912 29404
rect 17912 29348 17916 29404
rect 17852 29344 17916 29348
rect 22612 29404 22676 29408
rect 22612 29348 22616 29404
rect 22616 29348 22672 29404
rect 22672 29348 22676 29404
rect 22612 29344 22676 29348
rect 22692 29404 22756 29408
rect 22692 29348 22696 29404
rect 22696 29348 22752 29404
rect 22752 29348 22756 29404
rect 22692 29344 22756 29348
rect 22772 29404 22836 29408
rect 22772 29348 22776 29404
rect 22776 29348 22832 29404
rect 22832 29348 22836 29404
rect 22772 29344 22836 29348
rect 22852 29404 22916 29408
rect 22852 29348 22856 29404
rect 22856 29348 22912 29404
rect 22912 29348 22916 29404
rect 22852 29344 22916 29348
rect 27612 29404 27676 29408
rect 27612 29348 27616 29404
rect 27616 29348 27672 29404
rect 27672 29348 27676 29404
rect 27612 29344 27676 29348
rect 27692 29404 27756 29408
rect 27692 29348 27696 29404
rect 27696 29348 27752 29404
rect 27752 29348 27756 29404
rect 27692 29344 27756 29348
rect 27772 29404 27836 29408
rect 27772 29348 27776 29404
rect 27776 29348 27832 29404
rect 27832 29348 27836 29404
rect 27772 29344 27836 29348
rect 27852 29404 27916 29408
rect 27852 29348 27856 29404
rect 27856 29348 27912 29404
rect 27912 29348 27916 29404
rect 27852 29344 27916 29348
rect 32612 29404 32676 29408
rect 32612 29348 32616 29404
rect 32616 29348 32672 29404
rect 32672 29348 32676 29404
rect 32612 29344 32676 29348
rect 32692 29404 32756 29408
rect 32692 29348 32696 29404
rect 32696 29348 32752 29404
rect 32752 29348 32756 29404
rect 32692 29344 32756 29348
rect 32772 29404 32836 29408
rect 32772 29348 32776 29404
rect 32776 29348 32832 29404
rect 32832 29348 32836 29404
rect 32772 29344 32836 29348
rect 32852 29404 32916 29408
rect 32852 29348 32856 29404
rect 32856 29348 32912 29404
rect 32912 29348 32916 29404
rect 32852 29344 32916 29348
rect 37612 29404 37676 29408
rect 37612 29348 37616 29404
rect 37616 29348 37672 29404
rect 37672 29348 37676 29404
rect 37612 29344 37676 29348
rect 37692 29404 37756 29408
rect 37692 29348 37696 29404
rect 37696 29348 37752 29404
rect 37752 29348 37756 29404
rect 37692 29344 37756 29348
rect 37772 29404 37836 29408
rect 37772 29348 37776 29404
rect 37776 29348 37832 29404
rect 37832 29348 37836 29404
rect 37772 29344 37836 29348
rect 37852 29404 37916 29408
rect 37852 29348 37856 29404
rect 37856 29348 37912 29404
rect 37912 29348 37916 29404
rect 37852 29344 37916 29348
rect 1952 28860 2016 28864
rect 1952 28804 1956 28860
rect 1956 28804 2012 28860
rect 2012 28804 2016 28860
rect 1952 28800 2016 28804
rect 2032 28860 2096 28864
rect 2032 28804 2036 28860
rect 2036 28804 2092 28860
rect 2092 28804 2096 28860
rect 2032 28800 2096 28804
rect 2112 28860 2176 28864
rect 2112 28804 2116 28860
rect 2116 28804 2172 28860
rect 2172 28804 2176 28860
rect 2112 28800 2176 28804
rect 2192 28860 2256 28864
rect 2192 28804 2196 28860
rect 2196 28804 2252 28860
rect 2252 28804 2256 28860
rect 2192 28800 2256 28804
rect 6952 28860 7016 28864
rect 6952 28804 6956 28860
rect 6956 28804 7012 28860
rect 7012 28804 7016 28860
rect 6952 28800 7016 28804
rect 7032 28860 7096 28864
rect 7032 28804 7036 28860
rect 7036 28804 7092 28860
rect 7092 28804 7096 28860
rect 7032 28800 7096 28804
rect 7112 28860 7176 28864
rect 7112 28804 7116 28860
rect 7116 28804 7172 28860
rect 7172 28804 7176 28860
rect 7112 28800 7176 28804
rect 7192 28860 7256 28864
rect 7192 28804 7196 28860
rect 7196 28804 7252 28860
rect 7252 28804 7256 28860
rect 7192 28800 7256 28804
rect 11952 28860 12016 28864
rect 11952 28804 11956 28860
rect 11956 28804 12012 28860
rect 12012 28804 12016 28860
rect 11952 28800 12016 28804
rect 12032 28860 12096 28864
rect 12032 28804 12036 28860
rect 12036 28804 12092 28860
rect 12092 28804 12096 28860
rect 12032 28800 12096 28804
rect 12112 28860 12176 28864
rect 12112 28804 12116 28860
rect 12116 28804 12172 28860
rect 12172 28804 12176 28860
rect 12112 28800 12176 28804
rect 12192 28860 12256 28864
rect 12192 28804 12196 28860
rect 12196 28804 12252 28860
rect 12252 28804 12256 28860
rect 12192 28800 12256 28804
rect 16952 28860 17016 28864
rect 16952 28804 16956 28860
rect 16956 28804 17012 28860
rect 17012 28804 17016 28860
rect 16952 28800 17016 28804
rect 17032 28860 17096 28864
rect 17032 28804 17036 28860
rect 17036 28804 17092 28860
rect 17092 28804 17096 28860
rect 17032 28800 17096 28804
rect 17112 28860 17176 28864
rect 17112 28804 17116 28860
rect 17116 28804 17172 28860
rect 17172 28804 17176 28860
rect 17112 28800 17176 28804
rect 17192 28860 17256 28864
rect 17192 28804 17196 28860
rect 17196 28804 17252 28860
rect 17252 28804 17256 28860
rect 17192 28800 17256 28804
rect 21952 28860 22016 28864
rect 21952 28804 21956 28860
rect 21956 28804 22012 28860
rect 22012 28804 22016 28860
rect 21952 28800 22016 28804
rect 22032 28860 22096 28864
rect 22032 28804 22036 28860
rect 22036 28804 22092 28860
rect 22092 28804 22096 28860
rect 22032 28800 22096 28804
rect 22112 28860 22176 28864
rect 22112 28804 22116 28860
rect 22116 28804 22172 28860
rect 22172 28804 22176 28860
rect 22112 28800 22176 28804
rect 22192 28860 22256 28864
rect 22192 28804 22196 28860
rect 22196 28804 22252 28860
rect 22252 28804 22256 28860
rect 22192 28800 22256 28804
rect 26952 28860 27016 28864
rect 26952 28804 26956 28860
rect 26956 28804 27012 28860
rect 27012 28804 27016 28860
rect 26952 28800 27016 28804
rect 27032 28860 27096 28864
rect 27032 28804 27036 28860
rect 27036 28804 27092 28860
rect 27092 28804 27096 28860
rect 27032 28800 27096 28804
rect 27112 28860 27176 28864
rect 27112 28804 27116 28860
rect 27116 28804 27172 28860
rect 27172 28804 27176 28860
rect 27112 28800 27176 28804
rect 27192 28860 27256 28864
rect 27192 28804 27196 28860
rect 27196 28804 27252 28860
rect 27252 28804 27256 28860
rect 27192 28800 27256 28804
rect 31952 28860 32016 28864
rect 31952 28804 31956 28860
rect 31956 28804 32012 28860
rect 32012 28804 32016 28860
rect 31952 28800 32016 28804
rect 32032 28860 32096 28864
rect 32032 28804 32036 28860
rect 32036 28804 32092 28860
rect 32092 28804 32096 28860
rect 32032 28800 32096 28804
rect 32112 28860 32176 28864
rect 32112 28804 32116 28860
rect 32116 28804 32172 28860
rect 32172 28804 32176 28860
rect 32112 28800 32176 28804
rect 32192 28860 32256 28864
rect 32192 28804 32196 28860
rect 32196 28804 32252 28860
rect 32252 28804 32256 28860
rect 32192 28800 32256 28804
rect 36952 28860 37016 28864
rect 36952 28804 36956 28860
rect 36956 28804 37012 28860
rect 37012 28804 37016 28860
rect 36952 28800 37016 28804
rect 37032 28860 37096 28864
rect 37032 28804 37036 28860
rect 37036 28804 37092 28860
rect 37092 28804 37096 28860
rect 37032 28800 37096 28804
rect 37112 28860 37176 28864
rect 37112 28804 37116 28860
rect 37116 28804 37172 28860
rect 37172 28804 37176 28860
rect 37112 28800 37176 28804
rect 37192 28860 37256 28864
rect 37192 28804 37196 28860
rect 37196 28804 37252 28860
rect 37252 28804 37256 28860
rect 37192 28800 37256 28804
rect 2612 28316 2676 28320
rect 2612 28260 2616 28316
rect 2616 28260 2672 28316
rect 2672 28260 2676 28316
rect 2612 28256 2676 28260
rect 2692 28316 2756 28320
rect 2692 28260 2696 28316
rect 2696 28260 2752 28316
rect 2752 28260 2756 28316
rect 2692 28256 2756 28260
rect 2772 28316 2836 28320
rect 2772 28260 2776 28316
rect 2776 28260 2832 28316
rect 2832 28260 2836 28316
rect 2772 28256 2836 28260
rect 2852 28316 2916 28320
rect 2852 28260 2856 28316
rect 2856 28260 2912 28316
rect 2912 28260 2916 28316
rect 2852 28256 2916 28260
rect 7612 28316 7676 28320
rect 7612 28260 7616 28316
rect 7616 28260 7672 28316
rect 7672 28260 7676 28316
rect 7612 28256 7676 28260
rect 7692 28316 7756 28320
rect 7692 28260 7696 28316
rect 7696 28260 7752 28316
rect 7752 28260 7756 28316
rect 7692 28256 7756 28260
rect 7772 28316 7836 28320
rect 7772 28260 7776 28316
rect 7776 28260 7832 28316
rect 7832 28260 7836 28316
rect 7772 28256 7836 28260
rect 7852 28316 7916 28320
rect 7852 28260 7856 28316
rect 7856 28260 7912 28316
rect 7912 28260 7916 28316
rect 7852 28256 7916 28260
rect 12612 28316 12676 28320
rect 12612 28260 12616 28316
rect 12616 28260 12672 28316
rect 12672 28260 12676 28316
rect 12612 28256 12676 28260
rect 12692 28316 12756 28320
rect 12692 28260 12696 28316
rect 12696 28260 12752 28316
rect 12752 28260 12756 28316
rect 12692 28256 12756 28260
rect 12772 28316 12836 28320
rect 12772 28260 12776 28316
rect 12776 28260 12832 28316
rect 12832 28260 12836 28316
rect 12772 28256 12836 28260
rect 12852 28316 12916 28320
rect 12852 28260 12856 28316
rect 12856 28260 12912 28316
rect 12912 28260 12916 28316
rect 12852 28256 12916 28260
rect 17612 28316 17676 28320
rect 17612 28260 17616 28316
rect 17616 28260 17672 28316
rect 17672 28260 17676 28316
rect 17612 28256 17676 28260
rect 17692 28316 17756 28320
rect 17692 28260 17696 28316
rect 17696 28260 17752 28316
rect 17752 28260 17756 28316
rect 17692 28256 17756 28260
rect 17772 28316 17836 28320
rect 17772 28260 17776 28316
rect 17776 28260 17832 28316
rect 17832 28260 17836 28316
rect 17772 28256 17836 28260
rect 17852 28316 17916 28320
rect 17852 28260 17856 28316
rect 17856 28260 17912 28316
rect 17912 28260 17916 28316
rect 17852 28256 17916 28260
rect 22612 28316 22676 28320
rect 22612 28260 22616 28316
rect 22616 28260 22672 28316
rect 22672 28260 22676 28316
rect 22612 28256 22676 28260
rect 22692 28316 22756 28320
rect 22692 28260 22696 28316
rect 22696 28260 22752 28316
rect 22752 28260 22756 28316
rect 22692 28256 22756 28260
rect 22772 28316 22836 28320
rect 22772 28260 22776 28316
rect 22776 28260 22832 28316
rect 22832 28260 22836 28316
rect 22772 28256 22836 28260
rect 22852 28316 22916 28320
rect 22852 28260 22856 28316
rect 22856 28260 22912 28316
rect 22912 28260 22916 28316
rect 22852 28256 22916 28260
rect 27612 28316 27676 28320
rect 27612 28260 27616 28316
rect 27616 28260 27672 28316
rect 27672 28260 27676 28316
rect 27612 28256 27676 28260
rect 27692 28316 27756 28320
rect 27692 28260 27696 28316
rect 27696 28260 27752 28316
rect 27752 28260 27756 28316
rect 27692 28256 27756 28260
rect 27772 28316 27836 28320
rect 27772 28260 27776 28316
rect 27776 28260 27832 28316
rect 27832 28260 27836 28316
rect 27772 28256 27836 28260
rect 27852 28316 27916 28320
rect 27852 28260 27856 28316
rect 27856 28260 27912 28316
rect 27912 28260 27916 28316
rect 27852 28256 27916 28260
rect 32612 28316 32676 28320
rect 32612 28260 32616 28316
rect 32616 28260 32672 28316
rect 32672 28260 32676 28316
rect 32612 28256 32676 28260
rect 32692 28316 32756 28320
rect 32692 28260 32696 28316
rect 32696 28260 32752 28316
rect 32752 28260 32756 28316
rect 32692 28256 32756 28260
rect 32772 28316 32836 28320
rect 32772 28260 32776 28316
rect 32776 28260 32832 28316
rect 32832 28260 32836 28316
rect 32772 28256 32836 28260
rect 32852 28316 32916 28320
rect 32852 28260 32856 28316
rect 32856 28260 32912 28316
rect 32912 28260 32916 28316
rect 32852 28256 32916 28260
rect 37612 28316 37676 28320
rect 37612 28260 37616 28316
rect 37616 28260 37672 28316
rect 37672 28260 37676 28316
rect 37612 28256 37676 28260
rect 37692 28316 37756 28320
rect 37692 28260 37696 28316
rect 37696 28260 37752 28316
rect 37752 28260 37756 28316
rect 37692 28256 37756 28260
rect 37772 28316 37836 28320
rect 37772 28260 37776 28316
rect 37776 28260 37832 28316
rect 37832 28260 37836 28316
rect 37772 28256 37836 28260
rect 37852 28316 37916 28320
rect 37852 28260 37856 28316
rect 37856 28260 37912 28316
rect 37912 28260 37916 28316
rect 37852 28256 37916 28260
rect 1952 27772 2016 27776
rect 1952 27716 1956 27772
rect 1956 27716 2012 27772
rect 2012 27716 2016 27772
rect 1952 27712 2016 27716
rect 2032 27772 2096 27776
rect 2032 27716 2036 27772
rect 2036 27716 2092 27772
rect 2092 27716 2096 27772
rect 2032 27712 2096 27716
rect 2112 27772 2176 27776
rect 2112 27716 2116 27772
rect 2116 27716 2172 27772
rect 2172 27716 2176 27772
rect 2112 27712 2176 27716
rect 2192 27772 2256 27776
rect 2192 27716 2196 27772
rect 2196 27716 2252 27772
rect 2252 27716 2256 27772
rect 2192 27712 2256 27716
rect 6952 27772 7016 27776
rect 6952 27716 6956 27772
rect 6956 27716 7012 27772
rect 7012 27716 7016 27772
rect 6952 27712 7016 27716
rect 7032 27772 7096 27776
rect 7032 27716 7036 27772
rect 7036 27716 7092 27772
rect 7092 27716 7096 27772
rect 7032 27712 7096 27716
rect 7112 27772 7176 27776
rect 7112 27716 7116 27772
rect 7116 27716 7172 27772
rect 7172 27716 7176 27772
rect 7112 27712 7176 27716
rect 7192 27772 7256 27776
rect 7192 27716 7196 27772
rect 7196 27716 7252 27772
rect 7252 27716 7256 27772
rect 7192 27712 7256 27716
rect 11952 27772 12016 27776
rect 11952 27716 11956 27772
rect 11956 27716 12012 27772
rect 12012 27716 12016 27772
rect 11952 27712 12016 27716
rect 12032 27772 12096 27776
rect 12032 27716 12036 27772
rect 12036 27716 12092 27772
rect 12092 27716 12096 27772
rect 12032 27712 12096 27716
rect 12112 27772 12176 27776
rect 12112 27716 12116 27772
rect 12116 27716 12172 27772
rect 12172 27716 12176 27772
rect 12112 27712 12176 27716
rect 12192 27772 12256 27776
rect 12192 27716 12196 27772
rect 12196 27716 12252 27772
rect 12252 27716 12256 27772
rect 12192 27712 12256 27716
rect 16952 27772 17016 27776
rect 16952 27716 16956 27772
rect 16956 27716 17012 27772
rect 17012 27716 17016 27772
rect 16952 27712 17016 27716
rect 17032 27772 17096 27776
rect 17032 27716 17036 27772
rect 17036 27716 17092 27772
rect 17092 27716 17096 27772
rect 17032 27712 17096 27716
rect 17112 27772 17176 27776
rect 17112 27716 17116 27772
rect 17116 27716 17172 27772
rect 17172 27716 17176 27772
rect 17112 27712 17176 27716
rect 17192 27772 17256 27776
rect 17192 27716 17196 27772
rect 17196 27716 17252 27772
rect 17252 27716 17256 27772
rect 17192 27712 17256 27716
rect 21952 27772 22016 27776
rect 21952 27716 21956 27772
rect 21956 27716 22012 27772
rect 22012 27716 22016 27772
rect 21952 27712 22016 27716
rect 22032 27772 22096 27776
rect 22032 27716 22036 27772
rect 22036 27716 22092 27772
rect 22092 27716 22096 27772
rect 22032 27712 22096 27716
rect 22112 27772 22176 27776
rect 22112 27716 22116 27772
rect 22116 27716 22172 27772
rect 22172 27716 22176 27772
rect 22112 27712 22176 27716
rect 22192 27772 22256 27776
rect 22192 27716 22196 27772
rect 22196 27716 22252 27772
rect 22252 27716 22256 27772
rect 22192 27712 22256 27716
rect 26952 27772 27016 27776
rect 26952 27716 26956 27772
rect 26956 27716 27012 27772
rect 27012 27716 27016 27772
rect 26952 27712 27016 27716
rect 27032 27772 27096 27776
rect 27032 27716 27036 27772
rect 27036 27716 27092 27772
rect 27092 27716 27096 27772
rect 27032 27712 27096 27716
rect 27112 27772 27176 27776
rect 27112 27716 27116 27772
rect 27116 27716 27172 27772
rect 27172 27716 27176 27772
rect 27112 27712 27176 27716
rect 27192 27772 27256 27776
rect 27192 27716 27196 27772
rect 27196 27716 27252 27772
rect 27252 27716 27256 27772
rect 27192 27712 27256 27716
rect 31952 27772 32016 27776
rect 31952 27716 31956 27772
rect 31956 27716 32012 27772
rect 32012 27716 32016 27772
rect 31952 27712 32016 27716
rect 32032 27772 32096 27776
rect 32032 27716 32036 27772
rect 32036 27716 32092 27772
rect 32092 27716 32096 27772
rect 32032 27712 32096 27716
rect 32112 27772 32176 27776
rect 32112 27716 32116 27772
rect 32116 27716 32172 27772
rect 32172 27716 32176 27772
rect 32112 27712 32176 27716
rect 32192 27772 32256 27776
rect 32192 27716 32196 27772
rect 32196 27716 32252 27772
rect 32252 27716 32256 27772
rect 32192 27712 32256 27716
rect 36952 27772 37016 27776
rect 36952 27716 36956 27772
rect 36956 27716 37012 27772
rect 37012 27716 37016 27772
rect 36952 27712 37016 27716
rect 37032 27772 37096 27776
rect 37032 27716 37036 27772
rect 37036 27716 37092 27772
rect 37092 27716 37096 27772
rect 37032 27712 37096 27716
rect 37112 27772 37176 27776
rect 37112 27716 37116 27772
rect 37116 27716 37172 27772
rect 37172 27716 37176 27772
rect 37112 27712 37176 27716
rect 37192 27772 37256 27776
rect 37192 27716 37196 27772
rect 37196 27716 37252 27772
rect 37252 27716 37256 27772
rect 37192 27712 37256 27716
rect 2612 27228 2676 27232
rect 2612 27172 2616 27228
rect 2616 27172 2672 27228
rect 2672 27172 2676 27228
rect 2612 27168 2676 27172
rect 2692 27228 2756 27232
rect 2692 27172 2696 27228
rect 2696 27172 2752 27228
rect 2752 27172 2756 27228
rect 2692 27168 2756 27172
rect 2772 27228 2836 27232
rect 2772 27172 2776 27228
rect 2776 27172 2832 27228
rect 2832 27172 2836 27228
rect 2772 27168 2836 27172
rect 2852 27228 2916 27232
rect 2852 27172 2856 27228
rect 2856 27172 2912 27228
rect 2912 27172 2916 27228
rect 2852 27168 2916 27172
rect 7612 27228 7676 27232
rect 7612 27172 7616 27228
rect 7616 27172 7672 27228
rect 7672 27172 7676 27228
rect 7612 27168 7676 27172
rect 7692 27228 7756 27232
rect 7692 27172 7696 27228
rect 7696 27172 7752 27228
rect 7752 27172 7756 27228
rect 7692 27168 7756 27172
rect 7772 27228 7836 27232
rect 7772 27172 7776 27228
rect 7776 27172 7832 27228
rect 7832 27172 7836 27228
rect 7772 27168 7836 27172
rect 7852 27228 7916 27232
rect 7852 27172 7856 27228
rect 7856 27172 7912 27228
rect 7912 27172 7916 27228
rect 7852 27168 7916 27172
rect 12612 27228 12676 27232
rect 12612 27172 12616 27228
rect 12616 27172 12672 27228
rect 12672 27172 12676 27228
rect 12612 27168 12676 27172
rect 12692 27228 12756 27232
rect 12692 27172 12696 27228
rect 12696 27172 12752 27228
rect 12752 27172 12756 27228
rect 12692 27168 12756 27172
rect 12772 27228 12836 27232
rect 12772 27172 12776 27228
rect 12776 27172 12832 27228
rect 12832 27172 12836 27228
rect 12772 27168 12836 27172
rect 12852 27228 12916 27232
rect 12852 27172 12856 27228
rect 12856 27172 12912 27228
rect 12912 27172 12916 27228
rect 12852 27168 12916 27172
rect 17612 27228 17676 27232
rect 17612 27172 17616 27228
rect 17616 27172 17672 27228
rect 17672 27172 17676 27228
rect 17612 27168 17676 27172
rect 17692 27228 17756 27232
rect 17692 27172 17696 27228
rect 17696 27172 17752 27228
rect 17752 27172 17756 27228
rect 17692 27168 17756 27172
rect 17772 27228 17836 27232
rect 17772 27172 17776 27228
rect 17776 27172 17832 27228
rect 17832 27172 17836 27228
rect 17772 27168 17836 27172
rect 17852 27228 17916 27232
rect 17852 27172 17856 27228
rect 17856 27172 17912 27228
rect 17912 27172 17916 27228
rect 17852 27168 17916 27172
rect 22612 27228 22676 27232
rect 22612 27172 22616 27228
rect 22616 27172 22672 27228
rect 22672 27172 22676 27228
rect 22612 27168 22676 27172
rect 22692 27228 22756 27232
rect 22692 27172 22696 27228
rect 22696 27172 22752 27228
rect 22752 27172 22756 27228
rect 22692 27168 22756 27172
rect 22772 27228 22836 27232
rect 22772 27172 22776 27228
rect 22776 27172 22832 27228
rect 22832 27172 22836 27228
rect 22772 27168 22836 27172
rect 22852 27228 22916 27232
rect 22852 27172 22856 27228
rect 22856 27172 22912 27228
rect 22912 27172 22916 27228
rect 22852 27168 22916 27172
rect 27612 27228 27676 27232
rect 27612 27172 27616 27228
rect 27616 27172 27672 27228
rect 27672 27172 27676 27228
rect 27612 27168 27676 27172
rect 27692 27228 27756 27232
rect 27692 27172 27696 27228
rect 27696 27172 27752 27228
rect 27752 27172 27756 27228
rect 27692 27168 27756 27172
rect 27772 27228 27836 27232
rect 27772 27172 27776 27228
rect 27776 27172 27832 27228
rect 27832 27172 27836 27228
rect 27772 27168 27836 27172
rect 27852 27228 27916 27232
rect 27852 27172 27856 27228
rect 27856 27172 27912 27228
rect 27912 27172 27916 27228
rect 27852 27168 27916 27172
rect 32612 27228 32676 27232
rect 32612 27172 32616 27228
rect 32616 27172 32672 27228
rect 32672 27172 32676 27228
rect 32612 27168 32676 27172
rect 32692 27228 32756 27232
rect 32692 27172 32696 27228
rect 32696 27172 32752 27228
rect 32752 27172 32756 27228
rect 32692 27168 32756 27172
rect 32772 27228 32836 27232
rect 32772 27172 32776 27228
rect 32776 27172 32832 27228
rect 32832 27172 32836 27228
rect 32772 27168 32836 27172
rect 32852 27228 32916 27232
rect 32852 27172 32856 27228
rect 32856 27172 32912 27228
rect 32912 27172 32916 27228
rect 32852 27168 32916 27172
rect 37612 27228 37676 27232
rect 37612 27172 37616 27228
rect 37616 27172 37672 27228
rect 37672 27172 37676 27228
rect 37612 27168 37676 27172
rect 37692 27228 37756 27232
rect 37692 27172 37696 27228
rect 37696 27172 37752 27228
rect 37752 27172 37756 27228
rect 37692 27168 37756 27172
rect 37772 27228 37836 27232
rect 37772 27172 37776 27228
rect 37776 27172 37832 27228
rect 37832 27172 37836 27228
rect 37772 27168 37836 27172
rect 37852 27228 37916 27232
rect 37852 27172 37856 27228
rect 37856 27172 37912 27228
rect 37912 27172 37916 27228
rect 37852 27168 37916 27172
rect 1952 26684 2016 26688
rect 1952 26628 1956 26684
rect 1956 26628 2012 26684
rect 2012 26628 2016 26684
rect 1952 26624 2016 26628
rect 2032 26684 2096 26688
rect 2032 26628 2036 26684
rect 2036 26628 2092 26684
rect 2092 26628 2096 26684
rect 2032 26624 2096 26628
rect 2112 26684 2176 26688
rect 2112 26628 2116 26684
rect 2116 26628 2172 26684
rect 2172 26628 2176 26684
rect 2112 26624 2176 26628
rect 2192 26684 2256 26688
rect 2192 26628 2196 26684
rect 2196 26628 2252 26684
rect 2252 26628 2256 26684
rect 2192 26624 2256 26628
rect 6952 26684 7016 26688
rect 6952 26628 6956 26684
rect 6956 26628 7012 26684
rect 7012 26628 7016 26684
rect 6952 26624 7016 26628
rect 7032 26684 7096 26688
rect 7032 26628 7036 26684
rect 7036 26628 7092 26684
rect 7092 26628 7096 26684
rect 7032 26624 7096 26628
rect 7112 26684 7176 26688
rect 7112 26628 7116 26684
rect 7116 26628 7172 26684
rect 7172 26628 7176 26684
rect 7112 26624 7176 26628
rect 7192 26684 7256 26688
rect 7192 26628 7196 26684
rect 7196 26628 7252 26684
rect 7252 26628 7256 26684
rect 7192 26624 7256 26628
rect 11952 26684 12016 26688
rect 11952 26628 11956 26684
rect 11956 26628 12012 26684
rect 12012 26628 12016 26684
rect 11952 26624 12016 26628
rect 12032 26684 12096 26688
rect 12032 26628 12036 26684
rect 12036 26628 12092 26684
rect 12092 26628 12096 26684
rect 12032 26624 12096 26628
rect 12112 26684 12176 26688
rect 12112 26628 12116 26684
rect 12116 26628 12172 26684
rect 12172 26628 12176 26684
rect 12112 26624 12176 26628
rect 12192 26684 12256 26688
rect 12192 26628 12196 26684
rect 12196 26628 12252 26684
rect 12252 26628 12256 26684
rect 12192 26624 12256 26628
rect 16952 26684 17016 26688
rect 16952 26628 16956 26684
rect 16956 26628 17012 26684
rect 17012 26628 17016 26684
rect 16952 26624 17016 26628
rect 17032 26684 17096 26688
rect 17032 26628 17036 26684
rect 17036 26628 17092 26684
rect 17092 26628 17096 26684
rect 17032 26624 17096 26628
rect 17112 26684 17176 26688
rect 17112 26628 17116 26684
rect 17116 26628 17172 26684
rect 17172 26628 17176 26684
rect 17112 26624 17176 26628
rect 17192 26684 17256 26688
rect 17192 26628 17196 26684
rect 17196 26628 17252 26684
rect 17252 26628 17256 26684
rect 17192 26624 17256 26628
rect 21952 26684 22016 26688
rect 21952 26628 21956 26684
rect 21956 26628 22012 26684
rect 22012 26628 22016 26684
rect 21952 26624 22016 26628
rect 22032 26684 22096 26688
rect 22032 26628 22036 26684
rect 22036 26628 22092 26684
rect 22092 26628 22096 26684
rect 22032 26624 22096 26628
rect 22112 26684 22176 26688
rect 22112 26628 22116 26684
rect 22116 26628 22172 26684
rect 22172 26628 22176 26684
rect 22112 26624 22176 26628
rect 22192 26684 22256 26688
rect 22192 26628 22196 26684
rect 22196 26628 22252 26684
rect 22252 26628 22256 26684
rect 22192 26624 22256 26628
rect 26952 26684 27016 26688
rect 26952 26628 26956 26684
rect 26956 26628 27012 26684
rect 27012 26628 27016 26684
rect 26952 26624 27016 26628
rect 27032 26684 27096 26688
rect 27032 26628 27036 26684
rect 27036 26628 27092 26684
rect 27092 26628 27096 26684
rect 27032 26624 27096 26628
rect 27112 26684 27176 26688
rect 27112 26628 27116 26684
rect 27116 26628 27172 26684
rect 27172 26628 27176 26684
rect 27112 26624 27176 26628
rect 27192 26684 27256 26688
rect 27192 26628 27196 26684
rect 27196 26628 27252 26684
rect 27252 26628 27256 26684
rect 27192 26624 27256 26628
rect 31952 26684 32016 26688
rect 31952 26628 31956 26684
rect 31956 26628 32012 26684
rect 32012 26628 32016 26684
rect 31952 26624 32016 26628
rect 32032 26684 32096 26688
rect 32032 26628 32036 26684
rect 32036 26628 32092 26684
rect 32092 26628 32096 26684
rect 32032 26624 32096 26628
rect 32112 26684 32176 26688
rect 32112 26628 32116 26684
rect 32116 26628 32172 26684
rect 32172 26628 32176 26684
rect 32112 26624 32176 26628
rect 32192 26684 32256 26688
rect 32192 26628 32196 26684
rect 32196 26628 32252 26684
rect 32252 26628 32256 26684
rect 32192 26624 32256 26628
rect 36952 26684 37016 26688
rect 36952 26628 36956 26684
rect 36956 26628 37012 26684
rect 37012 26628 37016 26684
rect 36952 26624 37016 26628
rect 37032 26684 37096 26688
rect 37032 26628 37036 26684
rect 37036 26628 37092 26684
rect 37092 26628 37096 26684
rect 37032 26624 37096 26628
rect 37112 26684 37176 26688
rect 37112 26628 37116 26684
rect 37116 26628 37172 26684
rect 37172 26628 37176 26684
rect 37112 26624 37176 26628
rect 37192 26684 37256 26688
rect 37192 26628 37196 26684
rect 37196 26628 37252 26684
rect 37252 26628 37256 26684
rect 37192 26624 37256 26628
rect 18460 26284 18524 26348
rect 2612 26140 2676 26144
rect 2612 26084 2616 26140
rect 2616 26084 2672 26140
rect 2672 26084 2676 26140
rect 2612 26080 2676 26084
rect 2692 26140 2756 26144
rect 2692 26084 2696 26140
rect 2696 26084 2752 26140
rect 2752 26084 2756 26140
rect 2692 26080 2756 26084
rect 2772 26140 2836 26144
rect 2772 26084 2776 26140
rect 2776 26084 2832 26140
rect 2832 26084 2836 26140
rect 2772 26080 2836 26084
rect 2852 26140 2916 26144
rect 2852 26084 2856 26140
rect 2856 26084 2912 26140
rect 2912 26084 2916 26140
rect 2852 26080 2916 26084
rect 7612 26140 7676 26144
rect 7612 26084 7616 26140
rect 7616 26084 7672 26140
rect 7672 26084 7676 26140
rect 7612 26080 7676 26084
rect 7692 26140 7756 26144
rect 7692 26084 7696 26140
rect 7696 26084 7752 26140
rect 7752 26084 7756 26140
rect 7692 26080 7756 26084
rect 7772 26140 7836 26144
rect 7772 26084 7776 26140
rect 7776 26084 7832 26140
rect 7832 26084 7836 26140
rect 7772 26080 7836 26084
rect 7852 26140 7916 26144
rect 7852 26084 7856 26140
rect 7856 26084 7912 26140
rect 7912 26084 7916 26140
rect 7852 26080 7916 26084
rect 12612 26140 12676 26144
rect 12612 26084 12616 26140
rect 12616 26084 12672 26140
rect 12672 26084 12676 26140
rect 12612 26080 12676 26084
rect 12692 26140 12756 26144
rect 12692 26084 12696 26140
rect 12696 26084 12752 26140
rect 12752 26084 12756 26140
rect 12692 26080 12756 26084
rect 12772 26140 12836 26144
rect 12772 26084 12776 26140
rect 12776 26084 12832 26140
rect 12832 26084 12836 26140
rect 12772 26080 12836 26084
rect 12852 26140 12916 26144
rect 12852 26084 12856 26140
rect 12856 26084 12912 26140
rect 12912 26084 12916 26140
rect 12852 26080 12916 26084
rect 17612 26140 17676 26144
rect 17612 26084 17616 26140
rect 17616 26084 17672 26140
rect 17672 26084 17676 26140
rect 17612 26080 17676 26084
rect 17692 26140 17756 26144
rect 17692 26084 17696 26140
rect 17696 26084 17752 26140
rect 17752 26084 17756 26140
rect 17692 26080 17756 26084
rect 17772 26140 17836 26144
rect 17772 26084 17776 26140
rect 17776 26084 17832 26140
rect 17832 26084 17836 26140
rect 17772 26080 17836 26084
rect 17852 26140 17916 26144
rect 17852 26084 17856 26140
rect 17856 26084 17912 26140
rect 17912 26084 17916 26140
rect 17852 26080 17916 26084
rect 22612 26140 22676 26144
rect 22612 26084 22616 26140
rect 22616 26084 22672 26140
rect 22672 26084 22676 26140
rect 22612 26080 22676 26084
rect 22692 26140 22756 26144
rect 22692 26084 22696 26140
rect 22696 26084 22752 26140
rect 22752 26084 22756 26140
rect 22692 26080 22756 26084
rect 22772 26140 22836 26144
rect 22772 26084 22776 26140
rect 22776 26084 22832 26140
rect 22832 26084 22836 26140
rect 22772 26080 22836 26084
rect 22852 26140 22916 26144
rect 22852 26084 22856 26140
rect 22856 26084 22912 26140
rect 22912 26084 22916 26140
rect 22852 26080 22916 26084
rect 27612 26140 27676 26144
rect 27612 26084 27616 26140
rect 27616 26084 27672 26140
rect 27672 26084 27676 26140
rect 27612 26080 27676 26084
rect 27692 26140 27756 26144
rect 27692 26084 27696 26140
rect 27696 26084 27752 26140
rect 27752 26084 27756 26140
rect 27692 26080 27756 26084
rect 27772 26140 27836 26144
rect 27772 26084 27776 26140
rect 27776 26084 27832 26140
rect 27832 26084 27836 26140
rect 27772 26080 27836 26084
rect 27852 26140 27916 26144
rect 27852 26084 27856 26140
rect 27856 26084 27912 26140
rect 27912 26084 27916 26140
rect 27852 26080 27916 26084
rect 32612 26140 32676 26144
rect 32612 26084 32616 26140
rect 32616 26084 32672 26140
rect 32672 26084 32676 26140
rect 32612 26080 32676 26084
rect 32692 26140 32756 26144
rect 32692 26084 32696 26140
rect 32696 26084 32752 26140
rect 32752 26084 32756 26140
rect 32692 26080 32756 26084
rect 32772 26140 32836 26144
rect 32772 26084 32776 26140
rect 32776 26084 32832 26140
rect 32832 26084 32836 26140
rect 32772 26080 32836 26084
rect 32852 26140 32916 26144
rect 32852 26084 32856 26140
rect 32856 26084 32912 26140
rect 32912 26084 32916 26140
rect 32852 26080 32916 26084
rect 37612 26140 37676 26144
rect 37612 26084 37616 26140
rect 37616 26084 37672 26140
rect 37672 26084 37676 26140
rect 37612 26080 37676 26084
rect 37692 26140 37756 26144
rect 37692 26084 37696 26140
rect 37696 26084 37752 26140
rect 37752 26084 37756 26140
rect 37692 26080 37756 26084
rect 37772 26140 37836 26144
rect 37772 26084 37776 26140
rect 37776 26084 37832 26140
rect 37832 26084 37836 26140
rect 37772 26080 37836 26084
rect 37852 26140 37916 26144
rect 37852 26084 37856 26140
rect 37856 26084 37912 26140
rect 37912 26084 37916 26140
rect 37852 26080 37916 26084
rect 1952 25596 2016 25600
rect 1952 25540 1956 25596
rect 1956 25540 2012 25596
rect 2012 25540 2016 25596
rect 1952 25536 2016 25540
rect 2032 25596 2096 25600
rect 2032 25540 2036 25596
rect 2036 25540 2092 25596
rect 2092 25540 2096 25596
rect 2032 25536 2096 25540
rect 2112 25596 2176 25600
rect 2112 25540 2116 25596
rect 2116 25540 2172 25596
rect 2172 25540 2176 25596
rect 2112 25536 2176 25540
rect 2192 25596 2256 25600
rect 2192 25540 2196 25596
rect 2196 25540 2252 25596
rect 2252 25540 2256 25596
rect 2192 25536 2256 25540
rect 6952 25596 7016 25600
rect 6952 25540 6956 25596
rect 6956 25540 7012 25596
rect 7012 25540 7016 25596
rect 6952 25536 7016 25540
rect 7032 25596 7096 25600
rect 7032 25540 7036 25596
rect 7036 25540 7092 25596
rect 7092 25540 7096 25596
rect 7032 25536 7096 25540
rect 7112 25596 7176 25600
rect 7112 25540 7116 25596
rect 7116 25540 7172 25596
rect 7172 25540 7176 25596
rect 7112 25536 7176 25540
rect 7192 25596 7256 25600
rect 7192 25540 7196 25596
rect 7196 25540 7252 25596
rect 7252 25540 7256 25596
rect 7192 25536 7256 25540
rect 11952 25596 12016 25600
rect 11952 25540 11956 25596
rect 11956 25540 12012 25596
rect 12012 25540 12016 25596
rect 11952 25536 12016 25540
rect 12032 25596 12096 25600
rect 12032 25540 12036 25596
rect 12036 25540 12092 25596
rect 12092 25540 12096 25596
rect 12032 25536 12096 25540
rect 12112 25596 12176 25600
rect 12112 25540 12116 25596
rect 12116 25540 12172 25596
rect 12172 25540 12176 25596
rect 12112 25536 12176 25540
rect 12192 25596 12256 25600
rect 12192 25540 12196 25596
rect 12196 25540 12252 25596
rect 12252 25540 12256 25596
rect 12192 25536 12256 25540
rect 16952 25596 17016 25600
rect 16952 25540 16956 25596
rect 16956 25540 17012 25596
rect 17012 25540 17016 25596
rect 16952 25536 17016 25540
rect 17032 25596 17096 25600
rect 17032 25540 17036 25596
rect 17036 25540 17092 25596
rect 17092 25540 17096 25596
rect 17032 25536 17096 25540
rect 17112 25596 17176 25600
rect 17112 25540 17116 25596
rect 17116 25540 17172 25596
rect 17172 25540 17176 25596
rect 17112 25536 17176 25540
rect 17192 25596 17256 25600
rect 17192 25540 17196 25596
rect 17196 25540 17252 25596
rect 17252 25540 17256 25596
rect 17192 25536 17256 25540
rect 21952 25596 22016 25600
rect 21952 25540 21956 25596
rect 21956 25540 22012 25596
rect 22012 25540 22016 25596
rect 21952 25536 22016 25540
rect 22032 25596 22096 25600
rect 22032 25540 22036 25596
rect 22036 25540 22092 25596
rect 22092 25540 22096 25596
rect 22032 25536 22096 25540
rect 22112 25596 22176 25600
rect 22112 25540 22116 25596
rect 22116 25540 22172 25596
rect 22172 25540 22176 25596
rect 22112 25536 22176 25540
rect 22192 25596 22256 25600
rect 22192 25540 22196 25596
rect 22196 25540 22252 25596
rect 22252 25540 22256 25596
rect 22192 25536 22256 25540
rect 26952 25596 27016 25600
rect 26952 25540 26956 25596
rect 26956 25540 27012 25596
rect 27012 25540 27016 25596
rect 26952 25536 27016 25540
rect 27032 25596 27096 25600
rect 27032 25540 27036 25596
rect 27036 25540 27092 25596
rect 27092 25540 27096 25596
rect 27032 25536 27096 25540
rect 27112 25596 27176 25600
rect 27112 25540 27116 25596
rect 27116 25540 27172 25596
rect 27172 25540 27176 25596
rect 27112 25536 27176 25540
rect 27192 25596 27256 25600
rect 27192 25540 27196 25596
rect 27196 25540 27252 25596
rect 27252 25540 27256 25596
rect 27192 25536 27256 25540
rect 31952 25596 32016 25600
rect 31952 25540 31956 25596
rect 31956 25540 32012 25596
rect 32012 25540 32016 25596
rect 31952 25536 32016 25540
rect 32032 25596 32096 25600
rect 32032 25540 32036 25596
rect 32036 25540 32092 25596
rect 32092 25540 32096 25596
rect 32032 25536 32096 25540
rect 32112 25596 32176 25600
rect 32112 25540 32116 25596
rect 32116 25540 32172 25596
rect 32172 25540 32176 25596
rect 32112 25536 32176 25540
rect 32192 25596 32256 25600
rect 32192 25540 32196 25596
rect 32196 25540 32252 25596
rect 32252 25540 32256 25596
rect 32192 25536 32256 25540
rect 36952 25596 37016 25600
rect 36952 25540 36956 25596
rect 36956 25540 37012 25596
rect 37012 25540 37016 25596
rect 36952 25536 37016 25540
rect 37032 25596 37096 25600
rect 37032 25540 37036 25596
rect 37036 25540 37092 25596
rect 37092 25540 37096 25596
rect 37032 25536 37096 25540
rect 37112 25596 37176 25600
rect 37112 25540 37116 25596
rect 37116 25540 37172 25596
rect 37172 25540 37176 25596
rect 37112 25536 37176 25540
rect 37192 25596 37256 25600
rect 37192 25540 37196 25596
rect 37196 25540 37252 25596
rect 37252 25540 37256 25596
rect 37192 25536 37256 25540
rect 2612 25052 2676 25056
rect 2612 24996 2616 25052
rect 2616 24996 2672 25052
rect 2672 24996 2676 25052
rect 2612 24992 2676 24996
rect 2692 25052 2756 25056
rect 2692 24996 2696 25052
rect 2696 24996 2752 25052
rect 2752 24996 2756 25052
rect 2692 24992 2756 24996
rect 2772 25052 2836 25056
rect 2772 24996 2776 25052
rect 2776 24996 2832 25052
rect 2832 24996 2836 25052
rect 2772 24992 2836 24996
rect 2852 25052 2916 25056
rect 2852 24996 2856 25052
rect 2856 24996 2912 25052
rect 2912 24996 2916 25052
rect 2852 24992 2916 24996
rect 7612 25052 7676 25056
rect 7612 24996 7616 25052
rect 7616 24996 7672 25052
rect 7672 24996 7676 25052
rect 7612 24992 7676 24996
rect 7692 25052 7756 25056
rect 7692 24996 7696 25052
rect 7696 24996 7752 25052
rect 7752 24996 7756 25052
rect 7692 24992 7756 24996
rect 7772 25052 7836 25056
rect 7772 24996 7776 25052
rect 7776 24996 7832 25052
rect 7832 24996 7836 25052
rect 7772 24992 7836 24996
rect 7852 25052 7916 25056
rect 7852 24996 7856 25052
rect 7856 24996 7912 25052
rect 7912 24996 7916 25052
rect 7852 24992 7916 24996
rect 12612 25052 12676 25056
rect 12612 24996 12616 25052
rect 12616 24996 12672 25052
rect 12672 24996 12676 25052
rect 12612 24992 12676 24996
rect 12692 25052 12756 25056
rect 12692 24996 12696 25052
rect 12696 24996 12752 25052
rect 12752 24996 12756 25052
rect 12692 24992 12756 24996
rect 12772 25052 12836 25056
rect 12772 24996 12776 25052
rect 12776 24996 12832 25052
rect 12832 24996 12836 25052
rect 12772 24992 12836 24996
rect 12852 25052 12916 25056
rect 12852 24996 12856 25052
rect 12856 24996 12912 25052
rect 12912 24996 12916 25052
rect 12852 24992 12916 24996
rect 17612 25052 17676 25056
rect 17612 24996 17616 25052
rect 17616 24996 17672 25052
rect 17672 24996 17676 25052
rect 17612 24992 17676 24996
rect 17692 25052 17756 25056
rect 17692 24996 17696 25052
rect 17696 24996 17752 25052
rect 17752 24996 17756 25052
rect 17692 24992 17756 24996
rect 17772 25052 17836 25056
rect 17772 24996 17776 25052
rect 17776 24996 17832 25052
rect 17832 24996 17836 25052
rect 17772 24992 17836 24996
rect 17852 25052 17916 25056
rect 17852 24996 17856 25052
rect 17856 24996 17912 25052
rect 17912 24996 17916 25052
rect 17852 24992 17916 24996
rect 22612 25052 22676 25056
rect 22612 24996 22616 25052
rect 22616 24996 22672 25052
rect 22672 24996 22676 25052
rect 22612 24992 22676 24996
rect 22692 25052 22756 25056
rect 22692 24996 22696 25052
rect 22696 24996 22752 25052
rect 22752 24996 22756 25052
rect 22692 24992 22756 24996
rect 22772 25052 22836 25056
rect 22772 24996 22776 25052
rect 22776 24996 22832 25052
rect 22832 24996 22836 25052
rect 22772 24992 22836 24996
rect 22852 25052 22916 25056
rect 22852 24996 22856 25052
rect 22856 24996 22912 25052
rect 22912 24996 22916 25052
rect 22852 24992 22916 24996
rect 27612 25052 27676 25056
rect 27612 24996 27616 25052
rect 27616 24996 27672 25052
rect 27672 24996 27676 25052
rect 27612 24992 27676 24996
rect 27692 25052 27756 25056
rect 27692 24996 27696 25052
rect 27696 24996 27752 25052
rect 27752 24996 27756 25052
rect 27692 24992 27756 24996
rect 27772 25052 27836 25056
rect 27772 24996 27776 25052
rect 27776 24996 27832 25052
rect 27832 24996 27836 25052
rect 27772 24992 27836 24996
rect 27852 25052 27916 25056
rect 27852 24996 27856 25052
rect 27856 24996 27912 25052
rect 27912 24996 27916 25052
rect 27852 24992 27916 24996
rect 32612 25052 32676 25056
rect 32612 24996 32616 25052
rect 32616 24996 32672 25052
rect 32672 24996 32676 25052
rect 32612 24992 32676 24996
rect 32692 25052 32756 25056
rect 32692 24996 32696 25052
rect 32696 24996 32752 25052
rect 32752 24996 32756 25052
rect 32692 24992 32756 24996
rect 32772 25052 32836 25056
rect 32772 24996 32776 25052
rect 32776 24996 32832 25052
rect 32832 24996 32836 25052
rect 32772 24992 32836 24996
rect 32852 25052 32916 25056
rect 32852 24996 32856 25052
rect 32856 24996 32912 25052
rect 32912 24996 32916 25052
rect 32852 24992 32916 24996
rect 37612 25052 37676 25056
rect 37612 24996 37616 25052
rect 37616 24996 37672 25052
rect 37672 24996 37676 25052
rect 37612 24992 37676 24996
rect 37692 25052 37756 25056
rect 37692 24996 37696 25052
rect 37696 24996 37752 25052
rect 37752 24996 37756 25052
rect 37692 24992 37756 24996
rect 37772 25052 37836 25056
rect 37772 24996 37776 25052
rect 37776 24996 37832 25052
rect 37832 24996 37836 25052
rect 37772 24992 37836 24996
rect 37852 25052 37916 25056
rect 37852 24996 37856 25052
rect 37856 24996 37912 25052
rect 37912 24996 37916 25052
rect 37852 24992 37916 24996
rect 1952 24508 2016 24512
rect 1952 24452 1956 24508
rect 1956 24452 2012 24508
rect 2012 24452 2016 24508
rect 1952 24448 2016 24452
rect 2032 24508 2096 24512
rect 2032 24452 2036 24508
rect 2036 24452 2092 24508
rect 2092 24452 2096 24508
rect 2032 24448 2096 24452
rect 2112 24508 2176 24512
rect 2112 24452 2116 24508
rect 2116 24452 2172 24508
rect 2172 24452 2176 24508
rect 2112 24448 2176 24452
rect 2192 24508 2256 24512
rect 2192 24452 2196 24508
rect 2196 24452 2252 24508
rect 2252 24452 2256 24508
rect 2192 24448 2256 24452
rect 6952 24508 7016 24512
rect 6952 24452 6956 24508
rect 6956 24452 7012 24508
rect 7012 24452 7016 24508
rect 6952 24448 7016 24452
rect 7032 24508 7096 24512
rect 7032 24452 7036 24508
rect 7036 24452 7092 24508
rect 7092 24452 7096 24508
rect 7032 24448 7096 24452
rect 7112 24508 7176 24512
rect 7112 24452 7116 24508
rect 7116 24452 7172 24508
rect 7172 24452 7176 24508
rect 7112 24448 7176 24452
rect 7192 24508 7256 24512
rect 7192 24452 7196 24508
rect 7196 24452 7252 24508
rect 7252 24452 7256 24508
rect 7192 24448 7256 24452
rect 11952 24508 12016 24512
rect 11952 24452 11956 24508
rect 11956 24452 12012 24508
rect 12012 24452 12016 24508
rect 11952 24448 12016 24452
rect 12032 24508 12096 24512
rect 12032 24452 12036 24508
rect 12036 24452 12092 24508
rect 12092 24452 12096 24508
rect 12032 24448 12096 24452
rect 12112 24508 12176 24512
rect 12112 24452 12116 24508
rect 12116 24452 12172 24508
rect 12172 24452 12176 24508
rect 12112 24448 12176 24452
rect 12192 24508 12256 24512
rect 12192 24452 12196 24508
rect 12196 24452 12252 24508
rect 12252 24452 12256 24508
rect 12192 24448 12256 24452
rect 16952 24508 17016 24512
rect 16952 24452 16956 24508
rect 16956 24452 17012 24508
rect 17012 24452 17016 24508
rect 16952 24448 17016 24452
rect 17032 24508 17096 24512
rect 17032 24452 17036 24508
rect 17036 24452 17092 24508
rect 17092 24452 17096 24508
rect 17032 24448 17096 24452
rect 17112 24508 17176 24512
rect 17112 24452 17116 24508
rect 17116 24452 17172 24508
rect 17172 24452 17176 24508
rect 17112 24448 17176 24452
rect 17192 24508 17256 24512
rect 17192 24452 17196 24508
rect 17196 24452 17252 24508
rect 17252 24452 17256 24508
rect 17192 24448 17256 24452
rect 21952 24508 22016 24512
rect 21952 24452 21956 24508
rect 21956 24452 22012 24508
rect 22012 24452 22016 24508
rect 21952 24448 22016 24452
rect 22032 24508 22096 24512
rect 22032 24452 22036 24508
rect 22036 24452 22092 24508
rect 22092 24452 22096 24508
rect 22032 24448 22096 24452
rect 22112 24508 22176 24512
rect 22112 24452 22116 24508
rect 22116 24452 22172 24508
rect 22172 24452 22176 24508
rect 22112 24448 22176 24452
rect 22192 24508 22256 24512
rect 22192 24452 22196 24508
rect 22196 24452 22252 24508
rect 22252 24452 22256 24508
rect 22192 24448 22256 24452
rect 26952 24508 27016 24512
rect 26952 24452 26956 24508
rect 26956 24452 27012 24508
rect 27012 24452 27016 24508
rect 26952 24448 27016 24452
rect 27032 24508 27096 24512
rect 27032 24452 27036 24508
rect 27036 24452 27092 24508
rect 27092 24452 27096 24508
rect 27032 24448 27096 24452
rect 27112 24508 27176 24512
rect 27112 24452 27116 24508
rect 27116 24452 27172 24508
rect 27172 24452 27176 24508
rect 27112 24448 27176 24452
rect 27192 24508 27256 24512
rect 27192 24452 27196 24508
rect 27196 24452 27252 24508
rect 27252 24452 27256 24508
rect 27192 24448 27256 24452
rect 31952 24508 32016 24512
rect 31952 24452 31956 24508
rect 31956 24452 32012 24508
rect 32012 24452 32016 24508
rect 31952 24448 32016 24452
rect 32032 24508 32096 24512
rect 32032 24452 32036 24508
rect 32036 24452 32092 24508
rect 32092 24452 32096 24508
rect 32032 24448 32096 24452
rect 32112 24508 32176 24512
rect 32112 24452 32116 24508
rect 32116 24452 32172 24508
rect 32172 24452 32176 24508
rect 32112 24448 32176 24452
rect 32192 24508 32256 24512
rect 32192 24452 32196 24508
rect 32196 24452 32252 24508
rect 32252 24452 32256 24508
rect 32192 24448 32256 24452
rect 36952 24508 37016 24512
rect 36952 24452 36956 24508
rect 36956 24452 37012 24508
rect 37012 24452 37016 24508
rect 36952 24448 37016 24452
rect 37032 24508 37096 24512
rect 37032 24452 37036 24508
rect 37036 24452 37092 24508
rect 37092 24452 37096 24508
rect 37032 24448 37096 24452
rect 37112 24508 37176 24512
rect 37112 24452 37116 24508
rect 37116 24452 37172 24508
rect 37172 24452 37176 24508
rect 37112 24448 37176 24452
rect 37192 24508 37256 24512
rect 37192 24452 37196 24508
rect 37196 24452 37252 24508
rect 37252 24452 37256 24508
rect 37192 24448 37256 24452
rect 2612 23964 2676 23968
rect 2612 23908 2616 23964
rect 2616 23908 2672 23964
rect 2672 23908 2676 23964
rect 2612 23904 2676 23908
rect 2692 23964 2756 23968
rect 2692 23908 2696 23964
rect 2696 23908 2752 23964
rect 2752 23908 2756 23964
rect 2692 23904 2756 23908
rect 2772 23964 2836 23968
rect 2772 23908 2776 23964
rect 2776 23908 2832 23964
rect 2832 23908 2836 23964
rect 2772 23904 2836 23908
rect 2852 23964 2916 23968
rect 2852 23908 2856 23964
rect 2856 23908 2912 23964
rect 2912 23908 2916 23964
rect 2852 23904 2916 23908
rect 7612 23964 7676 23968
rect 7612 23908 7616 23964
rect 7616 23908 7672 23964
rect 7672 23908 7676 23964
rect 7612 23904 7676 23908
rect 7692 23964 7756 23968
rect 7692 23908 7696 23964
rect 7696 23908 7752 23964
rect 7752 23908 7756 23964
rect 7692 23904 7756 23908
rect 7772 23964 7836 23968
rect 7772 23908 7776 23964
rect 7776 23908 7832 23964
rect 7832 23908 7836 23964
rect 7772 23904 7836 23908
rect 7852 23964 7916 23968
rect 7852 23908 7856 23964
rect 7856 23908 7912 23964
rect 7912 23908 7916 23964
rect 7852 23904 7916 23908
rect 12612 23964 12676 23968
rect 12612 23908 12616 23964
rect 12616 23908 12672 23964
rect 12672 23908 12676 23964
rect 12612 23904 12676 23908
rect 12692 23964 12756 23968
rect 12692 23908 12696 23964
rect 12696 23908 12752 23964
rect 12752 23908 12756 23964
rect 12692 23904 12756 23908
rect 12772 23964 12836 23968
rect 12772 23908 12776 23964
rect 12776 23908 12832 23964
rect 12832 23908 12836 23964
rect 12772 23904 12836 23908
rect 12852 23964 12916 23968
rect 12852 23908 12856 23964
rect 12856 23908 12912 23964
rect 12912 23908 12916 23964
rect 12852 23904 12916 23908
rect 17612 23964 17676 23968
rect 17612 23908 17616 23964
rect 17616 23908 17672 23964
rect 17672 23908 17676 23964
rect 17612 23904 17676 23908
rect 17692 23964 17756 23968
rect 17692 23908 17696 23964
rect 17696 23908 17752 23964
rect 17752 23908 17756 23964
rect 17692 23904 17756 23908
rect 17772 23964 17836 23968
rect 17772 23908 17776 23964
rect 17776 23908 17832 23964
rect 17832 23908 17836 23964
rect 17772 23904 17836 23908
rect 17852 23964 17916 23968
rect 17852 23908 17856 23964
rect 17856 23908 17912 23964
rect 17912 23908 17916 23964
rect 17852 23904 17916 23908
rect 22612 23964 22676 23968
rect 22612 23908 22616 23964
rect 22616 23908 22672 23964
rect 22672 23908 22676 23964
rect 22612 23904 22676 23908
rect 22692 23964 22756 23968
rect 22692 23908 22696 23964
rect 22696 23908 22752 23964
rect 22752 23908 22756 23964
rect 22692 23904 22756 23908
rect 22772 23964 22836 23968
rect 22772 23908 22776 23964
rect 22776 23908 22832 23964
rect 22832 23908 22836 23964
rect 22772 23904 22836 23908
rect 22852 23964 22916 23968
rect 22852 23908 22856 23964
rect 22856 23908 22912 23964
rect 22912 23908 22916 23964
rect 22852 23904 22916 23908
rect 27612 23964 27676 23968
rect 27612 23908 27616 23964
rect 27616 23908 27672 23964
rect 27672 23908 27676 23964
rect 27612 23904 27676 23908
rect 27692 23964 27756 23968
rect 27692 23908 27696 23964
rect 27696 23908 27752 23964
rect 27752 23908 27756 23964
rect 27692 23904 27756 23908
rect 27772 23964 27836 23968
rect 27772 23908 27776 23964
rect 27776 23908 27832 23964
rect 27832 23908 27836 23964
rect 27772 23904 27836 23908
rect 27852 23964 27916 23968
rect 27852 23908 27856 23964
rect 27856 23908 27912 23964
rect 27912 23908 27916 23964
rect 27852 23904 27916 23908
rect 32612 23964 32676 23968
rect 32612 23908 32616 23964
rect 32616 23908 32672 23964
rect 32672 23908 32676 23964
rect 32612 23904 32676 23908
rect 32692 23964 32756 23968
rect 32692 23908 32696 23964
rect 32696 23908 32752 23964
rect 32752 23908 32756 23964
rect 32692 23904 32756 23908
rect 32772 23964 32836 23968
rect 32772 23908 32776 23964
rect 32776 23908 32832 23964
rect 32832 23908 32836 23964
rect 32772 23904 32836 23908
rect 32852 23964 32916 23968
rect 32852 23908 32856 23964
rect 32856 23908 32912 23964
rect 32912 23908 32916 23964
rect 32852 23904 32916 23908
rect 37612 23964 37676 23968
rect 37612 23908 37616 23964
rect 37616 23908 37672 23964
rect 37672 23908 37676 23964
rect 37612 23904 37676 23908
rect 37692 23964 37756 23968
rect 37692 23908 37696 23964
rect 37696 23908 37752 23964
rect 37752 23908 37756 23964
rect 37692 23904 37756 23908
rect 37772 23964 37836 23968
rect 37772 23908 37776 23964
rect 37776 23908 37832 23964
rect 37832 23908 37836 23964
rect 37772 23904 37836 23908
rect 37852 23964 37916 23968
rect 37852 23908 37856 23964
rect 37856 23908 37912 23964
rect 37912 23908 37916 23964
rect 37852 23904 37916 23908
rect 1952 23420 2016 23424
rect 1952 23364 1956 23420
rect 1956 23364 2012 23420
rect 2012 23364 2016 23420
rect 1952 23360 2016 23364
rect 2032 23420 2096 23424
rect 2032 23364 2036 23420
rect 2036 23364 2092 23420
rect 2092 23364 2096 23420
rect 2032 23360 2096 23364
rect 2112 23420 2176 23424
rect 2112 23364 2116 23420
rect 2116 23364 2172 23420
rect 2172 23364 2176 23420
rect 2112 23360 2176 23364
rect 2192 23420 2256 23424
rect 2192 23364 2196 23420
rect 2196 23364 2252 23420
rect 2252 23364 2256 23420
rect 2192 23360 2256 23364
rect 6952 23420 7016 23424
rect 6952 23364 6956 23420
rect 6956 23364 7012 23420
rect 7012 23364 7016 23420
rect 6952 23360 7016 23364
rect 7032 23420 7096 23424
rect 7032 23364 7036 23420
rect 7036 23364 7092 23420
rect 7092 23364 7096 23420
rect 7032 23360 7096 23364
rect 7112 23420 7176 23424
rect 7112 23364 7116 23420
rect 7116 23364 7172 23420
rect 7172 23364 7176 23420
rect 7112 23360 7176 23364
rect 7192 23420 7256 23424
rect 7192 23364 7196 23420
rect 7196 23364 7252 23420
rect 7252 23364 7256 23420
rect 7192 23360 7256 23364
rect 11952 23420 12016 23424
rect 11952 23364 11956 23420
rect 11956 23364 12012 23420
rect 12012 23364 12016 23420
rect 11952 23360 12016 23364
rect 12032 23420 12096 23424
rect 12032 23364 12036 23420
rect 12036 23364 12092 23420
rect 12092 23364 12096 23420
rect 12032 23360 12096 23364
rect 12112 23420 12176 23424
rect 12112 23364 12116 23420
rect 12116 23364 12172 23420
rect 12172 23364 12176 23420
rect 12112 23360 12176 23364
rect 12192 23420 12256 23424
rect 12192 23364 12196 23420
rect 12196 23364 12252 23420
rect 12252 23364 12256 23420
rect 12192 23360 12256 23364
rect 16952 23420 17016 23424
rect 16952 23364 16956 23420
rect 16956 23364 17012 23420
rect 17012 23364 17016 23420
rect 16952 23360 17016 23364
rect 17032 23420 17096 23424
rect 17032 23364 17036 23420
rect 17036 23364 17092 23420
rect 17092 23364 17096 23420
rect 17032 23360 17096 23364
rect 17112 23420 17176 23424
rect 17112 23364 17116 23420
rect 17116 23364 17172 23420
rect 17172 23364 17176 23420
rect 17112 23360 17176 23364
rect 17192 23420 17256 23424
rect 17192 23364 17196 23420
rect 17196 23364 17252 23420
rect 17252 23364 17256 23420
rect 17192 23360 17256 23364
rect 21952 23420 22016 23424
rect 21952 23364 21956 23420
rect 21956 23364 22012 23420
rect 22012 23364 22016 23420
rect 21952 23360 22016 23364
rect 22032 23420 22096 23424
rect 22032 23364 22036 23420
rect 22036 23364 22092 23420
rect 22092 23364 22096 23420
rect 22032 23360 22096 23364
rect 22112 23420 22176 23424
rect 22112 23364 22116 23420
rect 22116 23364 22172 23420
rect 22172 23364 22176 23420
rect 22112 23360 22176 23364
rect 22192 23420 22256 23424
rect 22192 23364 22196 23420
rect 22196 23364 22252 23420
rect 22252 23364 22256 23420
rect 22192 23360 22256 23364
rect 26952 23420 27016 23424
rect 26952 23364 26956 23420
rect 26956 23364 27012 23420
rect 27012 23364 27016 23420
rect 26952 23360 27016 23364
rect 27032 23420 27096 23424
rect 27032 23364 27036 23420
rect 27036 23364 27092 23420
rect 27092 23364 27096 23420
rect 27032 23360 27096 23364
rect 27112 23420 27176 23424
rect 27112 23364 27116 23420
rect 27116 23364 27172 23420
rect 27172 23364 27176 23420
rect 27112 23360 27176 23364
rect 27192 23420 27256 23424
rect 27192 23364 27196 23420
rect 27196 23364 27252 23420
rect 27252 23364 27256 23420
rect 27192 23360 27256 23364
rect 31952 23420 32016 23424
rect 31952 23364 31956 23420
rect 31956 23364 32012 23420
rect 32012 23364 32016 23420
rect 31952 23360 32016 23364
rect 32032 23420 32096 23424
rect 32032 23364 32036 23420
rect 32036 23364 32092 23420
rect 32092 23364 32096 23420
rect 32032 23360 32096 23364
rect 32112 23420 32176 23424
rect 32112 23364 32116 23420
rect 32116 23364 32172 23420
rect 32172 23364 32176 23420
rect 32112 23360 32176 23364
rect 32192 23420 32256 23424
rect 32192 23364 32196 23420
rect 32196 23364 32252 23420
rect 32252 23364 32256 23420
rect 32192 23360 32256 23364
rect 36952 23420 37016 23424
rect 36952 23364 36956 23420
rect 36956 23364 37012 23420
rect 37012 23364 37016 23420
rect 36952 23360 37016 23364
rect 37032 23420 37096 23424
rect 37032 23364 37036 23420
rect 37036 23364 37092 23420
rect 37092 23364 37096 23420
rect 37032 23360 37096 23364
rect 37112 23420 37176 23424
rect 37112 23364 37116 23420
rect 37116 23364 37172 23420
rect 37172 23364 37176 23420
rect 37112 23360 37176 23364
rect 37192 23420 37256 23424
rect 37192 23364 37196 23420
rect 37196 23364 37252 23420
rect 37252 23364 37256 23420
rect 37192 23360 37256 23364
rect 2612 22876 2676 22880
rect 2612 22820 2616 22876
rect 2616 22820 2672 22876
rect 2672 22820 2676 22876
rect 2612 22816 2676 22820
rect 2692 22876 2756 22880
rect 2692 22820 2696 22876
rect 2696 22820 2752 22876
rect 2752 22820 2756 22876
rect 2692 22816 2756 22820
rect 2772 22876 2836 22880
rect 2772 22820 2776 22876
rect 2776 22820 2832 22876
rect 2832 22820 2836 22876
rect 2772 22816 2836 22820
rect 2852 22876 2916 22880
rect 2852 22820 2856 22876
rect 2856 22820 2912 22876
rect 2912 22820 2916 22876
rect 2852 22816 2916 22820
rect 7612 22876 7676 22880
rect 7612 22820 7616 22876
rect 7616 22820 7672 22876
rect 7672 22820 7676 22876
rect 7612 22816 7676 22820
rect 7692 22876 7756 22880
rect 7692 22820 7696 22876
rect 7696 22820 7752 22876
rect 7752 22820 7756 22876
rect 7692 22816 7756 22820
rect 7772 22876 7836 22880
rect 7772 22820 7776 22876
rect 7776 22820 7832 22876
rect 7832 22820 7836 22876
rect 7772 22816 7836 22820
rect 7852 22876 7916 22880
rect 7852 22820 7856 22876
rect 7856 22820 7912 22876
rect 7912 22820 7916 22876
rect 7852 22816 7916 22820
rect 12612 22876 12676 22880
rect 12612 22820 12616 22876
rect 12616 22820 12672 22876
rect 12672 22820 12676 22876
rect 12612 22816 12676 22820
rect 12692 22876 12756 22880
rect 12692 22820 12696 22876
rect 12696 22820 12752 22876
rect 12752 22820 12756 22876
rect 12692 22816 12756 22820
rect 12772 22876 12836 22880
rect 12772 22820 12776 22876
rect 12776 22820 12832 22876
rect 12832 22820 12836 22876
rect 12772 22816 12836 22820
rect 12852 22876 12916 22880
rect 12852 22820 12856 22876
rect 12856 22820 12912 22876
rect 12912 22820 12916 22876
rect 12852 22816 12916 22820
rect 17612 22876 17676 22880
rect 17612 22820 17616 22876
rect 17616 22820 17672 22876
rect 17672 22820 17676 22876
rect 17612 22816 17676 22820
rect 17692 22876 17756 22880
rect 17692 22820 17696 22876
rect 17696 22820 17752 22876
rect 17752 22820 17756 22876
rect 17692 22816 17756 22820
rect 17772 22876 17836 22880
rect 17772 22820 17776 22876
rect 17776 22820 17832 22876
rect 17832 22820 17836 22876
rect 17772 22816 17836 22820
rect 17852 22876 17916 22880
rect 17852 22820 17856 22876
rect 17856 22820 17912 22876
rect 17912 22820 17916 22876
rect 17852 22816 17916 22820
rect 22612 22876 22676 22880
rect 22612 22820 22616 22876
rect 22616 22820 22672 22876
rect 22672 22820 22676 22876
rect 22612 22816 22676 22820
rect 22692 22876 22756 22880
rect 22692 22820 22696 22876
rect 22696 22820 22752 22876
rect 22752 22820 22756 22876
rect 22692 22816 22756 22820
rect 22772 22876 22836 22880
rect 22772 22820 22776 22876
rect 22776 22820 22832 22876
rect 22832 22820 22836 22876
rect 22772 22816 22836 22820
rect 22852 22876 22916 22880
rect 22852 22820 22856 22876
rect 22856 22820 22912 22876
rect 22912 22820 22916 22876
rect 22852 22816 22916 22820
rect 27612 22876 27676 22880
rect 27612 22820 27616 22876
rect 27616 22820 27672 22876
rect 27672 22820 27676 22876
rect 27612 22816 27676 22820
rect 27692 22876 27756 22880
rect 27692 22820 27696 22876
rect 27696 22820 27752 22876
rect 27752 22820 27756 22876
rect 27692 22816 27756 22820
rect 27772 22876 27836 22880
rect 27772 22820 27776 22876
rect 27776 22820 27832 22876
rect 27832 22820 27836 22876
rect 27772 22816 27836 22820
rect 27852 22876 27916 22880
rect 27852 22820 27856 22876
rect 27856 22820 27912 22876
rect 27912 22820 27916 22876
rect 27852 22816 27916 22820
rect 32612 22876 32676 22880
rect 32612 22820 32616 22876
rect 32616 22820 32672 22876
rect 32672 22820 32676 22876
rect 32612 22816 32676 22820
rect 32692 22876 32756 22880
rect 32692 22820 32696 22876
rect 32696 22820 32752 22876
rect 32752 22820 32756 22876
rect 32692 22816 32756 22820
rect 32772 22876 32836 22880
rect 32772 22820 32776 22876
rect 32776 22820 32832 22876
rect 32832 22820 32836 22876
rect 32772 22816 32836 22820
rect 32852 22876 32916 22880
rect 32852 22820 32856 22876
rect 32856 22820 32912 22876
rect 32912 22820 32916 22876
rect 32852 22816 32916 22820
rect 37612 22876 37676 22880
rect 37612 22820 37616 22876
rect 37616 22820 37672 22876
rect 37672 22820 37676 22876
rect 37612 22816 37676 22820
rect 37692 22876 37756 22880
rect 37692 22820 37696 22876
rect 37696 22820 37752 22876
rect 37752 22820 37756 22876
rect 37692 22816 37756 22820
rect 37772 22876 37836 22880
rect 37772 22820 37776 22876
rect 37776 22820 37832 22876
rect 37832 22820 37836 22876
rect 37772 22816 37836 22820
rect 37852 22876 37916 22880
rect 37852 22820 37856 22876
rect 37856 22820 37912 22876
rect 37912 22820 37916 22876
rect 37852 22816 37916 22820
rect 14964 22808 15028 22812
rect 14964 22752 14978 22808
rect 14978 22752 15028 22808
rect 14964 22748 15028 22752
rect 1952 22332 2016 22336
rect 1952 22276 1956 22332
rect 1956 22276 2012 22332
rect 2012 22276 2016 22332
rect 1952 22272 2016 22276
rect 2032 22332 2096 22336
rect 2032 22276 2036 22332
rect 2036 22276 2092 22332
rect 2092 22276 2096 22332
rect 2032 22272 2096 22276
rect 2112 22332 2176 22336
rect 2112 22276 2116 22332
rect 2116 22276 2172 22332
rect 2172 22276 2176 22332
rect 2112 22272 2176 22276
rect 2192 22332 2256 22336
rect 2192 22276 2196 22332
rect 2196 22276 2252 22332
rect 2252 22276 2256 22332
rect 2192 22272 2256 22276
rect 6952 22332 7016 22336
rect 6952 22276 6956 22332
rect 6956 22276 7012 22332
rect 7012 22276 7016 22332
rect 6952 22272 7016 22276
rect 7032 22332 7096 22336
rect 7032 22276 7036 22332
rect 7036 22276 7092 22332
rect 7092 22276 7096 22332
rect 7032 22272 7096 22276
rect 7112 22332 7176 22336
rect 7112 22276 7116 22332
rect 7116 22276 7172 22332
rect 7172 22276 7176 22332
rect 7112 22272 7176 22276
rect 7192 22332 7256 22336
rect 7192 22276 7196 22332
rect 7196 22276 7252 22332
rect 7252 22276 7256 22332
rect 7192 22272 7256 22276
rect 11952 22332 12016 22336
rect 11952 22276 11956 22332
rect 11956 22276 12012 22332
rect 12012 22276 12016 22332
rect 11952 22272 12016 22276
rect 12032 22332 12096 22336
rect 12032 22276 12036 22332
rect 12036 22276 12092 22332
rect 12092 22276 12096 22332
rect 12032 22272 12096 22276
rect 12112 22332 12176 22336
rect 12112 22276 12116 22332
rect 12116 22276 12172 22332
rect 12172 22276 12176 22332
rect 12112 22272 12176 22276
rect 12192 22332 12256 22336
rect 12192 22276 12196 22332
rect 12196 22276 12252 22332
rect 12252 22276 12256 22332
rect 12192 22272 12256 22276
rect 16952 22332 17016 22336
rect 16952 22276 16956 22332
rect 16956 22276 17012 22332
rect 17012 22276 17016 22332
rect 16952 22272 17016 22276
rect 17032 22332 17096 22336
rect 17032 22276 17036 22332
rect 17036 22276 17092 22332
rect 17092 22276 17096 22332
rect 17032 22272 17096 22276
rect 17112 22332 17176 22336
rect 17112 22276 17116 22332
rect 17116 22276 17172 22332
rect 17172 22276 17176 22332
rect 17112 22272 17176 22276
rect 17192 22332 17256 22336
rect 17192 22276 17196 22332
rect 17196 22276 17252 22332
rect 17252 22276 17256 22332
rect 17192 22272 17256 22276
rect 21952 22332 22016 22336
rect 21952 22276 21956 22332
rect 21956 22276 22012 22332
rect 22012 22276 22016 22332
rect 21952 22272 22016 22276
rect 22032 22332 22096 22336
rect 22032 22276 22036 22332
rect 22036 22276 22092 22332
rect 22092 22276 22096 22332
rect 22032 22272 22096 22276
rect 22112 22332 22176 22336
rect 22112 22276 22116 22332
rect 22116 22276 22172 22332
rect 22172 22276 22176 22332
rect 22112 22272 22176 22276
rect 22192 22332 22256 22336
rect 22192 22276 22196 22332
rect 22196 22276 22252 22332
rect 22252 22276 22256 22332
rect 22192 22272 22256 22276
rect 26952 22332 27016 22336
rect 26952 22276 26956 22332
rect 26956 22276 27012 22332
rect 27012 22276 27016 22332
rect 26952 22272 27016 22276
rect 27032 22332 27096 22336
rect 27032 22276 27036 22332
rect 27036 22276 27092 22332
rect 27092 22276 27096 22332
rect 27032 22272 27096 22276
rect 27112 22332 27176 22336
rect 27112 22276 27116 22332
rect 27116 22276 27172 22332
rect 27172 22276 27176 22332
rect 27112 22272 27176 22276
rect 27192 22332 27256 22336
rect 27192 22276 27196 22332
rect 27196 22276 27252 22332
rect 27252 22276 27256 22332
rect 27192 22272 27256 22276
rect 31952 22332 32016 22336
rect 31952 22276 31956 22332
rect 31956 22276 32012 22332
rect 32012 22276 32016 22332
rect 31952 22272 32016 22276
rect 32032 22332 32096 22336
rect 32032 22276 32036 22332
rect 32036 22276 32092 22332
rect 32092 22276 32096 22332
rect 32032 22272 32096 22276
rect 32112 22332 32176 22336
rect 32112 22276 32116 22332
rect 32116 22276 32172 22332
rect 32172 22276 32176 22332
rect 32112 22272 32176 22276
rect 32192 22332 32256 22336
rect 32192 22276 32196 22332
rect 32196 22276 32252 22332
rect 32252 22276 32256 22332
rect 32192 22272 32256 22276
rect 36952 22332 37016 22336
rect 36952 22276 36956 22332
rect 36956 22276 37012 22332
rect 37012 22276 37016 22332
rect 36952 22272 37016 22276
rect 37032 22332 37096 22336
rect 37032 22276 37036 22332
rect 37036 22276 37092 22332
rect 37092 22276 37096 22332
rect 37032 22272 37096 22276
rect 37112 22332 37176 22336
rect 37112 22276 37116 22332
rect 37116 22276 37172 22332
rect 37172 22276 37176 22332
rect 37112 22272 37176 22276
rect 37192 22332 37256 22336
rect 37192 22276 37196 22332
rect 37196 22276 37252 22332
rect 37252 22276 37256 22332
rect 37192 22272 37256 22276
rect 2612 21788 2676 21792
rect 2612 21732 2616 21788
rect 2616 21732 2672 21788
rect 2672 21732 2676 21788
rect 2612 21728 2676 21732
rect 2692 21788 2756 21792
rect 2692 21732 2696 21788
rect 2696 21732 2752 21788
rect 2752 21732 2756 21788
rect 2692 21728 2756 21732
rect 2772 21788 2836 21792
rect 2772 21732 2776 21788
rect 2776 21732 2832 21788
rect 2832 21732 2836 21788
rect 2772 21728 2836 21732
rect 2852 21788 2916 21792
rect 2852 21732 2856 21788
rect 2856 21732 2912 21788
rect 2912 21732 2916 21788
rect 2852 21728 2916 21732
rect 7612 21788 7676 21792
rect 7612 21732 7616 21788
rect 7616 21732 7672 21788
rect 7672 21732 7676 21788
rect 7612 21728 7676 21732
rect 7692 21788 7756 21792
rect 7692 21732 7696 21788
rect 7696 21732 7752 21788
rect 7752 21732 7756 21788
rect 7692 21728 7756 21732
rect 7772 21788 7836 21792
rect 7772 21732 7776 21788
rect 7776 21732 7832 21788
rect 7832 21732 7836 21788
rect 7772 21728 7836 21732
rect 7852 21788 7916 21792
rect 7852 21732 7856 21788
rect 7856 21732 7912 21788
rect 7912 21732 7916 21788
rect 7852 21728 7916 21732
rect 12612 21788 12676 21792
rect 12612 21732 12616 21788
rect 12616 21732 12672 21788
rect 12672 21732 12676 21788
rect 12612 21728 12676 21732
rect 12692 21788 12756 21792
rect 12692 21732 12696 21788
rect 12696 21732 12752 21788
rect 12752 21732 12756 21788
rect 12692 21728 12756 21732
rect 12772 21788 12836 21792
rect 12772 21732 12776 21788
rect 12776 21732 12832 21788
rect 12832 21732 12836 21788
rect 12772 21728 12836 21732
rect 12852 21788 12916 21792
rect 12852 21732 12856 21788
rect 12856 21732 12912 21788
rect 12912 21732 12916 21788
rect 12852 21728 12916 21732
rect 17612 21788 17676 21792
rect 17612 21732 17616 21788
rect 17616 21732 17672 21788
rect 17672 21732 17676 21788
rect 17612 21728 17676 21732
rect 17692 21788 17756 21792
rect 17692 21732 17696 21788
rect 17696 21732 17752 21788
rect 17752 21732 17756 21788
rect 17692 21728 17756 21732
rect 17772 21788 17836 21792
rect 17772 21732 17776 21788
rect 17776 21732 17832 21788
rect 17832 21732 17836 21788
rect 17772 21728 17836 21732
rect 17852 21788 17916 21792
rect 17852 21732 17856 21788
rect 17856 21732 17912 21788
rect 17912 21732 17916 21788
rect 17852 21728 17916 21732
rect 22612 21788 22676 21792
rect 22612 21732 22616 21788
rect 22616 21732 22672 21788
rect 22672 21732 22676 21788
rect 22612 21728 22676 21732
rect 22692 21788 22756 21792
rect 22692 21732 22696 21788
rect 22696 21732 22752 21788
rect 22752 21732 22756 21788
rect 22692 21728 22756 21732
rect 22772 21788 22836 21792
rect 22772 21732 22776 21788
rect 22776 21732 22832 21788
rect 22832 21732 22836 21788
rect 22772 21728 22836 21732
rect 22852 21788 22916 21792
rect 22852 21732 22856 21788
rect 22856 21732 22912 21788
rect 22912 21732 22916 21788
rect 22852 21728 22916 21732
rect 27612 21788 27676 21792
rect 27612 21732 27616 21788
rect 27616 21732 27672 21788
rect 27672 21732 27676 21788
rect 27612 21728 27676 21732
rect 27692 21788 27756 21792
rect 27692 21732 27696 21788
rect 27696 21732 27752 21788
rect 27752 21732 27756 21788
rect 27692 21728 27756 21732
rect 27772 21788 27836 21792
rect 27772 21732 27776 21788
rect 27776 21732 27832 21788
rect 27832 21732 27836 21788
rect 27772 21728 27836 21732
rect 27852 21788 27916 21792
rect 27852 21732 27856 21788
rect 27856 21732 27912 21788
rect 27912 21732 27916 21788
rect 27852 21728 27916 21732
rect 32612 21788 32676 21792
rect 32612 21732 32616 21788
rect 32616 21732 32672 21788
rect 32672 21732 32676 21788
rect 32612 21728 32676 21732
rect 32692 21788 32756 21792
rect 32692 21732 32696 21788
rect 32696 21732 32752 21788
rect 32752 21732 32756 21788
rect 32692 21728 32756 21732
rect 32772 21788 32836 21792
rect 32772 21732 32776 21788
rect 32776 21732 32832 21788
rect 32832 21732 32836 21788
rect 32772 21728 32836 21732
rect 32852 21788 32916 21792
rect 32852 21732 32856 21788
rect 32856 21732 32912 21788
rect 32912 21732 32916 21788
rect 32852 21728 32916 21732
rect 37612 21788 37676 21792
rect 37612 21732 37616 21788
rect 37616 21732 37672 21788
rect 37672 21732 37676 21788
rect 37612 21728 37676 21732
rect 37692 21788 37756 21792
rect 37692 21732 37696 21788
rect 37696 21732 37752 21788
rect 37752 21732 37756 21788
rect 37692 21728 37756 21732
rect 37772 21788 37836 21792
rect 37772 21732 37776 21788
rect 37776 21732 37832 21788
rect 37832 21732 37836 21788
rect 37772 21728 37836 21732
rect 37852 21788 37916 21792
rect 37852 21732 37856 21788
rect 37856 21732 37912 21788
rect 37912 21732 37916 21788
rect 37852 21728 37916 21732
rect 1952 21244 2016 21248
rect 1952 21188 1956 21244
rect 1956 21188 2012 21244
rect 2012 21188 2016 21244
rect 1952 21184 2016 21188
rect 2032 21244 2096 21248
rect 2032 21188 2036 21244
rect 2036 21188 2092 21244
rect 2092 21188 2096 21244
rect 2032 21184 2096 21188
rect 2112 21244 2176 21248
rect 2112 21188 2116 21244
rect 2116 21188 2172 21244
rect 2172 21188 2176 21244
rect 2112 21184 2176 21188
rect 2192 21244 2256 21248
rect 2192 21188 2196 21244
rect 2196 21188 2252 21244
rect 2252 21188 2256 21244
rect 2192 21184 2256 21188
rect 6952 21244 7016 21248
rect 6952 21188 6956 21244
rect 6956 21188 7012 21244
rect 7012 21188 7016 21244
rect 6952 21184 7016 21188
rect 7032 21244 7096 21248
rect 7032 21188 7036 21244
rect 7036 21188 7092 21244
rect 7092 21188 7096 21244
rect 7032 21184 7096 21188
rect 7112 21244 7176 21248
rect 7112 21188 7116 21244
rect 7116 21188 7172 21244
rect 7172 21188 7176 21244
rect 7112 21184 7176 21188
rect 7192 21244 7256 21248
rect 7192 21188 7196 21244
rect 7196 21188 7252 21244
rect 7252 21188 7256 21244
rect 7192 21184 7256 21188
rect 11952 21244 12016 21248
rect 11952 21188 11956 21244
rect 11956 21188 12012 21244
rect 12012 21188 12016 21244
rect 11952 21184 12016 21188
rect 12032 21244 12096 21248
rect 12032 21188 12036 21244
rect 12036 21188 12092 21244
rect 12092 21188 12096 21244
rect 12032 21184 12096 21188
rect 12112 21244 12176 21248
rect 12112 21188 12116 21244
rect 12116 21188 12172 21244
rect 12172 21188 12176 21244
rect 12112 21184 12176 21188
rect 12192 21244 12256 21248
rect 12192 21188 12196 21244
rect 12196 21188 12252 21244
rect 12252 21188 12256 21244
rect 12192 21184 12256 21188
rect 16952 21244 17016 21248
rect 16952 21188 16956 21244
rect 16956 21188 17012 21244
rect 17012 21188 17016 21244
rect 16952 21184 17016 21188
rect 17032 21244 17096 21248
rect 17032 21188 17036 21244
rect 17036 21188 17092 21244
rect 17092 21188 17096 21244
rect 17032 21184 17096 21188
rect 17112 21244 17176 21248
rect 17112 21188 17116 21244
rect 17116 21188 17172 21244
rect 17172 21188 17176 21244
rect 17112 21184 17176 21188
rect 17192 21244 17256 21248
rect 17192 21188 17196 21244
rect 17196 21188 17252 21244
rect 17252 21188 17256 21244
rect 17192 21184 17256 21188
rect 21952 21244 22016 21248
rect 21952 21188 21956 21244
rect 21956 21188 22012 21244
rect 22012 21188 22016 21244
rect 21952 21184 22016 21188
rect 22032 21244 22096 21248
rect 22032 21188 22036 21244
rect 22036 21188 22092 21244
rect 22092 21188 22096 21244
rect 22032 21184 22096 21188
rect 22112 21244 22176 21248
rect 22112 21188 22116 21244
rect 22116 21188 22172 21244
rect 22172 21188 22176 21244
rect 22112 21184 22176 21188
rect 22192 21244 22256 21248
rect 22192 21188 22196 21244
rect 22196 21188 22252 21244
rect 22252 21188 22256 21244
rect 22192 21184 22256 21188
rect 26952 21244 27016 21248
rect 26952 21188 26956 21244
rect 26956 21188 27012 21244
rect 27012 21188 27016 21244
rect 26952 21184 27016 21188
rect 27032 21244 27096 21248
rect 27032 21188 27036 21244
rect 27036 21188 27092 21244
rect 27092 21188 27096 21244
rect 27032 21184 27096 21188
rect 27112 21244 27176 21248
rect 27112 21188 27116 21244
rect 27116 21188 27172 21244
rect 27172 21188 27176 21244
rect 27112 21184 27176 21188
rect 27192 21244 27256 21248
rect 27192 21188 27196 21244
rect 27196 21188 27252 21244
rect 27252 21188 27256 21244
rect 27192 21184 27256 21188
rect 31952 21244 32016 21248
rect 31952 21188 31956 21244
rect 31956 21188 32012 21244
rect 32012 21188 32016 21244
rect 31952 21184 32016 21188
rect 32032 21244 32096 21248
rect 32032 21188 32036 21244
rect 32036 21188 32092 21244
rect 32092 21188 32096 21244
rect 32032 21184 32096 21188
rect 32112 21244 32176 21248
rect 32112 21188 32116 21244
rect 32116 21188 32172 21244
rect 32172 21188 32176 21244
rect 32112 21184 32176 21188
rect 32192 21244 32256 21248
rect 32192 21188 32196 21244
rect 32196 21188 32252 21244
rect 32252 21188 32256 21244
rect 32192 21184 32256 21188
rect 36952 21244 37016 21248
rect 36952 21188 36956 21244
rect 36956 21188 37012 21244
rect 37012 21188 37016 21244
rect 36952 21184 37016 21188
rect 37032 21244 37096 21248
rect 37032 21188 37036 21244
rect 37036 21188 37092 21244
rect 37092 21188 37096 21244
rect 37032 21184 37096 21188
rect 37112 21244 37176 21248
rect 37112 21188 37116 21244
rect 37116 21188 37172 21244
rect 37172 21188 37176 21244
rect 37112 21184 37176 21188
rect 37192 21244 37256 21248
rect 37192 21188 37196 21244
rect 37196 21188 37252 21244
rect 37252 21188 37256 21244
rect 37192 21184 37256 21188
rect 2612 20700 2676 20704
rect 2612 20644 2616 20700
rect 2616 20644 2672 20700
rect 2672 20644 2676 20700
rect 2612 20640 2676 20644
rect 2692 20700 2756 20704
rect 2692 20644 2696 20700
rect 2696 20644 2752 20700
rect 2752 20644 2756 20700
rect 2692 20640 2756 20644
rect 2772 20700 2836 20704
rect 2772 20644 2776 20700
rect 2776 20644 2832 20700
rect 2832 20644 2836 20700
rect 2772 20640 2836 20644
rect 2852 20700 2916 20704
rect 2852 20644 2856 20700
rect 2856 20644 2912 20700
rect 2912 20644 2916 20700
rect 2852 20640 2916 20644
rect 7612 20700 7676 20704
rect 7612 20644 7616 20700
rect 7616 20644 7672 20700
rect 7672 20644 7676 20700
rect 7612 20640 7676 20644
rect 7692 20700 7756 20704
rect 7692 20644 7696 20700
rect 7696 20644 7752 20700
rect 7752 20644 7756 20700
rect 7692 20640 7756 20644
rect 7772 20700 7836 20704
rect 7772 20644 7776 20700
rect 7776 20644 7832 20700
rect 7832 20644 7836 20700
rect 7772 20640 7836 20644
rect 7852 20700 7916 20704
rect 7852 20644 7856 20700
rect 7856 20644 7912 20700
rect 7912 20644 7916 20700
rect 7852 20640 7916 20644
rect 12612 20700 12676 20704
rect 12612 20644 12616 20700
rect 12616 20644 12672 20700
rect 12672 20644 12676 20700
rect 12612 20640 12676 20644
rect 12692 20700 12756 20704
rect 12692 20644 12696 20700
rect 12696 20644 12752 20700
rect 12752 20644 12756 20700
rect 12692 20640 12756 20644
rect 12772 20700 12836 20704
rect 12772 20644 12776 20700
rect 12776 20644 12832 20700
rect 12832 20644 12836 20700
rect 12772 20640 12836 20644
rect 12852 20700 12916 20704
rect 12852 20644 12856 20700
rect 12856 20644 12912 20700
rect 12912 20644 12916 20700
rect 12852 20640 12916 20644
rect 17612 20700 17676 20704
rect 17612 20644 17616 20700
rect 17616 20644 17672 20700
rect 17672 20644 17676 20700
rect 17612 20640 17676 20644
rect 17692 20700 17756 20704
rect 17692 20644 17696 20700
rect 17696 20644 17752 20700
rect 17752 20644 17756 20700
rect 17692 20640 17756 20644
rect 17772 20700 17836 20704
rect 17772 20644 17776 20700
rect 17776 20644 17832 20700
rect 17832 20644 17836 20700
rect 17772 20640 17836 20644
rect 17852 20700 17916 20704
rect 17852 20644 17856 20700
rect 17856 20644 17912 20700
rect 17912 20644 17916 20700
rect 17852 20640 17916 20644
rect 22612 20700 22676 20704
rect 22612 20644 22616 20700
rect 22616 20644 22672 20700
rect 22672 20644 22676 20700
rect 22612 20640 22676 20644
rect 22692 20700 22756 20704
rect 22692 20644 22696 20700
rect 22696 20644 22752 20700
rect 22752 20644 22756 20700
rect 22692 20640 22756 20644
rect 22772 20700 22836 20704
rect 22772 20644 22776 20700
rect 22776 20644 22832 20700
rect 22832 20644 22836 20700
rect 22772 20640 22836 20644
rect 22852 20700 22916 20704
rect 22852 20644 22856 20700
rect 22856 20644 22912 20700
rect 22912 20644 22916 20700
rect 22852 20640 22916 20644
rect 27612 20700 27676 20704
rect 27612 20644 27616 20700
rect 27616 20644 27672 20700
rect 27672 20644 27676 20700
rect 27612 20640 27676 20644
rect 27692 20700 27756 20704
rect 27692 20644 27696 20700
rect 27696 20644 27752 20700
rect 27752 20644 27756 20700
rect 27692 20640 27756 20644
rect 27772 20700 27836 20704
rect 27772 20644 27776 20700
rect 27776 20644 27832 20700
rect 27832 20644 27836 20700
rect 27772 20640 27836 20644
rect 27852 20700 27916 20704
rect 27852 20644 27856 20700
rect 27856 20644 27912 20700
rect 27912 20644 27916 20700
rect 27852 20640 27916 20644
rect 32612 20700 32676 20704
rect 32612 20644 32616 20700
rect 32616 20644 32672 20700
rect 32672 20644 32676 20700
rect 32612 20640 32676 20644
rect 32692 20700 32756 20704
rect 32692 20644 32696 20700
rect 32696 20644 32752 20700
rect 32752 20644 32756 20700
rect 32692 20640 32756 20644
rect 32772 20700 32836 20704
rect 32772 20644 32776 20700
rect 32776 20644 32832 20700
rect 32832 20644 32836 20700
rect 32772 20640 32836 20644
rect 32852 20700 32916 20704
rect 32852 20644 32856 20700
rect 32856 20644 32912 20700
rect 32912 20644 32916 20700
rect 32852 20640 32916 20644
rect 37612 20700 37676 20704
rect 37612 20644 37616 20700
rect 37616 20644 37672 20700
rect 37672 20644 37676 20700
rect 37612 20640 37676 20644
rect 37692 20700 37756 20704
rect 37692 20644 37696 20700
rect 37696 20644 37752 20700
rect 37752 20644 37756 20700
rect 37692 20640 37756 20644
rect 37772 20700 37836 20704
rect 37772 20644 37776 20700
rect 37776 20644 37832 20700
rect 37832 20644 37836 20700
rect 37772 20640 37836 20644
rect 37852 20700 37916 20704
rect 37852 20644 37856 20700
rect 37856 20644 37912 20700
rect 37912 20644 37916 20700
rect 37852 20640 37916 20644
rect 1952 20156 2016 20160
rect 1952 20100 1956 20156
rect 1956 20100 2012 20156
rect 2012 20100 2016 20156
rect 1952 20096 2016 20100
rect 2032 20156 2096 20160
rect 2032 20100 2036 20156
rect 2036 20100 2092 20156
rect 2092 20100 2096 20156
rect 2032 20096 2096 20100
rect 2112 20156 2176 20160
rect 2112 20100 2116 20156
rect 2116 20100 2172 20156
rect 2172 20100 2176 20156
rect 2112 20096 2176 20100
rect 2192 20156 2256 20160
rect 2192 20100 2196 20156
rect 2196 20100 2252 20156
rect 2252 20100 2256 20156
rect 2192 20096 2256 20100
rect 6952 20156 7016 20160
rect 6952 20100 6956 20156
rect 6956 20100 7012 20156
rect 7012 20100 7016 20156
rect 6952 20096 7016 20100
rect 7032 20156 7096 20160
rect 7032 20100 7036 20156
rect 7036 20100 7092 20156
rect 7092 20100 7096 20156
rect 7032 20096 7096 20100
rect 7112 20156 7176 20160
rect 7112 20100 7116 20156
rect 7116 20100 7172 20156
rect 7172 20100 7176 20156
rect 7112 20096 7176 20100
rect 7192 20156 7256 20160
rect 7192 20100 7196 20156
rect 7196 20100 7252 20156
rect 7252 20100 7256 20156
rect 7192 20096 7256 20100
rect 11952 20156 12016 20160
rect 11952 20100 11956 20156
rect 11956 20100 12012 20156
rect 12012 20100 12016 20156
rect 11952 20096 12016 20100
rect 12032 20156 12096 20160
rect 12032 20100 12036 20156
rect 12036 20100 12092 20156
rect 12092 20100 12096 20156
rect 12032 20096 12096 20100
rect 12112 20156 12176 20160
rect 12112 20100 12116 20156
rect 12116 20100 12172 20156
rect 12172 20100 12176 20156
rect 12112 20096 12176 20100
rect 12192 20156 12256 20160
rect 12192 20100 12196 20156
rect 12196 20100 12252 20156
rect 12252 20100 12256 20156
rect 12192 20096 12256 20100
rect 16952 20156 17016 20160
rect 16952 20100 16956 20156
rect 16956 20100 17012 20156
rect 17012 20100 17016 20156
rect 16952 20096 17016 20100
rect 17032 20156 17096 20160
rect 17032 20100 17036 20156
rect 17036 20100 17092 20156
rect 17092 20100 17096 20156
rect 17032 20096 17096 20100
rect 17112 20156 17176 20160
rect 17112 20100 17116 20156
rect 17116 20100 17172 20156
rect 17172 20100 17176 20156
rect 17112 20096 17176 20100
rect 17192 20156 17256 20160
rect 17192 20100 17196 20156
rect 17196 20100 17252 20156
rect 17252 20100 17256 20156
rect 17192 20096 17256 20100
rect 21952 20156 22016 20160
rect 21952 20100 21956 20156
rect 21956 20100 22012 20156
rect 22012 20100 22016 20156
rect 21952 20096 22016 20100
rect 22032 20156 22096 20160
rect 22032 20100 22036 20156
rect 22036 20100 22092 20156
rect 22092 20100 22096 20156
rect 22032 20096 22096 20100
rect 22112 20156 22176 20160
rect 22112 20100 22116 20156
rect 22116 20100 22172 20156
rect 22172 20100 22176 20156
rect 22112 20096 22176 20100
rect 22192 20156 22256 20160
rect 22192 20100 22196 20156
rect 22196 20100 22252 20156
rect 22252 20100 22256 20156
rect 22192 20096 22256 20100
rect 26952 20156 27016 20160
rect 26952 20100 26956 20156
rect 26956 20100 27012 20156
rect 27012 20100 27016 20156
rect 26952 20096 27016 20100
rect 27032 20156 27096 20160
rect 27032 20100 27036 20156
rect 27036 20100 27092 20156
rect 27092 20100 27096 20156
rect 27032 20096 27096 20100
rect 27112 20156 27176 20160
rect 27112 20100 27116 20156
rect 27116 20100 27172 20156
rect 27172 20100 27176 20156
rect 27112 20096 27176 20100
rect 27192 20156 27256 20160
rect 27192 20100 27196 20156
rect 27196 20100 27252 20156
rect 27252 20100 27256 20156
rect 27192 20096 27256 20100
rect 31952 20156 32016 20160
rect 31952 20100 31956 20156
rect 31956 20100 32012 20156
rect 32012 20100 32016 20156
rect 31952 20096 32016 20100
rect 32032 20156 32096 20160
rect 32032 20100 32036 20156
rect 32036 20100 32092 20156
rect 32092 20100 32096 20156
rect 32032 20096 32096 20100
rect 32112 20156 32176 20160
rect 32112 20100 32116 20156
rect 32116 20100 32172 20156
rect 32172 20100 32176 20156
rect 32112 20096 32176 20100
rect 32192 20156 32256 20160
rect 32192 20100 32196 20156
rect 32196 20100 32252 20156
rect 32252 20100 32256 20156
rect 32192 20096 32256 20100
rect 36952 20156 37016 20160
rect 36952 20100 36956 20156
rect 36956 20100 37012 20156
rect 37012 20100 37016 20156
rect 36952 20096 37016 20100
rect 37032 20156 37096 20160
rect 37032 20100 37036 20156
rect 37036 20100 37092 20156
rect 37092 20100 37096 20156
rect 37032 20096 37096 20100
rect 37112 20156 37176 20160
rect 37112 20100 37116 20156
rect 37116 20100 37172 20156
rect 37172 20100 37176 20156
rect 37112 20096 37176 20100
rect 37192 20156 37256 20160
rect 37192 20100 37196 20156
rect 37196 20100 37252 20156
rect 37252 20100 37256 20156
rect 37192 20096 37256 20100
rect 2612 19612 2676 19616
rect 2612 19556 2616 19612
rect 2616 19556 2672 19612
rect 2672 19556 2676 19612
rect 2612 19552 2676 19556
rect 2692 19612 2756 19616
rect 2692 19556 2696 19612
rect 2696 19556 2752 19612
rect 2752 19556 2756 19612
rect 2692 19552 2756 19556
rect 2772 19612 2836 19616
rect 2772 19556 2776 19612
rect 2776 19556 2832 19612
rect 2832 19556 2836 19612
rect 2772 19552 2836 19556
rect 2852 19612 2916 19616
rect 2852 19556 2856 19612
rect 2856 19556 2912 19612
rect 2912 19556 2916 19612
rect 2852 19552 2916 19556
rect 7612 19612 7676 19616
rect 7612 19556 7616 19612
rect 7616 19556 7672 19612
rect 7672 19556 7676 19612
rect 7612 19552 7676 19556
rect 7692 19612 7756 19616
rect 7692 19556 7696 19612
rect 7696 19556 7752 19612
rect 7752 19556 7756 19612
rect 7692 19552 7756 19556
rect 7772 19612 7836 19616
rect 7772 19556 7776 19612
rect 7776 19556 7832 19612
rect 7832 19556 7836 19612
rect 7772 19552 7836 19556
rect 7852 19612 7916 19616
rect 7852 19556 7856 19612
rect 7856 19556 7912 19612
rect 7912 19556 7916 19612
rect 7852 19552 7916 19556
rect 12612 19612 12676 19616
rect 12612 19556 12616 19612
rect 12616 19556 12672 19612
rect 12672 19556 12676 19612
rect 12612 19552 12676 19556
rect 12692 19612 12756 19616
rect 12692 19556 12696 19612
rect 12696 19556 12752 19612
rect 12752 19556 12756 19612
rect 12692 19552 12756 19556
rect 12772 19612 12836 19616
rect 12772 19556 12776 19612
rect 12776 19556 12832 19612
rect 12832 19556 12836 19612
rect 12772 19552 12836 19556
rect 12852 19612 12916 19616
rect 12852 19556 12856 19612
rect 12856 19556 12912 19612
rect 12912 19556 12916 19612
rect 12852 19552 12916 19556
rect 17612 19612 17676 19616
rect 17612 19556 17616 19612
rect 17616 19556 17672 19612
rect 17672 19556 17676 19612
rect 17612 19552 17676 19556
rect 17692 19612 17756 19616
rect 17692 19556 17696 19612
rect 17696 19556 17752 19612
rect 17752 19556 17756 19612
rect 17692 19552 17756 19556
rect 17772 19612 17836 19616
rect 17772 19556 17776 19612
rect 17776 19556 17832 19612
rect 17832 19556 17836 19612
rect 17772 19552 17836 19556
rect 17852 19612 17916 19616
rect 17852 19556 17856 19612
rect 17856 19556 17912 19612
rect 17912 19556 17916 19612
rect 17852 19552 17916 19556
rect 22612 19612 22676 19616
rect 22612 19556 22616 19612
rect 22616 19556 22672 19612
rect 22672 19556 22676 19612
rect 22612 19552 22676 19556
rect 22692 19612 22756 19616
rect 22692 19556 22696 19612
rect 22696 19556 22752 19612
rect 22752 19556 22756 19612
rect 22692 19552 22756 19556
rect 22772 19612 22836 19616
rect 22772 19556 22776 19612
rect 22776 19556 22832 19612
rect 22832 19556 22836 19612
rect 22772 19552 22836 19556
rect 22852 19612 22916 19616
rect 22852 19556 22856 19612
rect 22856 19556 22912 19612
rect 22912 19556 22916 19612
rect 22852 19552 22916 19556
rect 27612 19612 27676 19616
rect 27612 19556 27616 19612
rect 27616 19556 27672 19612
rect 27672 19556 27676 19612
rect 27612 19552 27676 19556
rect 27692 19612 27756 19616
rect 27692 19556 27696 19612
rect 27696 19556 27752 19612
rect 27752 19556 27756 19612
rect 27692 19552 27756 19556
rect 27772 19612 27836 19616
rect 27772 19556 27776 19612
rect 27776 19556 27832 19612
rect 27832 19556 27836 19612
rect 27772 19552 27836 19556
rect 27852 19612 27916 19616
rect 27852 19556 27856 19612
rect 27856 19556 27912 19612
rect 27912 19556 27916 19612
rect 27852 19552 27916 19556
rect 32612 19612 32676 19616
rect 32612 19556 32616 19612
rect 32616 19556 32672 19612
rect 32672 19556 32676 19612
rect 32612 19552 32676 19556
rect 32692 19612 32756 19616
rect 32692 19556 32696 19612
rect 32696 19556 32752 19612
rect 32752 19556 32756 19612
rect 32692 19552 32756 19556
rect 32772 19612 32836 19616
rect 32772 19556 32776 19612
rect 32776 19556 32832 19612
rect 32832 19556 32836 19612
rect 32772 19552 32836 19556
rect 32852 19612 32916 19616
rect 32852 19556 32856 19612
rect 32856 19556 32912 19612
rect 32912 19556 32916 19612
rect 32852 19552 32916 19556
rect 37612 19612 37676 19616
rect 37612 19556 37616 19612
rect 37616 19556 37672 19612
rect 37672 19556 37676 19612
rect 37612 19552 37676 19556
rect 37692 19612 37756 19616
rect 37692 19556 37696 19612
rect 37696 19556 37752 19612
rect 37752 19556 37756 19612
rect 37692 19552 37756 19556
rect 37772 19612 37836 19616
rect 37772 19556 37776 19612
rect 37776 19556 37832 19612
rect 37832 19556 37836 19612
rect 37772 19552 37836 19556
rect 37852 19612 37916 19616
rect 37852 19556 37856 19612
rect 37856 19556 37912 19612
rect 37912 19556 37916 19612
rect 37852 19552 37916 19556
rect 1952 19068 2016 19072
rect 1952 19012 1956 19068
rect 1956 19012 2012 19068
rect 2012 19012 2016 19068
rect 1952 19008 2016 19012
rect 2032 19068 2096 19072
rect 2032 19012 2036 19068
rect 2036 19012 2092 19068
rect 2092 19012 2096 19068
rect 2032 19008 2096 19012
rect 2112 19068 2176 19072
rect 2112 19012 2116 19068
rect 2116 19012 2172 19068
rect 2172 19012 2176 19068
rect 2112 19008 2176 19012
rect 2192 19068 2256 19072
rect 2192 19012 2196 19068
rect 2196 19012 2252 19068
rect 2252 19012 2256 19068
rect 2192 19008 2256 19012
rect 6952 19068 7016 19072
rect 6952 19012 6956 19068
rect 6956 19012 7012 19068
rect 7012 19012 7016 19068
rect 6952 19008 7016 19012
rect 7032 19068 7096 19072
rect 7032 19012 7036 19068
rect 7036 19012 7092 19068
rect 7092 19012 7096 19068
rect 7032 19008 7096 19012
rect 7112 19068 7176 19072
rect 7112 19012 7116 19068
rect 7116 19012 7172 19068
rect 7172 19012 7176 19068
rect 7112 19008 7176 19012
rect 7192 19068 7256 19072
rect 7192 19012 7196 19068
rect 7196 19012 7252 19068
rect 7252 19012 7256 19068
rect 7192 19008 7256 19012
rect 11952 19068 12016 19072
rect 11952 19012 11956 19068
rect 11956 19012 12012 19068
rect 12012 19012 12016 19068
rect 11952 19008 12016 19012
rect 12032 19068 12096 19072
rect 12032 19012 12036 19068
rect 12036 19012 12092 19068
rect 12092 19012 12096 19068
rect 12032 19008 12096 19012
rect 12112 19068 12176 19072
rect 12112 19012 12116 19068
rect 12116 19012 12172 19068
rect 12172 19012 12176 19068
rect 12112 19008 12176 19012
rect 12192 19068 12256 19072
rect 12192 19012 12196 19068
rect 12196 19012 12252 19068
rect 12252 19012 12256 19068
rect 12192 19008 12256 19012
rect 16952 19068 17016 19072
rect 16952 19012 16956 19068
rect 16956 19012 17012 19068
rect 17012 19012 17016 19068
rect 16952 19008 17016 19012
rect 17032 19068 17096 19072
rect 17032 19012 17036 19068
rect 17036 19012 17092 19068
rect 17092 19012 17096 19068
rect 17032 19008 17096 19012
rect 17112 19068 17176 19072
rect 17112 19012 17116 19068
rect 17116 19012 17172 19068
rect 17172 19012 17176 19068
rect 17112 19008 17176 19012
rect 17192 19068 17256 19072
rect 17192 19012 17196 19068
rect 17196 19012 17252 19068
rect 17252 19012 17256 19068
rect 17192 19008 17256 19012
rect 21952 19068 22016 19072
rect 21952 19012 21956 19068
rect 21956 19012 22012 19068
rect 22012 19012 22016 19068
rect 21952 19008 22016 19012
rect 22032 19068 22096 19072
rect 22032 19012 22036 19068
rect 22036 19012 22092 19068
rect 22092 19012 22096 19068
rect 22032 19008 22096 19012
rect 22112 19068 22176 19072
rect 22112 19012 22116 19068
rect 22116 19012 22172 19068
rect 22172 19012 22176 19068
rect 22112 19008 22176 19012
rect 22192 19068 22256 19072
rect 22192 19012 22196 19068
rect 22196 19012 22252 19068
rect 22252 19012 22256 19068
rect 22192 19008 22256 19012
rect 26952 19068 27016 19072
rect 26952 19012 26956 19068
rect 26956 19012 27012 19068
rect 27012 19012 27016 19068
rect 26952 19008 27016 19012
rect 27032 19068 27096 19072
rect 27032 19012 27036 19068
rect 27036 19012 27092 19068
rect 27092 19012 27096 19068
rect 27032 19008 27096 19012
rect 27112 19068 27176 19072
rect 27112 19012 27116 19068
rect 27116 19012 27172 19068
rect 27172 19012 27176 19068
rect 27112 19008 27176 19012
rect 27192 19068 27256 19072
rect 27192 19012 27196 19068
rect 27196 19012 27252 19068
rect 27252 19012 27256 19068
rect 27192 19008 27256 19012
rect 31952 19068 32016 19072
rect 31952 19012 31956 19068
rect 31956 19012 32012 19068
rect 32012 19012 32016 19068
rect 31952 19008 32016 19012
rect 32032 19068 32096 19072
rect 32032 19012 32036 19068
rect 32036 19012 32092 19068
rect 32092 19012 32096 19068
rect 32032 19008 32096 19012
rect 32112 19068 32176 19072
rect 32112 19012 32116 19068
rect 32116 19012 32172 19068
rect 32172 19012 32176 19068
rect 32112 19008 32176 19012
rect 32192 19068 32256 19072
rect 32192 19012 32196 19068
rect 32196 19012 32252 19068
rect 32252 19012 32256 19068
rect 32192 19008 32256 19012
rect 36952 19068 37016 19072
rect 36952 19012 36956 19068
rect 36956 19012 37012 19068
rect 37012 19012 37016 19068
rect 36952 19008 37016 19012
rect 37032 19068 37096 19072
rect 37032 19012 37036 19068
rect 37036 19012 37092 19068
rect 37092 19012 37096 19068
rect 37032 19008 37096 19012
rect 37112 19068 37176 19072
rect 37112 19012 37116 19068
rect 37116 19012 37172 19068
rect 37172 19012 37176 19068
rect 37112 19008 37176 19012
rect 37192 19068 37256 19072
rect 37192 19012 37196 19068
rect 37196 19012 37252 19068
rect 37252 19012 37256 19068
rect 37192 19008 37256 19012
rect 2612 18524 2676 18528
rect 2612 18468 2616 18524
rect 2616 18468 2672 18524
rect 2672 18468 2676 18524
rect 2612 18464 2676 18468
rect 2692 18524 2756 18528
rect 2692 18468 2696 18524
rect 2696 18468 2752 18524
rect 2752 18468 2756 18524
rect 2692 18464 2756 18468
rect 2772 18524 2836 18528
rect 2772 18468 2776 18524
rect 2776 18468 2832 18524
rect 2832 18468 2836 18524
rect 2772 18464 2836 18468
rect 2852 18524 2916 18528
rect 2852 18468 2856 18524
rect 2856 18468 2912 18524
rect 2912 18468 2916 18524
rect 2852 18464 2916 18468
rect 7612 18524 7676 18528
rect 7612 18468 7616 18524
rect 7616 18468 7672 18524
rect 7672 18468 7676 18524
rect 7612 18464 7676 18468
rect 7692 18524 7756 18528
rect 7692 18468 7696 18524
rect 7696 18468 7752 18524
rect 7752 18468 7756 18524
rect 7692 18464 7756 18468
rect 7772 18524 7836 18528
rect 7772 18468 7776 18524
rect 7776 18468 7832 18524
rect 7832 18468 7836 18524
rect 7772 18464 7836 18468
rect 7852 18524 7916 18528
rect 7852 18468 7856 18524
rect 7856 18468 7912 18524
rect 7912 18468 7916 18524
rect 7852 18464 7916 18468
rect 12612 18524 12676 18528
rect 12612 18468 12616 18524
rect 12616 18468 12672 18524
rect 12672 18468 12676 18524
rect 12612 18464 12676 18468
rect 12692 18524 12756 18528
rect 12692 18468 12696 18524
rect 12696 18468 12752 18524
rect 12752 18468 12756 18524
rect 12692 18464 12756 18468
rect 12772 18524 12836 18528
rect 12772 18468 12776 18524
rect 12776 18468 12832 18524
rect 12832 18468 12836 18524
rect 12772 18464 12836 18468
rect 12852 18524 12916 18528
rect 12852 18468 12856 18524
rect 12856 18468 12912 18524
rect 12912 18468 12916 18524
rect 12852 18464 12916 18468
rect 17612 18524 17676 18528
rect 17612 18468 17616 18524
rect 17616 18468 17672 18524
rect 17672 18468 17676 18524
rect 17612 18464 17676 18468
rect 17692 18524 17756 18528
rect 17692 18468 17696 18524
rect 17696 18468 17752 18524
rect 17752 18468 17756 18524
rect 17692 18464 17756 18468
rect 17772 18524 17836 18528
rect 17772 18468 17776 18524
rect 17776 18468 17832 18524
rect 17832 18468 17836 18524
rect 17772 18464 17836 18468
rect 17852 18524 17916 18528
rect 17852 18468 17856 18524
rect 17856 18468 17912 18524
rect 17912 18468 17916 18524
rect 17852 18464 17916 18468
rect 22612 18524 22676 18528
rect 22612 18468 22616 18524
rect 22616 18468 22672 18524
rect 22672 18468 22676 18524
rect 22612 18464 22676 18468
rect 22692 18524 22756 18528
rect 22692 18468 22696 18524
rect 22696 18468 22752 18524
rect 22752 18468 22756 18524
rect 22692 18464 22756 18468
rect 22772 18524 22836 18528
rect 22772 18468 22776 18524
rect 22776 18468 22832 18524
rect 22832 18468 22836 18524
rect 22772 18464 22836 18468
rect 22852 18524 22916 18528
rect 22852 18468 22856 18524
rect 22856 18468 22912 18524
rect 22912 18468 22916 18524
rect 22852 18464 22916 18468
rect 27612 18524 27676 18528
rect 27612 18468 27616 18524
rect 27616 18468 27672 18524
rect 27672 18468 27676 18524
rect 27612 18464 27676 18468
rect 27692 18524 27756 18528
rect 27692 18468 27696 18524
rect 27696 18468 27752 18524
rect 27752 18468 27756 18524
rect 27692 18464 27756 18468
rect 27772 18524 27836 18528
rect 27772 18468 27776 18524
rect 27776 18468 27832 18524
rect 27832 18468 27836 18524
rect 27772 18464 27836 18468
rect 27852 18524 27916 18528
rect 27852 18468 27856 18524
rect 27856 18468 27912 18524
rect 27912 18468 27916 18524
rect 27852 18464 27916 18468
rect 32612 18524 32676 18528
rect 32612 18468 32616 18524
rect 32616 18468 32672 18524
rect 32672 18468 32676 18524
rect 32612 18464 32676 18468
rect 32692 18524 32756 18528
rect 32692 18468 32696 18524
rect 32696 18468 32752 18524
rect 32752 18468 32756 18524
rect 32692 18464 32756 18468
rect 32772 18524 32836 18528
rect 32772 18468 32776 18524
rect 32776 18468 32832 18524
rect 32832 18468 32836 18524
rect 32772 18464 32836 18468
rect 32852 18524 32916 18528
rect 32852 18468 32856 18524
rect 32856 18468 32912 18524
rect 32912 18468 32916 18524
rect 32852 18464 32916 18468
rect 37612 18524 37676 18528
rect 37612 18468 37616 18524
rect 37616 18468 37672 18524
rect 37672 18468 37676 18524
rect 37612 18464 37676 18468
rect 37692 18524 37756 18528
rect 37692 18468 37696 18524
rect 37696 18468 37752 18524
rect 37752 18468 37756 18524
rect 37692 18464 37756 18468
rect 37772 18524 37836 18528
rect 37772 18468 37776 18524
rect 37776 18468 37832 18524
rect 37832 18468 37836 18524
rect 37772 18464 37836 18468
rect 37852 18524 37916 18528
rect 37852 18468 37856 18524
rect 37856 18468 37912 18524
rect 37912 18468 37916 18524
rect 37852 18464 37916 18468
rect 1952 17980 2016 17984
rect 1952 17924 1956 17980
rect 1956 17924 2012 17980
rect 2012 17924 2016 17980
rect 1952 17920 2016 17924
rect 2032 17980 2096 17984
rect 2032 17924 2036 17980
rect 2036 17924 2092 17980
rect 2092 17924 2096 17980
rect 2032 17920 2096 17924
rect 2112 17980 2176 17984
rect 2112 17924 2116 17980
rect 2116 17924 2172 17980
rect 2172 17924 2176 17980
rect 2112 17920 2176 17924
rect 2192 17980 2256 17984
rect 2192 17924 2196 17980
rect 2196 17924 2252 17980
rect 2252 17924 2256 17980
rect 2192 17920 2256 17924
rect 6952 17980 7016 17984
rect 6952 17924 6956 17980
rect 6956 17924 7012 17980
rect 7012 17924 7016 17980
rect 6952 17920 7016 17924
rect 7032 17980 7096 17984
rect 7032 17924 7036 17980
rect 7036 17924 7092 17980
rect 7092 17924 7096 17980
rect 7032 17920 7096 17924
rect 7112 17980 7176 17984
rect 7112 17924 7116 17980
rect 7116 17924 7172 17980
rect 7172 17924 7176 17980
rect 7112 17920 7176 17924
rect 7192 17980 7256 17984
rect 7192 17924 7196 17980
rect 7196 17924 7252 17980
rect 7252 17924 7256 17980
rect 7192 17920 7256 17924
rect 11952 17980 12016 17984
rect 11952 17924 11956 17980
rect 11956 17924 12012 17980
rect 12012 17924 12016 17980
rect 11952 17920 12016 17924
rect 12032 17980 12096 17984
rect 12032 17924 12036 17980
rect 12036 17924 12092 17980
rect 12092 17924 12096 17980
rect 12032 17920 12096 17924
rect 12112 17980 12176 17984
rect 12112 17924 12116 17980
rect 12116 17924 12172 17980
rect 12172 17924 12176 17980
rect 12112 17920 12176 17924
rect 12192 17980 12256 17984
rect 12192 17924 12196 17980
rect 12196 17924 12252 17980
rect 12252 17924 12256 17980
rect 12192 17920 12256 17924
rect 16952 17980 17016 17984
rect 16952 17924 16956 17980
rect 16956 17924 17012 17980
rect 17012 17924 17016 17980
rect 16952 17920 17016 17924
rect 17032 17980 17096 17984
rect 17032 17924 17036 17980
rect 17036 17924 17092 17980
rect 17092 17924 17096 17980
rect 17032 17920 17096 17924
rect 17112 17980 17176 17984
rect 17112 17924 17116 17980
rect 17116 17924 17172 17980
rect 17172 17924 17176 17980
rect 17112 17920 17176 17924
rect 17192 17980 17256 17984
rect 17192 17924 17196 17980
rect 17196 17924 17252 17980
rect 17252 17924 17256 17980
rect 17192 17920 17256 17924
rect 21952 17980 22016 17984
rect 21952 17924 21956 17980
rect 21956 17924 22012 17980
rect 22012 17924 22016 17980
rect 21952 17920 22016 17924
rect 22032 17980 22096 17984
rect 22032 17924 22036 17980
rect 22036 17924 22092 17980
rect 22092 17924 22096 17980
rect 22032 17920 22096 17924
rect 22112 17980 22176 17984
rect 22112 17924 22116 17980
rect 22116 17924 22172 17980
rect 22172 17924 22176 17980
rect 22112 17920 22176 17924
rect 22192 17980 22256 17984
rect 22192 17924 22196 17980
rect 22196 17924 22252 17980
rect 22252 17924 22256 17980
rect 22192 17920 22256 17924
rect 26952 17980 27016 17984
rect 26952 17924 26956 17980
rect 26956 17924 27012 17980
rect 27012 17924 27016 17980
rect 26952 17920 27016 17924
rect 27032 17980 27096 17984
rect 27032 17924 27036 17980
rect 27036 17924 27092 17980
rect 27092 17924 27096 17980
rect 27032 17920 27096 17924
rect 27112 17980 27176 17984
rect 27112 17924 27116 17980
rect 27116 17924 27172 17980
rect 27172 17924 27176 17980
rect 27112 17920 27176 17924
rect 27192 17980 27256 17984
rect 27192 17924 27196 17980
rect 27196 17924 27252 17980
rect 27252 17924 27256 17980
rect 27192 17920 27256 17924
rect 31952 17980 32016 17984
rect 31952 17924 31956 17980
rect 31956 17924 32012 17980
rect 32012 17924 32016 17980
rect 31952 17920 32016 17924
rect 32032 17980 32096 17984
rect 32032 17924 32036 17980
rect 32036 17924 32092 17980
rect 32092 17924 32096 17980
rect 32032 17920 32096 17924
rect 32112 17980 32176 17984
rect 32112 17924 32116 17980
rect 32116 17924 32172 17980
rect 32172 17924 32176 17980
rect 32112 17920 32176 17924
rect 32192 17980 32256 17984
rect 32192 17924 32196 17980
rect 32196 17924 32252 17980
rect 32252 17924 32256 17980
rect 32192 17920 32256 17924
rect 36952 17980 37016 17984
rect 36952 17924 36956 17980
rect 36956 17924 37012 17980
rect 37012 17924 37016 17980
rect 36952 17920 37016 17924
rect 37032 17980 37096 17984
rect 37032 17924 37036 17980
rect 37036 17924 37092 17980
rect 37092 17924 37096 17980
rect 37032 17920 37096 17924
rect 37112 17980 37176 17984
rect 37112 17924 37116 17980
rect 37116 17924 37172 17980
rect 37172 17924 37176 17980
rect 37112 17920 37176 17924
rect 37192 17980 37256 17984
rect 37192 17924 37196 17980
rect 37196 17924 37252 17980
rect 37252 17924 37256 17980
rect 37192 17920 37256 17924
rect 2612 17436 2676 17440
rect 2612 17380 2616 17436
rect 2616 17380 2672 17436
rect 2672 17380 2676 17436
rect 2612 17376 2676 17380
rect 2692 17436 2756 17440
rect 2692 17380 2696 17436
rect 2696 17380 2752 17436
rect 2752 17380 2756 17436
rect 2692 17376 2756 17380
rect 2772 17436 2836 17440
rect 2772 17380 2776 17436
rect 2776 17380 2832 17436
rect 2832 17380 2836 17436
rect 2772 17376 2836 17380
rect 2852 17436 2916 17440
rect 2852 17380 2856 17436
rect 2856 17380 2912 17436
rect 2912 17380 2916 17436
rect 2852 17376 2916 17380
rect 7612 17436 7676 17440
rect 7612 17380 7616 17436
rect 7616 17380 7672 17436
rect 7672 17380 7676 17436
rect 7612 17376 7676 17380
rect 7692 17436 7756 17440
rect 7692 17380 7696 17436
rect 7696 17380 7752 17436
rect 7752 17380 7756 17436
rect 7692 17376 7756 17380
rect 7772 17436 7836 17440
rect 7772 17380 7776 17436
rect 7776 17380 7832 17436
rect 7832 17380 7836 17436
rect 7772 17376 7836 17380
rect 7852 17436 7916 17440
rect 7852 17380 7856 17436
rect 7856 17380 7912 17436
rect 7912 17380 7916 17436
rect 7852 17376 7916 17380
rect 12612 17436 12676 17440
rect 12612 17380 12616 17436
rect 12616 17380 12672 17436
rect 12672 17380 12676 17436
rect 12612 17376 12676 17380
rect 12692 17436 12756 17440
rect 12692 17380 12696 17436
rect 12696 17380 12752 17436
rect 12752 17380 12756 17436
rect 12692 17376 12756 17380
rect 12772 17436 12836 17440
rect 12772 17380 12776 17436
rect 12776 17380 12832 17436
rect 12832 17380 12836 17436
rect 12772 17376 12836 17380
rect 12852 17436 12916 17440
rect 12852 17380 12856 17436
rect 12856 17380 12912 17436
rect 12912 17380 12916 17436
rect 12852 17376 12916 17380
rect 17612 17436 17676 17440
rect 17612 17380 17616 17436
rect 17616 17380 17672 17436
rect 17672 17380 17676 17436
rect 17612 17376 17676 17380
rect 17692 17436 17756 17440
rect 17692 17380 17696 17436
rect 17696 17380 17752 17436
rect 17752 17380 17756 17436
rect 17692 17376 17756 17380
rect 17772 17436 17836 17440
rect 17772 17380 17776 17436
rect 17776 17380 17832 17436
rect 17832 17380 17836 17436
rect 17772 17376 17836 17380
rect 17852 17436 17916 17440
rect 17852 17380 17856 17436
rect 17856 17380 17912 17436
rect 17912 17380 17916 17436
rect 17852 17376 17916 17380
rect 22612 17436 22676 17440
rect 22612 17380 22616 17436
rect 22616 17380 22672 17436
rect 22672 17380 22676 17436
rect 22612 17376 22676 17380
rect 22692 17436 22756 17440
rect 22692 17380 22696 17436
rect 22696 17380 22752 17436
rect 22752 17380 22756 17436
rect 22692 17376 22756 17380
rect 22772 17436 22836 17440
rect 22772 17380 22776 17436
rect 22776 17380 22832 17436
rect 22832 17380 22836 17436
rect 22772 17376 22836 17380
rect 22852 17436 22916 17440
rect 22852 17380 22856 17436
rect 22856 17380 22912 17436
rect 22912 17380 22916 17436
rect 22852 17376 22916 17380
rect 27612 17436 27676 17440
rect 27612 17380 27616 17436
rect 27616 17380 27672 17436
rect 27672 17380 27676 17436
rect 27612 17376 27676 17380
rect 27692 17436 27756 17440
rect 27692 17380 27696 17436
rect 27696 17380 27752 17436
rect 27752 17380 27756 17436
rect 27692 17376 27756 17380
rect 27772 17436 27836 17440
rect 27772 17380 27776 17436
rect 27776 17380 27832 17436
rect 27832 17380 27836 17436
rect 27772 17376 27836 17380
rect 27852 17436 27916 17440
rect 27852 17380 27856 17436
rect 27856 17380 27912 17436
rect 27912 17380 27916 17436
rect 27852 17376 27916 17380
rect 32612 17436 32676 17440
rect 32612 17380 32616 17436
rect 32616 17380 32672 17436
rect 32672 17380 32676 17436
rect 32612 17376 32676 17380
rect 32692 17436 32756 17440
rect 32692 17380 32696 17436
rect 32696 17380 32752 17436
rect 32752 17380 32756 17436
rect 32692 17376 32756 17380
rect 32772 17436 32836 17440
rect 32772 17380 32776 17436
rect 32776 17380 32832 17436
rect 32832 17380 32836 17436
rect 32772 17376 32836 17380
rect 32852 17436 32916 17440
rect 32852 17380 32856 17436
rect 32856 17380 32912 17436
rect 32912 17380 32916 17436
rect 32852 17376 32916 17380
rect 37612 17436 37676 17440
rect 37612 17380 37616 17436
rect 37616 17380 37672 17436
rect 37672 17380 37676 17436
rect 37612 17376 37676 17380
rect 37692 17436 37756 17440
rect 37692 17380 37696 17436
rect 37696 17380 37752 17436
rect 37752 17380 37756 17436
rect 37692 17376 37756 17380
rect 37772 17436 37836 17440
rect 37772 17380 37776 17436
rect 37776 17380 37832 17436
rect 37832 17380 37836 17436
rect 37772 17376 37836 17380
rect 37852 17436 37916 17440
rect 37852 17380 37856 17436
rect 37856 17380 37912 17436
rect 37912 17380 37916 17436
rect 37852 17376 37916 17380
rect 1952 16892 2016 16896
rect 1952 16836 1956 16892
rect 1956 16836 2012 16892
rect 2012 16836 2016 16892
rect 1952 16832 2016 16836
rect 2032 16892 2096 16896
rect 2032 16836 2036 16892
rect 2036 16836 2092 16892
rect 2092 16836 2096 16892
rect 2032 16832 2096 16836
rect 2112 16892 2176 16896
rect 2112 16836 2116 16892
rect 2116 16836 2172 16892
rect 2172 16836 2176 16892
rect 2112 16832 2176 16836
rect 2192 16892 2256 16896
rect 2192 16836 2196 16892
rect 2196 16836 2252 16892
rect 2252 16836 2256 16892
rect 2192 16832 2256 16836
rect 6952 16892 7016 16896
rect 6952 16836 6956 16892
rect 6956 16836 7012 16892
rect 7012 16836 7016 16892
rect 6952 16832 7016 16836
rect 7032 16892 7096 16896
rect 7032 16836 7036 16892
rect 7036 16836 7092 16892
rect 7092 16836 7096 16892
rect 7032 16832 7096 16836
rect 7112 16892 7176 16896
rect 7112 16836 7116 16892
rect 7116 16836 7172 16892
rect 7172 16836 7176 16892
rect 7112 16832 7176 16836
rect 7192 16892 7256 16896
rect 7192 16836 7196 16892
rect 7196 16836 7252 16892
rect 7252 16836 7256 16892
rect 7192 16832 7256 16836
rect 11952 16892 12016 16896
rect 11952 16836 11956 16892
rect 11956 16836 12012 16892
rect 12012 16836 12016 16892
rect 11952 16832 12016 16836
rect 12032 16892 12096 16896
rect 12032 16836 12036 16892
rect 12036 16836 12092 16892
rect 12092 16836 12096 16892
rect 12032 16832 12096 16836
rect 12112 16892 12176 16896
rect 12112 16836 12116 16892
rect 12116 16836 12172 16892
rect 12172 16836 12176 16892
rect 12112 16832 12176 16836
rect 12192 16892 12256 16896
rect 12192 16836 12196 16892
rect 12196 16836 12252 16892
rect 12252 16836 12256 16892
rect 12192 16832 12256 16836
rect 16952 16892 17016 16896
rect 16952 16836 16956 16892
rect 16956 16836 17012 16892
rect 17012 16836 17016 16892
rect 16952 16832 17016 16836
rect 17032 16892 17096 16896
rect 17032 16836 17036 16892
rect 17036 16836 17092 16892
rect 17092 16836 17096 16892
rect 17032 16832 17096 16836
rect 17112 16892 17176 16896
rect 17112 16836 17116 16892
rect 17116 16836 17172 16892
rect 17172 16836 17176 16892
rect 17112 16832 17176 16836
rect 17192 16892 17256 16896
rect 17192 16836 17196 16892
rect 17196 16836 17252 16892
rect 17252 16836 17256 16892
rect 17192 16832 17256 16836
rect 21952 16892 22016 16896
rect 21952 16836 21956 16892
rect 21956 16836 22012 16892
rect 22012 16836 22016 16892
rect 21952 16832 22016 16836
rect 22032 16892 22096 16896
rect 22032 16836 22036 16892
rect 22036 16836 22092 16892
rect 22092 16836 22096 16892
rect 22032 16832 22096 16836
rect 22112 16892 22176 16896
rect 22112 16836 22116 16892
rect 22116 16836 22172 16892
rect 22172 16836 22176 16892
rect 22112 16832 22176 16836
rect 22192 16892 22256 16896
rect 22192 16836 22196 16892
rect 22196 16836 22252 16892
rect 22252 16836 22256 16892
rect 22192 16832 22256 16836
rect 26952 16892 27016 16896
rect 26952 16836 26956 16892
rect 26956 16836 27012 16892
rect 27012 16836 27016 16892
rect 26952 16832 27016 16836
rect 27032 16892 27096 16896
rect 27032 16836 27036 16892
rect 27036 16836 27092 16892
rect 27092 16836 27096 16892
rect 27032 16832 27096 16836
rect 27112 16892 27176 16896
rect 27112 16836 27116 16892
rect 27116 16836 27172 16892
rect 27172 16836 27176 16892
rect 27112 16832 27176 16836
rect 27192 16892 27256 16896
rect 27192 16836 27196 16892
rect 27196 16836 27252 16892
rect 27252 16836 27256 16892
rect 27192 16832 27256 16836
rect 31952 16892 32016 16896
rect 31952 16836 31956 16892
rect 31956 16836 32012 16892
rect 32012 16836 32016 16892
rect 31952 16832 32016 16836
rect 32032 16892 32096 16896
rect 32032 16836 32036 16892
rect 32036 16836 32092 16892
rect 32092 16836 32096 16892
rect 32032 16832 32096 16836
rect 32112 16892 32176 16896
rect 32112 16836 32116 16892
rect 32116 16836 32172 16892
rect 32172 16836 32176 16892
rect 32112 16832 32176 16836
rect 32192 16892 32256 16896
rect 32192 16836 32196 16892
rect 32196 16836 32252 16892
rect 32252 16836 32256 16892
rect 32192 16832 32256 16836
rect 36952 16892 37016 16896
rect 36952 16836 36956 16892
rect 36956 16836 37012 16892
rect 37012 16836 37016 16892
rect 36952 16832 37016 16836
rect 37032 16892 37096 16896
rect 37032 16836 37036 16892
rect 37036 16836 37092 16892
rect 37092 16836 37096 16892
rect 37032 16832 37096 16836
rect 37112 16892 37176 16896
rect 37112 16836 37116 16892
rect 37116 16836 37172 16892
rect 37172 16836 37176 16892
rect 37112 16832 37176 16836
rect 37192 16892 37256 16896
rect 37192 16836 37196 16892
rect 37196 16836 37252 16892
rect 37252 16836 37256 16892
rect 37192 16832 37256 16836
rect 2612 16348 2676 16352
rect 2612 16292 2616 16348
rect 2616 16292 2672 16348
rect 2672 16292 2676 16348
rect 2612 16288 2676 16292
rect 2692 16348 2756 16352
rect 2692 16292 2696 16348
rect 2696 16292 2752 16348
rect 2752 16292 2756 16348
rect 2692 16288 2756 16292
rect 2772 16348 2836 16352
rect 2772 16292 2776 16348
rect 2776 16292 2832 16348
rect 2832 16292 2836 16348
rect 2772 16288 2836 16292
rect 2852 16348 2916 16352
rect 2852 16292 2856 16348
rect 2856 16292 2912 16348
rect 2912 16292 2916 16348
rect 2852 16288 2916 16292
rect 7612 16348 7676 16352
rect 7612 16292 7616 16348
rect 7616 16292 7672 16348
rect 7672 16292 7676 16348
rect 7612 16288 7676 16292
rect 7692 16348 7756 16352
rect 7692 16292 7696 16348
rect 7696 16292 7752 16348
rect 7752 16292 7756 16348
rect 7692 16288 7756 16292
rect 7772 16348 7836 16352
rect 7772 16292 7776 16348
rect 7776 16292 7832 16348
rect 7832 16292 7836 16348
rect 7772 16288 7836 16292
rect 7852 16348 7916 16352
rect 7852 16292 7856 16348
rect 7856 16292 7912 16348
rect 7912 16292 7916 16348
rect 7852 16288 7916 16292
rect 12612 16348 12676 16352
rect 12612 16292 12616 16348
rect 12616 16292 12672 16348
rect 12672 16292 12676 16348
rect 12612 16288 12676 16292
rect 12692 16348 12756 16352
rect 12692 16292 12696 16348
rect 12696 16292 12752 16348
rect 12752 16292 12756 16348
rect 12692 16288 12756 16292
rect 12772 16348 12836 16352
rect 12772 16292 12776 16348
rect 12776 16292 12832 16348
rect 12832 16292 12836 16348
rect 12772 16288 12836 16292
rect 12852 16348 12916 16352
rect 12852 16292 12856 16348
rect 12856 16292 12912 16348
rect 12912 16292 12916 16348
rect 12852 16288 12916 16292
rect 17612 16348 17676 16352
rect 17612 16292 17616 16348
rect 17616 16292 17672 16348
rect 17672 16292 17676 16348
rect 17612 16288 17676 16292
rect 17692 16348 17756 16352
rect 17692 16292 17696 16348
rect 17696 16292 17752 16348
rect 17752 16292 17756 16348
rect 17692 16288 17756 16292
rect 17772 16348 17836 16352
rect 17772 16292 17776 16348
rect 17776 16292 17832 16348
rect 17832 16292 17836 16348
rect 17772 16288 17836 16292
rect 17852 16348 17916 16352
rect 17852 16292 17856 16348
rect 17856 16292 17912 16348
rect 17912 16292 17916 16348
rect 17852 16288 17916 16292
rect 22612 16348 22676 16352
rect 22612 16292 22616 16348
rect 22616 16292 22672 16348
rect 22672 16292 22676 16348
rect 22612 16288 22676 16292
rect 22692 16348 22756 16352
rect 22692 16292 22696 16348
rect 22696 16292 22752 16348
rect 22752 16292 22756 16348
rect 22692 16288 22756 16292
rect 22772 16348 22836 16352
rect 22772 16292 22776 16348
rect 22776 16292 22832 16348
rect 22832 16292 22836 16348
rect 22772 16288 22836 16292
rect 22852 16348 22916 16352
rect 22852 16292 22856 16348
rect 22856 16292 22912 16348
rect 22912 16292 22916 16348
rect 22852 16288 22916 16292
rect 27612 16348 27676 16352
rect 27612 16292 27616 16348
rect 27616 16292 27672 16348
rect 27672 16292 27676 16348
rect 27612 16288 27676 16292
rect 27692 16348 27756 16352
rect 27692 16292 27696 16348
rect 27696 16292 27752 16348
rect 27752 16292 27756 16348
rect 27692 16288 27756 16292
rect 27772 16348 27836 16352
rect 27772 16292 27776 16348
rect 27776 16292 27832 16348
rect 27832 16292 27836 16348
rect 27772 16288 27836 16292
rect 27852 16348 27916 16352
rect 27852 16292 27856 16348
rect 27856 16292 27912 16348
rect 27912 16292 27916 16348
rect 27852 16288 27916 16292
rect 32612 16348 32676 16352
rect 32612 16292 32616 16348
rect 32616 16292 32672 16348
rect 32672 16292 32676 16348
rect 32612 16288 32676 16292
rect 32692 16348 32756 16352
rect 32692 16292 32696 16348
rect 32696 16292 32752 16348
rect 32752 16292 32756 16348
rect 32692 16288 32756 16292
rect 32772 16348 32836 16352
rect 32772 16292 32776 16348
rect 32776 16292 32832 16348
rect 32832 16292 32836 16348
rect 32772 16288 32836 16292
rect 32852 16348 32916 16352
rect 32852 16292 32856 16348
rect 32856 16292 32912 16348
rect 32912 16292 32916 16348
rect 32852 16288 32916 16292
rect 37612 16348 37676 16352
rect 37612 16292 37616 16348
rect 37616 16292 37672 16348
rect 37672 16292 37676 16348
rect 37612 16288 37676 16292
rect 37692 16348 37756 16352
rect 37692 16292 37696 16348
rect 37696 16292 37752 16348
rect 37752 16292 37756 16348
rect 37692 16288 37756 16292
rect 37772 16348 37836 16352
rect 37772 16292 37776 16348
rect 37776 16292 37832 16348
rect 37832 16292 37836 16348
rect 37772 16288 37836 16292
rect 37852 16348 37916 16352
rect 37852 16292 37856 16348
rect 37856 16292 37912 16348
rect 37912 16292 37916 16348
rect 37852 16288 37916 16292
rect 1952 15804 2016 15808
rect 1952 15748 1956 15804
rect 1956 15748 2012 15804
rect 2012 15748 2016 15804
rect 1952 15744 2016 15748
rect 2032 15804 2096 15808
rect 2032 15748 2036 15804
rect 2036 15748 2092 15804
rect 2092 15748 2096 15804
rect 2032 15744 2096 15748
rect 2112 15804 2176 15808
rect 2112 15748 2116 15804
rect 2116 15748 2172 15804
rect 2172 15748 2176 15804
rect 2112 15744 2176 15748
rect 2192 15804 2256 15808
rect 2192 15748 2196 15804
rect 2196 15748 2252 15804
rect 2252 15748 2256 15804
rect 2192 15744 2256 15748
rect 6952 15804 7016 15808
rect 6952 15748 6956 15804
rect 6956 15748 7012 15804
rect 7012 15748 7016 15804
rect 6952 15744 7016 15748
rect 7032 15804 7096 15808
rect 7032 15748 7036 15804
rect 7036 15748 7092 15804
rect 7092 15748 7096 15804
rect 7032 15744 7096 15748
rect 7112 15804 7176 15808
rect 7112 15748 7116 15804
rect 7116 15748 7172 15804
rect 7172 15748 7176 15804
rect 7112 15744 7176 15748
rect 7192 15804 7256 15808
rect 7192 15748 7196 15804
rect 7196 15748 7252 15804
rect 7252 15748 7256 15804
rect 7192 15744 7256 15748
rect 11952 15804 12016 15808
rect 11952 15748 11956 15804
rect 11956 15748 12012 15804
rect 12012 15748 12016 15804
rect 11952 15744 12016 15748
rect 12032 15804 12096 15808
rect 12032 15748 12036 15804
rect 12036 15748 12092 15804
rect 12092 15748 12096 15804
rect 12032 15744 12096 15748
rect 12112 15804 12176 15808
rect 12112 15748 12116 15804
rect 12116 15748 12172 15804
rect 12172 15748 12176 15804
rect 12112 15744 12176 15748
rect 12192 15804 12256 15808
rect 12192 15748 12196 15804
rect 12196 15748 12252 15804
rect 12252 15748 12256 15804
rect 12192 15744 12256 15748
rect 16952 15804 17016 15808
rect 16952 15748 16956 15804
rect 16956 15748 17012 15804
rect 17012 15748 17016 15804
rect 16952 15744 17016 15748
rect 17032 15804 17096 15808
rect 17032 15748 17036 15804
rect 17036 15748 17092 15804
rect 17092 15748 17096 15804
rect 17032 15744 17096 15748
rect 17112 15804 17176 15808
rect 17112 15748 17116 15804
rect 17116 15748 17172 15804
rect 17172 15748 17176 15804
rect 17112 15744 17176 15748
rect 17192 15804 17256 15808
rect 17192 15748 17196 15804
rect 17196 15748 17252 15804
rect 17252 15748 17256 15804
rect 17192 15744 17256 15748
rect 21952 15804 22016 15808
rect 21952 15748 21956 15804
rect 21956 15748 22012 15804
rect 22012 15748 22016 15804
rect 21952 15744 22016 15748
rect 22032 15804 22096 15808
rect 22032 15748 22036 15804
rect 22036 15748 22092 15804
rect 22092 15748 22096 15804
rect 22032 15744 22096 15748
rect 22112 15804 22176 15808
rect 22112 15748 22116 15804
rect 22116 15748 22172 15804
rect 22172 15748 22176 15804
rect 22112 15744 22176 15748
rect 22192 15804 22256 15808
rect 22192 15748 22196 15804
rect 22196 15748 22252 15804
rect 22252 15748 22256 15804
rect 22192 15744 22256 15748
rect 26952 15804 27016 15808
rect 26952 15748 26956 15804
rect 26956 15748 27012 15804
rect 27012 15748 27016 15804
rect 26952 15744 27016 15748
rect 27032 15804 27096 15808
rect 27032 15748 27036 15804
rect 27036 15748 27092 15804
rect 27092 15748 27096 15804
rect 27032 15744 27096 15748
rect 27112 15804 27176 15808
rect 27112 15748 27116 15804
rect 27116 15748 27172 15804
rect 27172 15748 27176 15804
rect 27112 15744 27176 15748
rect 27192 15804 27256 15808
rect 27192 15748 27196 15804
rect 27196 15748 27252 15804
rect 27252 15748 27256 15804
rect 27192 15744 27256 15748
rect 31952 15804 32016 15808
rect 31952 15748 31956 15804
rect 31956 15748 32012 15804
rect 32012 15748 32016 15804
rect 31952 15744 32016 15748
rect 32032 15804 32096 15808
rect 32032 15748 32036 15804
rect 32036 15748 32092 15804
rect 32092 15748 32096 15804
rect 32032 15744 32096 15748
rect 32112 15804 32176 15808
rect 32112 15748 32116 15804
rect 32116 15748 32172 15804
rect 32172 15748 32176 15804
rect 32112 15744 32176 15748
rect 32192 15804 32256 15808
rect 32192 15748 32196 15804
rect 32196 15748 32252 15804
rect 32252 15748 32256 15804
rect 32192 15744 32256 15748
rect 36952 15804 37016 15808
rect 36952 15748 36956 15804
rect 36956 15748 37012 15804
rect 37012 15748 37016 15804
rect 36952 15744 37016 15748
rect 37032 15804 37096 15808
rect 37032 15748 37036 15804
rect 37036 15748 37092 15804
rect 37092 15748 37096 15804
rect 37032 15744 37096 15748
rect 37112 15804 37176 15808
rect 37112 15748 37116 15804
rect 37116 15748 37172 15804
rect 37172 15748 37176 15804
rect 37112 15744 37176 15748
rect 37192 15804 37256 15808
rect 37192 15748 37196 15804
rect 37196 15748 37252 15804
rect 37252 15748 37256 15804
rect 37192 15744 37256 15748
rect 2612 15260 2676 15264
rect 2612 15204 2616 15260
rect 2616 15204 2672 15260
rect 2672 15204 2676 15260
rect 2612 15200 2676 15204
rect 2692 15260 2756 15264
rect 2692 15204 2696 15260
rect 2696 15204 2752 15260
rect 2752 15204 2756 15260
rect 2692 15200 2756 15204
rect 2772 15260 2836 15264
rect 2772 15204 2776 15260
rect 2776 15204 2832 15260
rect 2832 15204 2836 15260
rect 2772 15200 2836 15204
rect 2852 15260 2916 15264
rect 2852 15204 2856 15260
rect 2856 15204 2912 15260
rect 2912 15204 2916 15260
rect 2852 15200 2916 15204
rect 7612 15260 7676 15264
rect 7612 15204 7616 15260
rect 7616 15204 7672 15260
rect 7672 15204 7676 15260
rect 7612 15200 7676 15204
rect 7692 15260 7756 15264
rect 7692 15204 7696 15260
rect 7696 15204 7752 15260
rect 7752 15204 7756 15260
rect 7692 15200 7756 15204
rect 7772 15260 7836 15264
rect 7772 15204 7776 15260
rect 7776 15204 7832 15260
rect 7832 15204 7836 15260
rect 7772 15200 7836 15204
rect 7852 15260 7916 15264
rect 7852 15204 7856 15260
rect 7856 15204 7912 15260
rect 7912 15204 7916 15260
rect 7852 15200 7916 15204
rect 12612 15260 12676 15264
rect 12612 15204 12616 15260
rect 12616 15204 12672 15260
rect 12672 15204 12676 15260
rect 12612 15200 12676 15204
rect 12692 15260 12756 15264
rect 12692 15204 12696 15260
rect 12696 15204 12752 15260
rect 12752 15204 12756 15260
rect 12692 15200 12756 15204
rect 12772 15260 12836 15264
rect 12772 15204 12776 15260
rect 12776 15204 12832 15260
rect 12832 15204 12836 15260
rect 12772 15200 12836 15204
rect 12852 15260 12916 15264
rect 12852 15204 12856 15260
rect 12856 15204 12912 15260
rect 12912 15204 12916 15260
rect 12852 15200 12916 15204
rect 17612 15260 17676 15264
rect 17612 15204 17616 15260
rect 17616 15204 17672 15260
rect 17672 15204 17676 15260
rect 17612 15200 17676 15204
rect 17692 15260 17756 15264
rect 17692 15204 17696 15260
rect 17696 15204 17752 15260
rect 17752 15204 17756 15260
rect 17692 15200 17756 15204
rect 17772 15260 17836 15264
rect 17772 15204 17776 15260
rect 17776 15204 17832 15260
rect 17832 15204 17836 15260
rect 17772 15200 17836 15204
rect 17852 15260 17916 15264
rect 17852 15204 17856 15260
rect 17856 15204 17912 15260
rect 17912 15204 17916 15260
rect 17852 15200 17916 15204
rect 22612 15260 22676 15264
rect 22612 15204 22616 15260
rect 22616 15204 22672 15260
rect 22672 15204 22676 15260
rect 22612 15200 22676 15204
rect 22692 15260 22756 15264
rect 22692 15204 22696 15260
rect 22696 15204 22752 15260
rect 22752 15204 22756 15260
rect 22692 15200 22756 15204
rect 22772 15260 22836 15264
rect 22772 15204 22776 15260
rect 22776 15204 22832 15260
rect 22832 15204 22836 15260
rect 22772 15200 22836 15204
rect 22852 15260 22916 15264
rect 22852 15204 22856 15260
rect 22856 15204 22912 15260
rect 22912 15204 22916 15260
rect 22852 15200 22916 15204
rect 27612 15260 27676 15264
rect 27612 15204 27616 15260
rect 27616 15204 27672 15260
rect 27672 15204 27676 15260
rect 27612 15200 27676 15204
rect 27692 15260 27756 15264
rect 27692 15204 27696 15260
rect 27696 15204 27752 15260
rect 27752 15204 27756 15260
rect 27692 15200 27756 15204
rect 27772 15260 27836 15264
rect 27772 15204 27776 15260
rect 27776 15204 27832 15260
rect 27832 15204 27836 15260
rect 27772 15200 27836 15204
rect 27852 15260 27916 15264
rect 27852 15204 27856 15260
rect 27856 15204 27912 15260
rect 27912 15204 27916 15260
rect 27852 15200 27916 15204
rect 32612 15260 32676 15264
rect 32612 15204 32616 15260
rect 32616 15204 32672 15260
rect 32672 15204 32676 15260
rect 32612 15200 32676 15204
rect 32692 15260 32756 15264
rect 32692 15204 32696 15260
rect 32696 15204 32752 15260
rect 32752 15204 32756 15260
rect 32692 15200 32756 15204
rect 32772 15260 32836 15264
rect 32772 15204 32776 15260
rect 32776 15204 32832 15260
rect 32832 15204 32836 15260
rect 32772 15200 32836 15204
rect 32852 15260 32916 15264
rect 32852 15204 32856 15260
rect 32856 15204 32912 15260
rect 32912 15204 32916 15260
rect 32852 15200 32916 15204
rect 37612 15260 37676 15264
rect 37612 15204 37616 15260
rect 37616 15204 37672 15260
rect 37672 15204 37676 15260
rect 37612 15200 37676 15204
rect 37692 15260 37756 15264
rect 37692 15204 37696 15260
rect 37696 15204 37752 15260
rect 37752 15204 37756 15260
rect 37692 15200 37756 15204
rect 37772 15260 37836 15264
rect 37772 15204 37776 15260
rect 37776 15204 37832 15260
rect 37832 15204 37836 15260
rect 37772 15200 37836 15204
rect 37852 15260 37916 15264
rect 37852 15204 37856 15260
rect 37856 15204 37912 15260
rect 37912 15204 37916 15260
rect 37852 15200 37916 15204
rect 24900 14996 24964 15060
rect 1952 14716 2016 14720
rect 1952 14660 1956 14716
rect 1956 14660 2012 14716
rect 2012 14660 2016 14716
rect 1952 14656 2016 14660
rect 2032 14716 2096 14720
rect 2032 14660 2036 14716
rect 2036 14660 2092 14716
rect 2092 14660 2096 14716
rect 2032 14656 2096 14660
rect 2112 14716 2176 14720
rect 2112 14660 2116 14716
rect 2116 14660 2172 14716
rect 2172 14660 2176 14716
rect 2112 14656 2176 14660
rect 2192 14716 2256 14720
rect 2192 14660 2196 14716
rect 2196 14660 2252 14716
rect 2252 14660 2256 14716
rect 2192 14656 2256 14660
rect 6952 14716 7016 14720
rect 6952 14660 6956 14716
rect 6956 14660 7012 14716
rect 7012 14660 7016 14716
rect 6952 14656 7016 14660
rect 7032 14716 7096 14720
rect 7032 14660 7036 14716
rect 7036 14660 7092 14716
rect 7092 14660 7096 14716
rect 7032 14656 7096 14660
rect 7112 14716 7176 14720
rect 7112 14660 7116 14716
rect 7116 14660 7172 14716
rect 7172 14660 7176 14716
rect 7112 14656 7176 14660
rect 7192 14716 7256 14720
rect 7192 14660 7196 14716
rect 7196 14660 7252 14716
rect 7252 14660 7256 14716
rect 7192 14656 7256 14660
rect 11952 14716 12016 14720
rect 11952 14660 11956 14716
rect 11956 14660 12012 14716
rect 12012 14660 12016 14716
rect 11952 14656 12016 14660
rect 12032 14716 12096 14720
rect 12032 14660 12036 14716
rect 12036 14660 12092 14716
rect 12092 14660 12096 14716
rect 12032 14656 12096 14660
rect 12112 14716 12176 14720
rect 12112 14660 12116 14716
rect 12116 14660 12172 14716
rect 12172 14660 12176 14716
rect 12112 14656 12176 14660
rect 12192 14716 12256 14720
rect 12192 14660 12196 14716
rect 12196 14660 12252 14716
rect 12252 14660 12256 14716
rect 12192 14656 12256 14660
rect 16952 14716 17016 14720
rect 16952 14660 16956 14716
rect 16956 14660 17012 14716
rect 17012 14660 17016 14716
rect 16952 14656 17016 14660
rect 17032 14716 17096 14720
rect 17032 14660 17036 14716
rect 17036 14660 17092 14716
rect 17092 14660 17096 14716
rect 17032 14656 17096 14660
rect 17112 14716 17176 14720
rect 17112 14660 17116 14716
rect 17116 14660 17172 14716
rect 17172 14660 17176 14716
rect 17112 14656 17176 14660
rect 17192 14716 17256 14720
rect 17192 14660 17196 14716
rect 17196 14660 17252 14716
rect 17252 14660 17256 14716
rect 17192 14656 17256 14660
rect 21952 14716 22016 14720
rect 21952 14660 21956 14716
rect 21956 14660 22012 14716
rect 22012 14660 22016 14716
rect 21952 14656 22016 14660
rect 22032 14716 22096 14720
rect 22032 14660 22036 14716
rect 22036 14660 22092 14716
rect 22092 14660 22096 14716
rect 22032 14656 22096 14660
rect 22112 14716 22176 14720
rect 22112 14660 22116 14716
rect 22116 14660 22172 14716
rect 22172 14660 22176 14716
rect 22112 14656 22176 14660
rect 22192 14716 22256 14720
rect 22192 14660 22196 14716
rect 22196 14660 22252 14716
rect 22252 14660 22256 14716
rect 22192 14656 22256 14660
rect 26952 14716 27016 14720
rect 26952 14660 26956 14716
rect 26956 14660 27012 14716
rect 27012 14660 27016 14716
rect 26952 14656 27016 14660
rect 27032 14716 27096 14720
rect 27032 14660 27036 14716
rect 27036 14660 27092 14716
rect 27092 14660 27096 14716
rect 27032 14656 27096 14660
rect 27112 14716 27176 14720
rect 27112 14660 27116 14716
rect 27116 14660 27172 14716
rect 27172 14660 27176 14716
rect 27112 14656 27176 14660
rect 27192 14716 27256 14720
rect 27192 14660 27196 14716
rect 27196 14660 27252 14716
rect 27252 14660 27256 14716
rect 27192 14656 27256 14660
rect 31952 14716 32016 14720
rect 31952 14660 31956 14716
rect 31956 14660 32012 14716
rect 32012 14660 32016 14716
rect 31952 14656 32016 14660
rect 32032 14716 32096 14720
rect 32032 14660 32036 14716
rect 32036 14660 32092 14716
rect 32092 14660 32096 14716
rect 32032 14656 32096 14660
rect 32112 14716 32176 14720
rect 32112 14660 32116 14716
rect 32116 14660 32172 14716
rect 32172 14660 32176 14716
rect 32112 14656 32176 14660
rect 32192 14716 32256 14720
rect 32192 14660 32196 14716
rect 32196 14660 32252 14716
rect 32252 14660 32256 14716
rect 32192 14656 32256 14660
rect 36952 14716 37016 14720
rect 36952 14660 36956 14716
rect 36956 14660 37012 14716
rect 37012 14660 37016 14716
rect 36952 14656 37016 14660
rect 37032 14716 37096 14720
rect 37032 14660 37036 14716
rect 37036 14660 37092 14716
rect 37092 14660 37096 14716
rect 37032 14656 37096 14660
rect 37112 14716 37176 14720
rect 37112 14660 37116 14716
rect 37116 14660 37172 14716
rect 37172 14660 37176 14716
rect 37112 14656 37176 14660
rect 37192 14716 37256 14720
rect 37192 14660 37196 14716
rect 37196 14660 37252 14716
rect 37252 14660 37256 14716
rect 37192 14656 37256 14660
rect 2612 14172 2676 14176
rect 2612 14116 2616 14172
rect 2616 14116 2672 14172
rect 2672 14116 2676 14172
rect 2612 14112 2676 14116
rect 2692 14172 2756 14176
rect 2692 14116 2696 14172
rect 2696 14116 2752 14172
rect 2752 14116 2756 14172
rect 2692 14112 2756 14116
rect 2772 14172 2836 14176
rect 2772 14116 2776 14172
rect 2776 14116 2832 14172
rect 2832 14116 2836 14172
rect 2772 14112 2836 14116
rect 2852 14172 2916 14176
rect 2852 14116 2856 14172
rect 2856 14116 2912 14172
rect 2912 14116 2916 14172
rect 2852 14112 2916 14116
rect 7612 14172 7676 14176
rect 7612 14116 7616 14172
rect 7616 14116 7672 14172
rect 7672 14116 7676 14172
rect 7612 14112 7676 14116
rect 7692 14172 7756 14176
rect 7692 14116 7696 14172
rect 7696 14116 7752 14172
rect 7752 14116 7756 14172
rect 7692 14112 7756 14116
rect 7772 14172 7836 14176
rect 7772 14116 7776 14172
rect 7776 14116 7832 14172
rect 7832 14116 7836 14172
rect 7772 14112 7836 14116
rect 7852 14172 7916 14176
rect 7852 14116 7856 14172
rect 7856 14116 7912 14172
rect 7912 14116 7916 14172
rect 7852 14112 7916 14116
rect 12612 14172 12676 14176
rect 12612 14116 12616 14172
rect 12616 14116 12672 14172
rect 12672 14116 12676 14172
rect 12612 14112 12676 14116
rect 12692 14172 12756 14176
rect 12692 14116 12696 14172
rect 12696 14116 12752 14172
rect 12752 14116 12756 14172
rect 12692 14112 12756 14116
rect 12772 14172 12836 14176
rect 12772 14116 12776 14172
rect 12776 14116 12832 14172
rect 12832 14116 12836 14172
rect 12772 14112 12836 14116
rect 12852 14172 12916 14176
rect 12852 14116 12856 14172
rect 12856 14116 12912 14172
rect 12912 14116 12916 14172
rect 12852 14112 12916 14116
rect 17612 14172 17676 14176
rect 17612 14116 17616 14172
rect 17616 14116 17672 14172
rect 17672 14116 17676 14172
rect 17612 14112 17676 14116
rect 17692 14172 17756 14176
rect 17692 14116 17696 14172
rect 17696 14116 17752 14172
rect 17752 14116 17756 14172
rect 17692 14112 17756 14116
rect 17772 14172 17836 14176
rect 17772 14116 17776 14172
rect 17776 14116 17832 14172
rect 17832 14116 17836 14172
rect 17772 14112 17836 14116
rect 17852 14172 17916 14176
rect 17852 14116 17856 14172
rect 17856 14116 17912 14172
rect 17912 14116 17916 14172
rect 17852 14112 17916 14116
rect 22612 14172 22676 14176
rect 22612 14116 22616 14172
rect 22616 14116 22672 14172
rect 22672 14116 22676 14172
rect 22612 14112 22676 14116
rect 22692 14172 22756 14176
rect 22692 14116 22696 14172
rect 22696 14116 22752 14172
rect 22752 14116 22756 14172
rect 22692 14112 22756 14116
rect 22772 14172 22836 14176
rect 22772 14116 22776 14172
rect 22776 14116 22832 14172
rect 22832 14116 22836 14172
rect 22772 14112 22836 14116
rect 22852 14172 22916 14176
rect 22852 14116 22856 14172
rect 22856 14116 22912 14172
rect 22912 14116 22916 14172
rect 22852 14112 22916 14116
rect 27612 14172 27676 14176
rect 27612 14116 27616 14172
rect 27616 14116 27672 14172
rect 27672 14116 27676 14172
rect 27612 14112 27676 14116
rect 27692 14172 27756 14176
rect 27692 14116 27696 14172
rect 27696 14116 27752 14172
rect 27752 14116 27756 14172
rect 27692 14112 27756 14116
rect 27772 14172 27836 14176
rect 27772 14116 27776 14172
rect 27776 14116 27832 14172
rect 27832 14116 27836 14172
rect 27772 14112 27836 14116
rect 27852 14172 27916 14176
rect 27852 14116 27856 14172
rect 27856 14116 27912 14172
rect 27912 14116 27916 14172
rect 27852 14112 27916 14116
rect 32612 14172 32676 14176
rect 32612 14116 32616 14172
rect 32616 14116 32672 14172
rect 32672 14116 32676 14172
rect 32612 14112 32676 14116
rect 32692 14172 32756 14176
rect 32692 14116 32696 14172
rect 32696 14116 32752 14172
rect 32752 14116 32756 14172
rect 32692 14112 32756 14116
rect 32772 14172 32836 14176
rect 32772 14116 32776 14172
rect 32776 14116 32832 14172
rect 32832 14116 32836 14172
rect 32772 14112 32836 14116
rect 32852 14172 32916 14176
rect 32852 14116 32856 14172
rect 32856 14116 32912 14172
rect 32912 14116 32916 14172
rect 32852 14112 32916 14116
rect 37612 14172 37676 14176
rect 37612 14116 37616 14172
rect 37616 14116 37672 14172
rect 37672 14116 37676 14172
rect 37612 14112 37676 14116
rect 37692 14172 37756 14176
rect 37692 14116 37696 14172
rect 37696 14116 37752 14172
rect 37752 14116 37756 14172
rect 37692 14112 37756 14116
rect 37772 14172 37836 14176
rect 37772 14116 37776 14172
rect 37776 14116 37832 14172
rect 37832 14116 37836 14172
rect 37772 14112 37836 14116
rect 37852 14172 37916 14176
rect 37852 14116 37856 14172
rect 37856 14116 37912 14172
rect 37912 14116 37916 14172
rect 37852 14112 37916 14116
rect 1952 13628 2016 13632
rect 1952 13572 1956 13628
rect 1956 13572 2012 13628
rect 2012 13572 2016 13628
rect 1952 13568 2016 13572
rect 2032 13628 2096 13632
rect 2032 13572 2036 13628
rect 2036 13572 2092 13628
rect 2092 13572 2096 13628
rect 2032 13568 2096 13572
rect 2112 13628 2176 13632
rect 2112 13572 2116 13628
rect 2116 13572 2172 13628
rect 2172 13572 2176 13628
rect 2112 13568 2176 13572
rect 2192 13628 2256 13632
rect 2192 13572 2196 13628
rect 2196 13572 2252 13628
rect 2252 13572 2256 13628
rect 2192 13568 2256 13572
rect 6952 13628 7016 13632
rect 6952 13572 6956 13628
rect 6956 13572 7012 13628
rect 7012 13572 7016 13628
rect 6952 13568 7016 13572
rect 7032 13628 7096 13632
rect 7032 13572 7036 13628
rect 7036 13572 7092 13628
rect 7092 13572 7096 13628
rect 7032 13568 7096 13572
rect 7112 13628 7176 13632
rect 7112 13572 7116 13628
rect 7116 13572 7172 13628
rect 7172 13572 7176 13628
rect 7112 13568 7176 13572
rect 7192 13628 7256 13632
rect 7192 13572 7196 13628
rect 7196 13572 7252 13628
rect 7252 13572 7256 13628
rect 7192 13568 7256 13572
rect 11952 13628 12016 13632
rect 11952 13572 11956 13628
rect 11956 13572 12012 13628
rect 12012 13572 12016 13628
rect 11952 13568 12016 13572
rect 12032 13628 12096 13632
rect 12032 13572 12036 13628
rect 12036 13572 12092 13628
rect 12092 13572 12096 13628
rect 12032 13568 12096 13572
rect 12112 13628 12176 13632
rect 12112 13572 12116 13628
rect 12116 13572 12172 13628
rect 12172 13572 12176 13628
rect 12112 13568 12176 13572
rect 12192 13628 12256 13632
rect 12192 13572 12196 13628
rect 12196 13572 12252 13628
rect 12252 13572 12256 13628
rect 12192 13568 12256 13572
rect 16952 13628 17016 13632
rect 16952 13572 16956 13628
rect 16956 13572 17012 13628
rect 17012 13572 17016 13628
rect 16952 13568 17016 13572
rect 17032 13628 17096 13632
rect 17032 13572 17036 13628
rect 17036 13572 17092 13628
rect 17092 13572 17096 13628
rect 17032 13568 17096 13572
rect 17112 13628 17176 13632
rect 17112 13572 17116 13628
rect 17116 13572 17172 13628
rect 17172 13572 17176 13628
rect 17112 13568 17176 13572
rect 17192 13628 17256 13632
rect 17192 13572 17196 13628
rect 17196 13572 17252 13628
rect 17252 13572 17256 13628
rect 17192 13568 17256 13572
rect 21952 13628 22016 13632
rect 21952 13572 21956 13628
rect 21956 13572 22012 13628
rect 22012 13572 22016 13628
rect 21952 13568 22016 13572
rect 22032 13628 22096 13632
rect 22032 13572 22036 13628
rect 22036 13572 22092 13628
rect 22092 13572 22096 13628
rect 22032 13568 22096 13572
rect 22112 13628 22176 13632
rect 22112 13572 22116 13628
rect 22116 13572 22172 13628
rect 22172 13572 22176 13628
rect 22112 13568 22176 13572
rect 22192 13628 22256 13632
rect 22192 13572 22196 13628
rect 22196 13572 22252 13628
rect 22252 13572 22256 13628
rect 22192 13568 22256 13572
rect 26952 13628 27016 13632
rect 26952 13572 26956 13628
rect 26956 13572 27012 13628
rect 27012 13572 27016 13628
rect 26952 13568 27016 13572
rect 27032 13628 27096 13632
rect 27032 13572 27036 13628
rect 27036 13572 27092 13628
rect 27092 13572 27096 13628
rect 27032 13568 27096 13572
rect 27112 13628 27176 13632
rect 27112 13572 27116 13628
rect 27116 13572 27172 13628
rect 27172 13572 27176 13628
rect 27112 13568 27176 13572
rect 27192 13628 27256 13632
rect 27192 13572 27196 13628
rect 27196 13572 27252 13628
rect 27252 13572 27256 13628
rect 27192 13568 27256 13572
rect 31952 13628 32016 13632
rect 31952 13572 31956 13628
rect 31956 13572 32012 13628
rect 32012 13572 32016 13628
rect 31952 13568 32016 13572
rect 32032 13628 32096 13632
rect 32032 13572 32036 13628
rect 32036 13572 32092 13628
rect 32092 13572 32096 13628
rect 32032 13568 32096 13572
rect 32112 13628 32176 13632
rect 32112 13572 32116 13628
rect 32116 13572 32172 13628
rect 32172 13572 32176 13628
rect 32112 13568 32176 13572
rect 32192 13628 32256 13632
rect 32192 13572 32196 13628
rect 32196 13572 32252 13628
rect 32252 13572 32256 13628
rect 32192 13568 32256 13572
rect 36952 13628 37016 13632
rect 36952 13572 36956 13628
rect 36956 13572 37012 13628
rect 37012 13572 37016 13628
rect 36952 13568 37016 13572
rect 37032 13628 37096 13632
rect 37032 13572 37036 13628
rect 37036 13572 37092 13628
rect 37092 13572 37096 13628
rect 37032 13568 37096 13572
rect 37112 13628 37176 13632
rect 37112 13572 37116 13628
rect 37116 13572 37172 13628
rect 37172 13572 37176 13628
rect 37112 13568 37176 13572
rect 37192 13628 37256 13632
rect 37192 13572 37196 13628
rect 37196 13572 37252 13628
rect 37252 13572 37256 13628
rect 37192 13568 37256 13572
rect 21588 13364 21652 13428
rect 2612 13084 2676 13088
rect 2612 13028 2616 13084
rect 2616 13028 2672 13084
rect 2672 13028 2676 13084
rect 2612 13024 2676 13028
rect 2692 13084 2756 13088
rect 2692 13028 2696 13084
rect 2696 13028 2752 13084
rect 2752 13028 2756 13084
rect 2692 13024 2756 13028
rect 2772 13084 2836 13088
rect 2772 13028 2776 13084
rect 2776 13028 2832 13084
rect 2832 13028 2836 13084
rect 2772 13024 2836 13028
rect 2852 13084 2916 13088
rect 2852 13028 2856 13084
rect 2856 13028 2912 13084
rect 2912 13028 2916 13084
rect 2852 13024 2916 13028
rect 7612 13084 7676 13088
rect 7612 13028 7616 13084
rect 7616 13028 7672 13084
rect 7672 13028 7676 13084
rect 7612 13024 7676 13028
rect 7692 13084 7756 13088
rect 7692 13028 7696 13084
rect 7696 13028 7752 13084
rect 7752 13028 7756 13084
rect 7692 13024 7756 13028
rect 7772 13084 7836 13088
rect 7772 13028 7776 13084
rect 7776 13028 7832 13084
rect 7832 13028 7836 13084
rect 7772 13024 7836 13028
rect 7852 13084 7916 13088
rect 7852 13028 7856 13084
rect 7856 13028 7912 13084
rect 7912 13028 7916 13084
rect 7852 13024 7916 13028
rect 12612 13084 12676 13088
rect 12612 13028 12616 13084
rect 12616 13028 12672 13084
rect 12672 13028 12676 13084
rect 12612 13024 12676 13028
rect 12692 13084 12756 13088
rect 12692 13028 12696 13084
rect 12696 13028 12752 13084
rect 12752 13028 12756 13084
rect 12692 13024 12756 13028
rect 12772 13084 12836 13088
rect 12772 13028 12776 13084
rect 12776 13028 12832 13084
rect 12832 13028 12836 13084
rect 12772 13024 12836 13028
rect 12852 13084 12916 13088
rect 12852 13028 12856 13084
rect 12856 13028 12912 13084
rect 12912 13028 12916 13084
rect 12852 13024 12916 13028
rect 17612 13084 17676 13088
rect 17612 13028 17616 13084
rect 17616 13028 17672 13084
rect 17672 13028 17676 13084
rect 17612 13024 17676 13028
rect 17692 13084 17756 13088
rect 17692 13028 17696 13084
rect 17696 13028 17752 13084
rect 17752 13028 17756 13084
rect 17692 13024 17756 13028
rect 17772 13084 17836 13088
rect 17772 13028 17776 13084
rect 17776 13028 17832 13084
rect 17832 13028 17836 13084
rect 17772 13024 17836 13028
rect 17852 13084 17916 13088
rect 17852 13028 17856 13084
rect 17856 13028 17912 13084
rect 17912 13028 17916 13084
rect 17852 13024 17916 13028
rect 22612 13084 22676 13088
rect 22612 13028 22616 13084
rect 22616 13028 22672 13084
rect 22672 13028 22676 13084
rect 22612 13024 22676 13028
rect 22692 13084 22756 13088
rect 22692 13028 22696 13084
rect 22696 13028 22752 13084
rect 22752 13028 22756 13084
rect 22692 13024 22756 13028
rect 22772 13084 22836 13088
rect 22772 13028 22776 13084
rect 22776 13028 22832 13084
rect 22832 13028 22836 13084
rect 22772 13024 22836 13028
rect 22852 13084 22916 13088
rect 22852 13028 22856 13084
rect 22856 13028 22912 13084
rect 22912 13028 22916 13084
rect 22852 13024 22916 13028
rect 27612 13084 27676 13088
rect 27612 13028 27616 13084
rect 27616 13028 27672 13084
rect 27672 13028 27676 13084
rect 27612 13024 27676 13028
rect 27692 13084 27756 13088
rect 27692 13028 27696 13084
rect 27696 13028 27752 13084
rect 27752 13028 27756 13084
rect 27692 13024 27756 13028
rect 27772 13084 27836 13088
rect 27772 13028 27776 13084
rect 27776 13028 27832 13084
rect 27832 13028 27836 13084
rect 27772 13024 27836 13028
rect 27852 13084 27916 13088
rect 27852 13028 27856 13084
rect 27856 13028 27912 13084
rect 27912 13028 27916 13084
rect 27852 13024 27916 13028
rect 32612 13084 32676 13088
rect 32612 13028 32616 13084
rect 32616 13028 32672 13084
rect 32672 13028 32676 13084
rect 32612 13024 32676 13028
rect 32692 13084 32756 13088
rect 32692 13028 32696 13084
rect 32696 13028 32752 13084
rect 32752 13028 32756 13084
rect 32692 13024 32756 13028
rect 32772 13084 32836 13088
rect 32772 13028 32776 13084
rect 32776 13028 32832 13084
rect 32832 13028 32836 13084
rect 32772 13024 32836 13028
rect 32852 13084 32916 13088
rect 32852 13028 32856 13084
rect 32856 13028 32912 13084
rect 32912 13028 32916 13084
rect 32852 13024 32916 13028
rect 37612 13084 37676 13088
rect 37612 13028 37616 13084
rect 37616 13028 37672 13084
rect 37672 13028 37676 13084
rect 37612 13024 37676 13028
rect 37692 13084 37756 13088
rect 37692 13028 37696 13084
rect 37696 13028 37752 13084
rect 37752 13028 37756 13084
rect 37692 13024 37756 13028
rect 37772 13084 37836 13088
rect 37772 13028 37776 13084
rect 37776 13028 37832 13084
rect 37832 13028 37836 13084
rect 37772 13024 37836 13028
rect 37852 13084 37916 13088
rect 37852 13028 37856 13084
rect 37856 13028 37912 13084
rect 37912 13028 37916 13084
rect 37852 13024 37916 13028
rect 1952 12540 2016 12544
rect 1952 12484 1956 12540
rect 1956 12484 2012 12540
rect 2012 12484 2016 12540
rect 1952 12480 2016 12484
rect 2032 12540 2096 12544
rect 2032 12484 2036 12540
rect 2036 12484 2092 12540
rect 2092 12484 2096 12540
rect 2032 12480 2096 12484
rect 2112 12540 2176 12544
rect 2112 12484 2116 12540
rect 2116 12484 2172 12540
rect 2172 12484 2176 12540
rect 2112 12480 2176 12484
rect 2192 12540 2256 12544
rect 2192 12484 2196 12540
rect 2196 12484 2252 12540
rect 2252 12484 2256 12540
rect 2192 12480 2256 12484
rect 6952 12540 7016 12544
rect 6952 12484 6956 12540
rect 6956 12484 7012 12540
rect 7012 12484 7016 12540
rect 6952 12480 7016 12484
rect 7032 12540 7096 12544
rect 7032 12484 7036 12540
rect 7036 12484 7092 12540
rect 7092 12484 7096 12540
rect 7032 12480 7096 12484
rect 7112 12540 7176 12544
rect 7112 12484 7116 12540
rect 7116 12484 7172 12540
rect 7172 12484 7176 12540
rect 7112 12480 7176 12484
rect 7192 12540 7256 12544
rect 7192 12484 7196 12540
rect 7196 12484 7252 12540
rect 7252 12484 7256 12540
rect 7192 12480 7256 12484
rect 11952 12540 12016 12544
rect 11952 12484 11956 12540
rect 11956 12484 12012 12540
rect 12012 12484 12016 12540
rect 11952 12480 12016 12484
rect 12032 12540 12096 12544
rect 12032 12484 12036 12540
rect 12036 12484 12092 12540
rect 12092 12484 12096 12540
rect 12032 12480 12096 12484
rect 12112 12540 12176 12544
rect 12112 12484 12116 12540
rect 12116 12484 12172 12540
rect 12172 12484 12176 12540
rect 12112 12480 12176 12484
rect 12192 12540 12256 12544
rect 12192 12484 12196 12540
rect 12196 12484 12252 12540
rect 12252 12484 12256 12540
rect 12192 12480 12256 12484
rect 16952 12540 17016 12544
rect 16952 12484 16956 12540
rect 16956 12484 17012 12540
rect 17012 12484 17016 12540
rect 16952 12480 17016 12484
rect 17032 12540 17096 12544
rect 17032 12484 17036 12540
rect 17036 12484 17092 12540
rect 17092 12484 17096 12540
rect 17032 12480 17096 12484
rect 17112 12540 17176 12544
rect 17112 12484 17116 12540
rect 17116 12484 17172 12540
rect 17172 12484 17176 12540
rect 17112 12480 17176 12484
rect 17192 12540 17256 12544
rect 17192 12484 17196 12540
rect 17196 12484 17252 12540
rect 17252 12484 17256 12540
rect 17192 12480 17256 12484
rect 21952 12540 22016 12544
rect 21952 12484 21956 12540
rect 21956 12484 22012 12540
rect 22012 12484 22016 12540
rect 21952 12480 22016 12484
rect 22032 12540 22096 12544
rect 22032 12484 22036 12540
rect 22036 12484 22092 12540
rect 22092 12484 22096 12540
rect 22032 12480 22096 12484
rect 22112 12540 22176 12544
rect 22112 12484 22116 12540
rect 22116 12484 22172 12540
rect 22172 12484 22176 12540
rect 22112 12480 22176 12484
rect 22192 12540 22256 12544
rect 22192 12484 22196 12540
rect 22196 12484 22252 12540
rect 22252 12484 22256 12540
rect 22192 12480 22256 12484
rect 26952 12540 27016 12544
rect 26952 12484 26956 12540
rect 26956 12484 27012 12540
rect 27012 12484 27016 12540
rect 26952 12480 27016 12484
rect 27032 12540 27096 12544
rect 27032 12484 27036 12540
rect 27036 12484 27092 12540
rect 27092 12484 27096 12540
rect 27032 12480 27096 12484
rect 27112 12540 27176 12544
rect 27112 12484 27116 12540
rect 27116 12484 27172 12540
rect 27172 12484 27176 12540
rect 27112 12480 27176 12484
rect 27192 12540 27256 12544
rect 27192 12484 27196 12540
rect 27196 12484 27252 12540
rect 27252 12484 27256 12540
rect 27192 12480 27256 12484
rect 31952 12540 32016 12544
rect 31952 12484 31956 12540
rect 31956 12484 32012 12540
rect 32012 12484 32016 12540
rect 31952 12480 32016 12484
rect 32032 12540 32096 12544
rect 32032 12484 32036 12540
rect 32036 12484 32092 12540
rect 32092 12484 32096 12540
rect 32032 12480 32096 12484
rect 32112 12540 32176 12544
rect 32112 12484 32116 12540
rect 32116 12484 32172 12540
rect 32172 12484 32176 12540
rect 32112 12480 32176 12484
rect 32192 12540 32256 12544
rect 32192 12484 32196 12540
rect 32196 12484 32252 12540
rect 32252 12484 32256 12540
rect 32192 12480 32256 12484
rect 36952 12540 37016 12544
rect 36952 12484 36956 12540
rect 36956 12484 37012 12540
rect 37012 12484 37016 12540
rect 36952 12480 37016 12484
rect 37032 12540 37096 12544
rect 37032 12484 37036 12540
rect 37036 12484 37092 12540
rect 37092 12484 37096 12540
rect 37032 12480 37096 12484
rect 37112 12540 37176 12544
rect 37112 12484 37116 12540
rect 37116 12484 37172 12540
rect 37172 12484 37176 12540
rect 37112 12480 37176 12484
rect 37192 12540 37256 12544
rect 37192 12484 37196 12540
rect 37196 12484 37252 12540
rect 37252 12484 37256 12540
rect 37192 12480 37256 12484
rect 20484 12140 20548 12204
rect 2612 11996 2676 12000
rect 2612 11940 2616 11996
rect 2616 11940 2672 11996
rect 2672 11940 2676 11996
rect 2612 11936 2676 11940
rect 2692 11996 2756 12000
rect 2692 11940 2696 11996
rect 2696 11940 2752 11996
rect 2752 11940 2756 11996
rect 2692 11936 2756 11940
rect 2772 11996 2836 12000
rect 2772 11940 2776 11996
rect 2776 11940 2832 11996
rect 2832 11940 2836 11996
rect 2772 11936 2836 11940
rect 2852 11996 2916 12000
rect 2852 11940 2856 11996
rect 2856 11940 2912 11996
rect 2912 11940 2916 11996
rect 2852 11936 2916 11940
rect 7612 11996 7676 12000
rect 7612 11940 7616 11996
rect 7616 11940 7672 11996
rect 7672 11940 7676 11996
rect 7612 11936 7676 11940
rect 7692 11996 7756 12000
rect 7692 11940 7696 11996
rect 7696 11940 7752 11996
rect 7752 11940 7756 11996
rect 7692 11936 7756 11940
rect 7772 11996 7836 12000
rect 7772 11940 7776 11996
rect 7776 11940 7832 11996
rect 7832 11940 7836 11996
rect 7772 11936 7836 11940
rect 7852 11996 7916 12000
rect 7852 11940 7856 11996
rect 7856 11940 7912 11996
rect 7912 11940 7916 11996
rect 7852 11936 7916 11940
rect 12612 11996 12676 12000
rect 12612 11940 12616 11996
rect 12616 11940 12672 11996
rect 12672 11940 12676 11996
rect 12612 11936 12676 11940
rect 12692 11996 12756 12000
rect 12692 11940 12696 11996
rect 12696 11940 12752 11996
rect 12752 11940 12756 11996
rect 12692 11936 12756 11940
rect 12772 11996 12836 12000
rect 12772 11940 12776 11996
rect 12776 11940 12832 11996
rect 12832 11940 12836 11996
rect 12772 11936 12836 11940
rect 12852 11996 12916 12000
rect 12852 11940 12856 11996
rect 12856 11940 12912 11996
rect 12912 11940 12916 11996
rect 12852 11936 12916 11940
rect 17612 11996 17676 12000
rect 17612 11940 17616 11996
rect 17616 11940 17672 11996
rect 17672 11940 17676 11996
rect 17612 11936 17676 11940
rect 17692 11996 17756 12000
rect 17692 11940 17696 11996
rect 17696 11940 17752 11996
rect 17752 11940 17756 11996
rect 17692 11936 17756 11940
rect 17772 11996 17836 12000
rect 17772 11940 17776 11996
rect 17776 11940 17832 11996
rect 17832 11940 17836 11996
rect 17772 11936 17836 11940
rect 17852 11996 17916 12000
rect 17852 11940 17856 11996
rect 17856 11940 17912 11996
rect 17912 11940 17916 11996
rect 17852 11936 17916 11940
rect 22612 11996 22676 12000
rect 22612 11940 22616 11996
rect 22616 11940 22672 11996
rect 22672 11940 22676 11996
rect 22612 11936 22676 11940
rect 22692 11996 22756 12000
rect 22692 11940 22696 11996
rect 22696 11940 22752 11996
rect 22752 11940 22756 11996
rect 22692 11936 22756 11940
rect 22772 11996 22836 12000
rect 22772 11940 22776 11996
rect 22776 11940 22832 11996
rect 22832 11940 22836 11996
rect 22772 11936 22836 11940
rect 22852 11996 22916 12000
rect 22852 11940 22856 11996
rect 22856 11940 22912 11996
rect 22912 11940 22916 11996
rect 22852 11936 22916 11940
rect 27612 11996 27676 12000
rect 27612 11940 27616 11996
rect 27616 11940 27672 11996
rect 27672 11940 27676 11996
rect 27612 11936 27676 11940
rect 27692 11996 27756 12000
rect 27692 11940 27696 11996
rect 27696 11940 27752 11996
rect 27752 11940 27756 11996
rect 27692 11936 27756 11940
rect 27772 11996 27836 12000
rect 27772 11940 27776 11996
rect 27776 11940 27832 11996
rect 27832 11940 27836 11996
rect 27772 11936 27836 11940
rect 27852 11996 27916 12000
rect 27852 11940 27856 11996
rect 27856 11940 27912 11996
rect 27912 11940 27916 11996
rect 27852 11936 27916 11940
rect 32612 11996 32676 12000
rect 32612 11940 32616 11996
rect 32616 11940 32672 11996
rect 32672 11940 32676 11996
rect 32612 11936 32676 11940
rect 32692 11996 32756 12000
rect 32692 11940 32696 11996
rect 32696 11940 32752 11996
rect 32752 11940 32756 11996
rect 32692 11936 32756 11940
rect 32772 11996 32836 12000
rect 32772 11940 32776 11996
rect 32776 11940 32832 11996
rect 32832 11940 32836 11996
rect 32772 11936 32836 11940
rect 32852 11996 32916 12000
rect 32852 11940 32856 11996
rect 32856 11940 32912 11996
rect 32912 11940 32916 11996
rect 32852 11936 32916 11940
rect 37612 11996 37676 12000
rect 37612 11940 37616 11996
rect 37616 11940 37672 11996
rect 37672 11940 37676 11996
rect 37612 11936 37676 11940
rect 37692 11996 37756 12000
rect 37692 11940 37696 11996
rect 37696 11940 37752 11996
rect 37752 11940 37756 11996
rect 37692 11936 37756 11940
rect 37772 11996 37836 12000
rect 37772 11940 37776 11996
rect 37776 11940 37832 11996
rect 37832 11940 37836 11996
rect 37772 11936 37836 11940
rect 37852 11996 37916 12000
rect 37852 11940 37856 11996
rect 37856 11940 37912 11996
rect 37912 11940 37916 11996
rect 37852 11936 37916 11940
rect 34836 11596 34900 11660
rect 1952 11452 2016 11456
rect 1952 11396 1956 11452
rect 1956 11396 2012 11452
rect 2012 11396 2016 11452
rect 1952 11392 2016 11396
rect 2032 11452 2096 11456
rect 2032 11396 2036 11452
rect 2036 11396 2092 11452
rect 2092 11396 2096 11452
rect 2032 11392 2096 11396
rect 2112 11452 2176 11456
rect 2112 11396 2116 11452
rect 2116 11396 2172 11452
rect 2172 11396 2176 11452
rect 2112 11392 2176 11396
rect 2192 11452 2256 11456
rect 2192 11396 2196 11452
rect 2196 11396 2252 11452
rect 2252 11396 2256 11452
rect 2192 11392 2256 11396
rect 6952 11452 7016 11456
rect 6952 11396 6956 11452
rect 6956 11396 7012 11452
rect 7012 11396 7016 11452
rect 6952 11392 7016 11396
rect 7032 11452 7096 11456
rect 7032 11396 7036 11452
rect 7036 11396 7092 11452
rect 7092 11396 7096 11452
rect 7032 11392 7096 11396
rect 7112 11452 7176 11456
rect 7112 11396 7116 11452
rect 7116 11396 7172 11452
rect 7172 11396 7176 11452
rect 7112 11392 7176 11396
rect 7192 11452 7256 11456
rect 7192 11396 7196 11452
rect 7196 11396 7252 11452
rect 7252 11396 7256 11452
rect 7192 11392 7256 11396
rect 11952 11452 12016 11456
rect 11952 11396 11956 11452
rect 11956 11396 12012 11452
rect 12012 11396 12016 11452
rect 11952 11392 12016 11396
rect 12032 11452 12096 11456
rect 12032 11396 12036 11452
rect 12036 11396 12092 11452
rect 12092 11396 12096 11452
rect 12032 11392 12096 11396
rect 12112 11452 12176 11456
rect 12112 11396 12116 11452
rect 12116 11396 12172 11452
rect 12172 11396 12176 11452
rect 12112 11392 12176 11396
rect 12192 11452 12256 11456
rect 12192 11396 12196 11452
rect 12196 11396 12252 11452
rect 12252 11396 12256 11452
rect 12192 11392 12256 11396
rect 16952 11452 17016 11456
rect 16952 11396 16956 11452
rect 16956 11396 17012 11452
rect 17012 11396 17016 11452
rect 16952 11392 17016 11396
rect 17032 11452 17096 11456
rect 17032 11396 17036 11452
rect 17036 11396 17092 11452
rect 17092 11396 17096 11452
rect 17032 11392 17096 11396
rect 17112 11452 17176 11456
rect 17112 11396 17116 11452
rect 17116 11396 17172 11452
rect 17172 11396 17176 11452
rect 17112 11392 17176 11396
rect 17192 11452 17256 11456
rect 17192 11396 17196 11452
rect 17196 11396 17252 11452
rect 17252 11396 17256 11452
rect 17192 11392 17256 11396
rect 21952 11452 22016 11456
rect 21952 11396 21956 11452
rect 21956 11396 22012 11452
rect 22012 11396 22016 11452
rect 21952 11392 22016 11396
rect 22032 11452 22096 11456
rect 22032 11396 22036 11452
rect 22036 11396 22092 11452
rect 22092 11396 22096 11452
rect 22032 11392 22096 11396
rect 22112 11452 22176 11456
rect 22112 11396 22116 11452
rect 22116 11396 22172 11452
rect 22172 11396 22176 11452
rect 22112 11392 22176 11396
rect 22192 11452 22256 11456
rect 22192 11396 22196 11452
rect 22196 11396 22252 11452
rect 22252 11396 22256 11452
rect 22192 11392 22256 11396
rect 26952 11452 27016 11456
rect 26952 11396 26956 11452
rect 26956 11396 27012 11452
rect 27012 11396 27016 11452
rect 26952 11392 27016 11396
rect 27032 11452 27096 11456
rect 27032 11396 27036 11452
rect 27036 11396 27092 11452
rect 27092 11396 27096 11452
rect 27032 11392 27096 11396
rect 27112 11452 27176 11456
rect 27112 11396 27116 11452
rect 27116 11396 27172 11452
rect 27172 11396 27176 11452
rect 27112 11392 27176 11396
rect 27192 11452 27256 11456
rect 27192 11396 27196 11452
rect 27196 11396 27252 11452
rect 27252 11396 27256 11452
rect 27192 11392 27256 11396
rect 31952 11452 32016 11456
rect 31952 11396 31956 11452
rect 31956 11396 32012 11452
rect 32012 11396 32016 11452
rect 31952 11392 32016 11396
rect 32032 11452 32096 11456
rect 32032 11396 32036 11452
rect 32036 11396 32092 11452
rect 32092 11396 32096 11452
rect 32032 11392 32096 11396
rect 32112 11452 32176 11456
rect 32112 11396 32116 11452
rect 32116 11396 32172 11452
rect 32172 11396 32176 11452
rect 32112 11392 32176 11396
rect 32192 11452 32256 11456
rect 32192 11396 32196 11452
rect 32196 11396 32252 11452
rect 32252 11396 32256 11452
rect 32192 11392 32256 11396
rect 36952 11452 37016 11456
rect 36952 11396 36956 11452
rect 36956 11396 37012 11452
rect 37012 11396 37016 11452
rect 36952 11392 37016 11396
rect 37032 11452 37096 11456
rect 37032 11396 37036 11452
rect 37036 11396 37092 11452
rect 37092 11396 37096 11452
rect 37032 11392 37096 11396
rect 37112 11452 37176 11456
rect 37112 11396 37116 11452
rect 37116 11396 37172 11452
rect 37172 11396 37176 11452
rect 37112 11392 37176 11396
rect 37192 11452 37256 11456
rect 37192 11396 37196 11452
rect 37196 11396 37252 11452
rect 37252 11396 37256 11452
rect 37192 11392 37256 11396
rect 3372 11052 3436 11116
rect 2612 10908 2676 10912
rect 2612 10852 2616 10908
rect 2616 10852 2672 10908
rect 2672 10852 2676 10908
rect 2612 10848 2676 10852
rect 2692 10908 2756 10912
rect 2692 10852 2696 10908
rect 2696 10852 2752 10908
rect 2752 10852 2756 10908
rect 2692 10848 2756 10852
rect 2772 10908 2836 10912
rect 2772 10852 2776 10908
rect 2776 10852 2832 10908
rect 2832 10852 2836 10908
rect 2772 10848 2836 10852
rect 2852 10908 2916 10912
rect 2852 10852 2856 10908
rect 2856 10852 2912 10908
rect 2912 10852 2916 10908
rect 2852 10848 2916 10852
rect 7612 10908 7676 10912
rect 7612 10852 7616 10908
rect 7616 10852 7672 10908
rect 7672 10852 7676 10908
rect 7612 10848 7676 10852
rect 7692 10908 7756 10912
rect 7692 10852 7696 10908
rect 7696 10852 7752 10908
rect 7752 10852 7756 10908
rect 7692 10848 7756 10852
rect 7772 10908 7836 10912
rect 7772 10852 7776 10908
rect 7776 10852 7832 10908
rect 7832 10852 7836 10908
rect 7772 10848 7836 10852
rect 7852 10908 7916 10912
rect 7852 10852 7856 10908
rect 7856 10852 7912 10908
rect 7912 10852 7916 10908
rect 7852 10848 7916 10852
rect 12612 10908 12676 10912
rect 12612 10852 12616 10908
rect 12616 10852 12672 10908
rect 12672 10852 12676 10908
rect 12612 10848 12676 10852
rect 12692 10908 12756 10912
rect 12692 10852 12696 10908
rect 12696 10852 12752 10908
rect 12752 10852 12756 10908
rect 12692 10848 12756 10852
rect 12772 10908 12836 10912
rect 12772 10852 12776 10908
rect 12776 10852 12832 10908
rect 12832 10852 12836 10908
rect 12772 10848 12836 10852
rect 12852 10908 12916 10912
rect 12852 10852 12856 10908
rect 12856 10852 12912 10908
rect 12912 10852 12916 10908
rect 12852 10848 12916 10852
rect 17612 10908 17676 10912
rect 17612 10852 17616 10908
rect 17616 10852 17672 10908
rect 17672 10852 17676 10908
rect 17612 10848 17676 10852
rect 17692 10908 17756 10912
rect 17692 10852 17696 10908
rect 17696 10852 17752 10908
rect 17752 10852 17756 10908
rect 17692 10848 17756 10852
rect 17772 10908 17836 10912
rect 17772 10852 17776 10908
rect 17776 10852 17832 10908
rect 17832 10852 17836 10908
rect 17772 10848 17836 10852
rect 17852 10908 17916 10912
rect 17852 10852 17856 10908
rect 17856 10852 17912 10908
rect 17912 10852 17916 10908
rect 17852 10848 17916 10852
rect 22612 10908 22676 10912
rect 22612 10852 22616 10908
rect 22616 10852 22672 10908
rect 22672 10852 22676 10908
rect 22612 10848 22676 10852
rect 22692 10908 22756 10912
rect 22692 10852 22696 10908
rect 22696 10852 22752 10908
rect 22752 10852 22756 10908
rect 22692 10848 22756 10852
rect 22772 10908 22836 10912
rect 22772 10852 22776 10908
rect 22776 10852 22832 10908
rect 22832 10852 22836 10908
rect 22772 10848 22836 10852
rect 22852 10908 22916 10912
rect 22852 10852 22856 10908
rect 22856 10852 22912 10908
rect 22912 10852 22916 10908
rect 22852 10848 22916 10852
rect 27612 10908 27676 10912
rect 27612 10852 27616 10908
rect 27616 10852 27672 10908
rect 27672 10852 27676 10908
rect 27612 10848 27676 10852
rect 27692 10908 27756 10912
rect 27692 10852 27696 10908
rect 27696 10852 27752 10908
rect 27752 10852 27756 10908
rect 27692 10848 27756 10852
rect 27772 10908 27836 10912
rect 27772 10852 27776 10908
rect 27776 10852 27832 10908
rect 27832 10852 27836 10908
rect 27772 10848 27836 10852
rect 27852 10908 27916 10912
rect 27852 10852 27856 10908
rect 27856 10852 27912 10908
rect 27912 10852 27916 10908
rect 27852 10848 27916 10852
rect 32612 10908 32676 10912
rect 32612 10852 32616 10908
rect 32616 10852 32672 10908
rect 32672 10852 32676 10908
rect 32612 10848 32676 10852
rect 32692 10908 32756 10912
rect 32692 10852 32696 10908
rect 32696 10852 32752 10908
rect 32752 10852 32756 10908
rect 32692 10848 32756 10852
rect 32772 10908 32836 10912
rect 32772 10852 32776 10908
rect 32776 10852 32832 10908
rect 32832 10852 32836 10908
rect 32772 10848 32836 10852
rect 32852 10908 32916 10912
rect 32852 10852 32856 10908
rect 32856 10852 32912 10908
rect 32912 10852 32916 10908
rect 32852 10848 32916 10852
rect 37612 10908 37676 10912
rect 37612 10852 37616 10908
rect 37616 10852 37672 10908
rect 37672 10852 37676 10908
rect 37612 10848 37676 10852
rect 37692 10908 37756 10912
rect 37692 10852 37696 10908
rect 37696 10852 37752 10908
rect 37752 10852 37756 10908
rect 37692 10848 37756 10852
rect 37772 10908 37836 10912
rect 37772 10852 37776 10908
rect 37776 10852 37832 10908
rect 37832 10852 37836 10908
rect 37772 10848 37836 10852
rect 37852 10908 37916 10912
rect 37852 10852 37856 10908
rect 37856 10852 37912 10908
rect 37912 10852 37916 10908
rect 37852 10848 37916 10852
rect 1952 10364 2016 10368
rect 1952 10308 1956 10364
rect 1956 10308 2012 10364
rect 2012 10308 2016 10364
rect 1952 10304 2016 10308
rect 2032 10364 2096 10368
rect 2032 10308 2036 10364
rect 2036 10308 2092 10364
rect 2092 10308 2096 10364
rect 2032 10304 2096 10308
rect 2112 10364 2176 10368
rect 2112 10308 2116 10364
rect 2116 10308 2172 10364
rect 2172 10308 2176 10364
rect 2112 10304 2176 10308
rect 2192 10364 2256 10368
rect 2192 10308 2196 10364
rect 2196 10308 2252 10364
rect 2252 10308 2256 10364
rect 2192 10304 2256 10308
rect 6952 10364 7016 10368
rect 6952 10308 6956 10364
rect 6956 10308 7012 10364
rect 7012 10308 7016 10364
rect 6952 10304 7016 10308
rect 7032 10364 7096 10368
rect 7032 10308 7036 10364
rect 7036 10308 7092 10364
rect 7092 10308 7096 10364
rect 7032 10304 7096 10308
rect 7112 10364 7176 10368
rect 7112 10308 7116 10364
rect 7116 10308 7172 10364
rect 7172 10308 7176 10364
rect 7112 10304 7176 10308
rect 7192 10364 7256 10368
rect 7192 10308 7196 10364
rect 7196 10308 7252 10364
rect 7252 10308 7256 10364
rect 7192 10304 7256 10308
rect 11952 10364 12016 10368
rect 11952 10308 11956 10364
rect 11956 10308 12012 10364
rect 12012 10308 12016 10364
rect 11952 10304 12016 10308
rect 12032 10364 12096 10368
rect 12032 10308 12036 10364
rect 12036 10308 12092 10364
rect 12092 10308 12096 10364
rect 12032 10304 12096 10308
rect 12112 10364 12176 10368
rect 12112 10308 12116 10364
rect 12116 10308 12172 10364
rect 12172 10308 12176 10364
rect 12112 10304 12176 10308
rect 12192 10364 12256 10368
rect 12192 10308 12196 10364
rect 12196 10308 12252 10364
rect 12252 10308 12256 10364
rect 12192 10304 12256 10308
rect 16952 10364 17016 10368
rect 16952 10308 16956 10364
rect 16956 10308 17012 10364
rect 17012 10308 17016 10364
rect 16952 10304 17016 10308
rect 17032 10364 17096 10368
rect 17032 10308 17036 10364
rect 17036 10308 17092 10364
rect 17092 10308 17096 10364
rect 17032 10304 17096 10308
rect 17112 10364 17176 10368
rect 17112 10308 17116 10364
rect 17116 10308 17172 10364
rect 17172 10308 17176 10364
rect 17112 10304 17176 10308
rect 17192 10364 17256 10368
rect 17192 10308 17196 10364
rect 17196 10308 17252 10364
rect 17252 10308 17256 10364
rect 17192 10304 17256 10308
rect 21952 10364 22016 10368
rect 21952 10308 21956 10364
rect 21956 10308 22012 10364
rect 22012 10308 22016 10364
rect 21952 10304 22016 10308
rect 22032 10364 22096 10368
rect 22032 10308 22036 10364
rect 22036 10308 22092 10364
rect 22092 10308 22096 10364
rect 22032 10304 22096 10308
rect 22112 10364 22176 10368
rect 22112 10308 22116 10364
rect 22116 10308 22172 10364
rect 22172 10308 22176 10364
rect 22112 10304 22176 10308
rect 22192 10364 22256 10368
rect 22192 10308 22196 10364
rect 22196 10308 22252 10364
rect 22252 10308 22256 10364
rect 22192 10304 22256 10308
rect 26952 10364 27016 10368
rect 26952 10308 26956 10364
rect 26956 10308 27012 10364
rect 27012 10308 27016 10364
rect 26952 10304 27016 10308
rect 27032 10364 27096 10368
rect 27032 10308 27036 10364
rect 27036 10308 27092 10364
rect 27092 10308 27096 10364
rect 27032 10304 27096 10308
rect 27112 10364 27176 10368
rect 27112 10308 27116 10364
rect 27116 10308 27172 10364
rect 27172 10308 27176 10364
rect 27112 10304 27176 10308
rect 27192 10364 27256 10368
rect 27192 10308 27196 10364
rect 27196 10308 27252 10364
rect 27252 10308 27256 10364
rect 27192 10304 27256 10308
rect 31952 10364 32016 10368
rect 31952 10308 31956 10364
rect 31956 10308 32012 10364
rect 32012 10308 32016 10364
rect 31952 10304 32016 10308
rect 32032 10364 32096 10368
rect 32032 10308 32036 10364
rect 32036 10308 32092 10364
rect 32092 10308 32096 10364
rect 32032 10304 32096 10308
rect 32112 10364 32176 10368
rect 32112 10308 32116 10364
rect 32116 10308 32172 10364
rect 32172 10308 32176 10364
rect 32112 10304 32176 10308
rect 32192 10364 32256 10368
rect 32192 10308 32196 10364
rect 32196 10308 32252 10364
rect 32252 10308 32256 10364
rect 32192 10304 32256 10308
rect 36952 10364 37016 10368
rect 36952 10308 36956 10364
rect 36956 10308 37012 10364
rect 37012 10308 37016 10364
rect 36952 10304 37016 10308
rect 37032 10364 37096 10368
rect 37032 10308 37036 10364
rect 37036 10308 37092 10364
rect 37092 10308 37096 10364
rect 37032 10304 37096 10308
rect 37112 10364 37176 10368
rect 37112 10308 37116 10364
rect 37116 10308 37172 10364
rect 37172 10308 37176 10364
rect 37112 10304 37176 10308
rect 37192 10364 37256 10368
rect 37192 10308 37196 10364
rect 37196 10308 37252 10364
rect 37252 10308 37256 10364
rect 37192 10304 37256 10308
rect 2612 9820 2676 9824
rect 2612 9764 2616 9820
rect 2616 9764 2672 9820
rect 2672 9764 2676 9820
rect 2612 9760 2676 9764
rect 2692 9820 2756 9824
rect 2692 9764 2696 9820
rect 2696 9764 2752 9820
rect 2752 9764 2756 9820
rect 2692 9760 2756 9764
rect 2772 9820 2836 9824
rect 2772 9764 2776 9820
rect 2776 9764 2832 9820
rect 2832 9764 2836 9820
rect 2772 9760 2836 9764
rect 2852 9820 2916 9824
rect 2852 9764 2856 9820
rect 2856 9764 2912 9820
rect 2912 9764 2916 9820
rect 2852 9760 2916 9764
rect 7612 9820 7676 9824
rect 7612 9764 7616 9820
rect 7616 9764 7672 9820
rect 7672 9764 7676 9820
rect 7612 9760 7676 9764
rect 7692 9820 7756 9824
rect 7692 9764 7696 9820
rect 7696 9764 7752 9820
rect 7752 9764 7756 9820
rect 7692 9760 7756 9764
rect 7772 9820 7836 9824
rect 7772 9764 7776 9820
rect 7776 9764 7832 9820
rect 7832 9764 7836 9820
rect 7772 9760 7836 9764
rect 7852 9820 7916 9824
rect 7852 9764 7856 9820
rect 7856 9764 7912 9820
rect 7912 9764 7916 9820
rect 7852 9760 7916 9764
rect 12612 9820 12676 9824
rect 12612 9764 12616 9820
rect 12616 9764 12672 9820
rect 12672 9764 12676 9820
rect 12612 9760 12676 9764
rect 12692 9820 12756 9824
rect 12692 9764 12696 9820
rect 12696 9764 12752 9820
rect 12752 9764 12756 9820
rect 12692 9760 12756 9764
rect 12772 9820 12836 9824
rect 12772 9764 12776 9820
rect 12776 9764 12832 9820
rect 12832 9764 12836 9820
rect 12772 9760 12836 9764
rect 12852 9820 12916 9824
rect 12852 9764 12856 9820
rect 12856 9764 12912 9820
rect 12912 9764 12916 9820
rect 12852 9760 12916 9764
rect 17612 9820 17676 9824
rect 17612 9764 17616 9820
rect 17616 9764 17672 9820
rect 17672 9764 17676 9820
rect 17612 9760 17676 9764
rect 17692 9820 17756 9824
rect 17692 9764 17696 9820
rect 17696 9764 17752 9820
rect 17752 9764 17756 9820
rect 17692 9760 17756 9764
rect 17772 9820 17836 9824
rect 17772 9764 17776 9820
rect 17776 9764 17832 9820
rect 17832 9764 17836 9820
rect 17772 9760 17836 9764
rect 17852 9820 17916 9824
rect 17852 9764 17856 9820
rect 17856 9764 17912 9820
rect 17912 9764 17916 9820
rect 17852 9760 17916 9764
rect 22612 9820 22676 9824
rect 22612 9764 22616 9820
rect 22616 9764 22672 9820
rect 22672 9764 22676 9820
rect 22612 9760 22676 9764
rect 22692 9820 22756 9824
rect 22692 9764 22696 9820
rect 22696 9764 22752 9820
rect 22752 9764 22756 9820
rect 22692 9760 22756 9764
rect 22772 9820 22836 9824
rect 22772 9764 22776 9820
rect 22776 9764 22832 9820
rect 22832 9764 22836 9820
rect 22772 9760 22836 9764
rect 22852 9820 22916 9824
rect 22852 9764 22856 9820
rect 22856 9764 22912 9820
rect 22912 9764 22916 9820
rect 22852 9760 22916 9764
rect 27612 9820 27676 9824
rect 27612 9764 27616 9820
rect 27616 9764 27672 9820
rect 27672 9764 27676 9820
rect 27612 9760 27676 9764
rect 27692 9820 27756 9824
rect 27692 9764 27696 9820
rect 27696 9764 27752 9820
rect 27752 9764 27756 9820
rect 27692 9760 27756 9764
rect 27772 9820 27836 9824
rect 27772 9764 27776 9820
rect 27776 9764 27832 9820
rect 27832 9764 27836 9820
rect 27772 9760 27836 9764
rect 27852 9820 27916 9824
rect 27852 9764 27856 9820
rect 27856 9764 27912 9820
rect 27912 9764 27916 9820
rect 27852 9760 27916 9764
rect 32612 9820 32676 9824
rect 32612 9764 32616 9820
rect 32616 9764 32672 9820
rect 32672 9764 32676 9820
rect 32612 9760 32676 9764
rect 32692 9820 32756 9824
rect 32692 9764 32696 9820
rect 32696 9764 32752 9820
rect 32752 9764 32756 9820
rect 32692 9760 32756 9764
rect 32772 9820 32836 9824
rect 32772 9764 32776 9820
rect 32776 9764 32832 9820
rect 32832 9764 32836 9820
rect 32772 9760 32836 9764
rect 32852 9820 32916 9824
rect 32852 9764 32856 9820
rect 32856 9764 32912 9820
rect 32912 9764 32916 9820
rect 32852 9760 32916 9764
rect 37612 9820 37676 9824
rect 37612 9764 37616 9820
rect 37616 9764 37672 9820
rect 37672 9764 37676 9820
rect 37612 9760 37676 9764
rect 37692 9820 37756 9824
rect 37692 9764 37696 9820
rect 37696 9764 37752 9820
rect 37752 9764 37756 9820
rect 37692 9760 37756 9764
rect 37772 9820 37836 9824
rect 37772 9764 37776 9820
rect 37776 9764 37832 9820
rect 37832 9764 37836 9820
rect 37772 9760 37836 9764
rect 37852 9820 37916 9824
rect 37852 9764 37856 9820
rect 37856 9764 37912 9820
rect 37912 9764 37916 9820
rect 37852 9760 37916 9764
rect 1952 9276 2016 9280
rect 1952 9220 1956 9276
rect 1956 9220 2012 9276
rect 2012 9220 2016 9276
rect 1952 9216 2016 9220
rect 2032 9276 2096 9280
rect 2032 9220 2036 9276
rect 2036 9220 2092 9276
rect 2092 9220 2096 9276
rect 2032 9216 2096 9220
rect 2112 9276 2176 9280
rect 2112 9220 2116 9276
rect 2116 9220 2172 9276
rect 2172 9220 2176 9276
rect 2112 9216 2176 9220
rect 2192 9276 2256 9280
rect 2192 9220 2196 9276
rect 2196 9220 2252 9276
rect 2252 9220 2256 9276
rect 2192 9216 2256 9220
rect 6952 9276 7016 9280
rect 6952 9220 6956 9276
rect 6956 9220 7012 9276
rect 7012 9220 7016 9276
rect 6952 9216 7016 9220
rect 7032 9276 7096 9280
rect 7032 9220 7036 9276
rect 7036 9220 7092 9276
rect 7092 9220 7096 9276
rect 7032 9216 7096 9220
rect 7112 9276 7176 9280
rect 7112 9220 7116 9276
rect 7116 9220 7172 9276
rect 7172 9220 7176 9276
rect 7112 9216 7176 9220
rect 7192 9276 7256 9280
rect 7192 9220 7196 9276
rect 7196 9220 7252 9276
rect 7252 9220 7256 9276
rect 7192 9216 7256 9220
rect 11952 9276 12016 9280
rect 11952 9220 11956 9276
rect 11956 9220 12012 9276
rect 12012 9220 12016 9276
rect 11952 9216 12016 9220
rect 12032 9276 12096 9280
rect 12032 9220 12036 9276
rect 12036 9220 12092 9276
rect 12092 9220 12096 9276
rect 12032 9216 12096 9220
rect 12112 9276 12176 9280
rect 12112 9220 12116 9276
rect 12116 9220 12172 9276
rect 12172 9220 12176 9276
rect 12112 9216 12176 9220
rect 12192 9276 12256 9280
rect 12192 9220 12196 9276
rect 12196 9220 12252 9276
rect 12252 9220 12256 9276
rect 12192 9216 12256 9220
rect 16952 9276 17016 9280
rect 16952 9220 16956 9276
rect 16956 9220 17012 9276
rect 17012 9220 17016 9276
rect 16952 9216 17016 9220
rect 17032 9276 17096 9280
rect 17032 9220 17036 9276
rect 17036 9220 17092 9276
rect 17092 9220 17096 9276
rect 17032 9216 17096 9220
rect 17112 9276 17176 9280
rect 17112 9220 17116 9276
rect 17116 9220 17172 9276
rect 17172 9220 17176 9276
rect 17112 9216 17176 9220
rect 17192 9276 17256 9280
rect 17192 9220 17196 9276
rect 17196 9220 17252 9276
rect 17252 9220 17256 9276
rect 17192 9216 17256 9220
rect 21952 9276 22016 9280
rect 21952 9220 21956 9276
rect 21956 9220 22012 9276
rect 22012 9220 22016 9276
rect 21952 9216 22016 9220
rect 22032 9276 22096 9280
rect 22032 9220 22036 9276
rect 22036 9220 22092 9276
rect 22092 9220 22096 9276
rect 22032 9216 22096 9220
rect 22112 9276 22176 9280
rect 22112 9220 22116 9276
rect 22116 9220 22172 9276
rect 22172 9220 22176 9276
rect 22112 9216 22176 9220
rect 22192 9276 22256 9280
rect 22192 9220 22196 9276
rect 22196 9220 22252 9276
rect 22252 9220 22256 9276
rect 22192 9216 22256 9220
rect 26952 9276 27016 9280
rect 26952 9220 26956 9276
rect 26956 9220 27012 9276
rect 27012 9220 27016 9276
rect 26952 9216 27016 9220
rect 27032 9276 27096 9280
rect 27032 9220 27036 9276
rect 27036 9220 27092 9276
rect 27092 9220 27096 9276
rect 27032 9216 27096 9220
rect 27112 9276 27176 9280
rect 27112 9220 27116 9276
rect 27116 9220 27172 9276
rect 27172 9220 27176 9276
rect 27112 9216 27176 9220
rect 27192 9276 27256 9280
rect 27192 9220 27196 9276
rect 27196 9220 27252 9276
rect 27252 9220 27256 9276
rect 27192 9216 27256 9220
rect 31952 9276 32016 9280
rect 31952 9220 31956 9276
rect 31956 9220 32012 9276
rect 32012 9220 32016 9276
rect 31952 9216 32016 9220
rect 32032 9276 32096 9280
rect 32032 9220 32036 9276
rect 32036 9220 32092 9276
rect 32092 9220 32096 9276
rect 32032 9216 32096 9220
rect 32112 9276 32176 9280
rect 32112 9220 32116 9276
rect 32116 9220 32172 9276
rect 32172 9220 32176 9276
rect 32112 9216 32176 9220
rect 32192 9276 32256 9280
rect 32192 9220 32196 9276
rect 32196 9220 32252 9276
rect 32252 9220 32256 9276
rect 32192 9216 32256 9220
rect 36952 9276 37016 9280
rect 36952 9220 36956 9276
rect 36956 9220 37012 9276
rect 37012 9220 37016 9276
rect 36952 9216 37016 9220
rect 37032 9276 37096 9280
rect 37032 9220 37036 9276
rect 37036 9220 37092 9276
rect 37092 9220 37096 9276
rect 37032 9216 37096 9220
rect 37112 9276 37176 9280
rect 37112 9220 37116 9276
rect 37116 9220 37172 9276
rect 37172 9220 37176 9276
rect 37112 9216 37176 9220
rect 37192 9276 37256 9280
rect 37192 9220 37196 9276
rect 37196 9220 37252 9276
rect 37252 9220 37256 9276
rect 37192 9216 37256 9220
rect 2612 8732 2676 8736
rect 2612 8676 2616 8732
rect 2616 8676 2672 8732
rect 2672 8676 2676 8732
rect 2612 8672 2676 8676
rect 2692 8732 2756 8736
rect 2692 8676 2696 8732
rect 2696 8676 2752 8732
rect 2752 8676 2756 8732
rect 2692 8672 2756 8676
rect 2772 8732 2836 8736
rect 2772 8676 2776 8732
rect 2776 8676 2832 8732
rect 2832 8676 2836 8732
rect 2772 8672 2836 8676
rect 2852 8732 2916 8736
rect 2852 8676 2856 8732
rect 2856 8676 2912 8732
rect 2912 8676 2916 8732
rect 2852 8672 2916 8676
rect 7612 8732 7676 8736
rect 7612 8676 7616 8732
rect 7616 8676 7672 8732
rect 7672 8676 7676 8732
rect 7612 8672 7676 8676
rect 7692 8732 7756 8736
rect 7692 8676 7696 8732
rect 7696 8676 7752 8732
rect 7752 8676 7756 8732
rect 7692 8672 7756 8676
rect 7772 8732 7836 8736
rect 7772 8676 7776 8732
rect 7776 8676 7832 8732
rect 7832 8676 7836 8732
rect 7772 8672 7836 8676
rect 7852 8732 7916 8736
rect 7852 8676 7856 8732
rect 7856 8676 7912 8732
rect 7912 8676 7916 8732
rect 7852 8672 7916 8676
rect 12612 8732 12676 8736
rect 12612 8676 12616 8732
rect 12616 8676 12672 8732
rect 12672 8676 12676 8732
rect 12612 8672 12676 8676
rect 12692 8732 12756 8736
rect 12692 8676 12696 8732
rect 12696 8676 12752 8732
rect 12752 8676 12756 8732
rect 12692 8672 12756 8676
rect 12772 8732 12836 8736
rect 12772 8676 12776 8732
rect 12776 8676 12832 8732
rect 12832 8676 12836 8732
rect 12772 8672 12836 8676
rect 12852 8732 12916 8736
rect 12852 8676 12856 8732
rect 12856 8676 12912 8732
rect 12912 8676 12916 8732
rect 12852 8672 12916 8676
rect 17612 8732 17676 8736
rect 17612 8676 17616 8732
rect 17616 8676 17672 8732
rect 17672 8676 17676 8732
rect 17612 8672 17676 8676
rect 17692 8732 17756 8736
rect 17692 8676 17696 8732
rect 17696 8676 17752 8732
rect 17752 8676 17756 8732
rect 17692 8672 17756 8676
rect 17772 8732 17836 8736
rect 17772 8676 17776 8732
rect 17776 8676 17832 8732
rect 17832 8676 17836 8732
rect 17772 8672 17836 8676
rect 17852 8732 17916 8736
rect 17852 8676 17856 8732
rect 17856 8676 17912 8732
rect 17912 8676 17916 8732
rect 17852 8672 17916 8676
rect 22612 8732 22676 8736
rect 22612 8676 22616 8732
rect 22616 8676 22672 8732
rect 22672 8676 22676 8732
rect 22612 8672 22676 8676
rect 22692 8732 22756 8736
rect 22692 8676 22696 8732
rect 22696 8676 22752 8732
rect 22752 8676 22756 8732
rect 22692 8672 22756 8676
rect 22772 8732 22836 8736
rect 22772 8676 22776 8732
rect 22776 8676 22832 8732
rect 22832 8676 22836 8732
rect 22772 8672 22836 8676
rect 22852 8732 22916 8736
rect 22852 8676 22856 8732
rect 22856 8676 22912 8732
rect 22912 8676 22916 8732
rect 22852 8672 22916 8676
rect 27612 8732 27676 8736
rect 27612 8676 27616 8732
rect 27616 8676 27672 8732
rect 27672 8676 27676 8732
rect 27612 8672 27676 8676
rect 27692 8732 27756 8736
rect 27692 8676 27696 8732
rect 27696 8676 27752 8732
rect 27752 8676 27756 8732
rect 27692 8672 27756 8676
rect 27772 8732 27836 8736
rect 27772 8676 27776 8732
rect 27776 8676 27832 8732
rect 27832 8676 27836 8732
rect 27772 8672 27836 8676
rect 27852 8732 27916 8736
rect 27852 8676 27856 8732
rect 27856 8676 27912 8732
rect 27912 8676 27916 8732
rect 27852 8672 27916 8676
rect 32612 8732 32676 8736
rect 32612 8676 32616 8732
rect 32616 8676 32672 8732
rect 32672 8676 32676 8732
rect 32612 8672 32676 8676
rect 32692 8732 32756 8736
rect 32692 8676 32696 8732
rect 32696 8676 32752 8732
rect 32752 8676 32756 8732
rect 32692 8672 32756 8676
rect 32772 8732 32836 8736
rect 32772 8676 32776 8732
rect 32776 8676 32832 8732
rect 32832 8676 32836 8732
rect 32772 8672 32836 8676
rect 32852 8732 32916 8736
rect 32852 8676 32856 8732
rect 32856 8676 32912 8732
rect 32912 8676 32916 8732
rect 32852 8672 32916 8676
rect 37612 8732 37676 8736
rect 37612 8676 37616 8732
rect 37616 8676 37672 8732
rect 37672 8676 37676 8732
rect 37612 8672 37676 8676
rect 37692 8732 37756 8736
rect 37692 8676 37696 8732
rect 37696 8676 37752 8732
rect 37752 8676 37756 8732
rect 37692 8672 37756 8676
rect 37772 8732 37836 8736
rect 37772 8676 37776 8732
rect 37776 8676 37832 8732
rect 37832 8676 37836 8732
rect 37772 8672 37836 8676
rect 37852 8732 37916 8736
rect 37852 8676 37856 8732
rect 37856 8676 37912 8732
rect 37912 8676 37916 8732
rect 37852 8672 37916 8676
rect 1952 8188 2016 8192
rect 1952 8132 1956 8188
rect 1956 8132 2012 8188
rect 2012 8132 2016 8188
rect 1952 8128 2016 8132
rect 2032 8188 2096 8192
rect 2032 8132 2036 8188
rect 2036 8132 2092 8188
rect 2092 8132 2096 8188
rect 2032 8128 2096 8132
rect 2112 8188 2176 8192
rect 2112 8132 2116 8188
rect 2116 8132 2172 8188
rect 2172 8132 2176 8188
rect 2112 8128 2176 8132
rect 2192 8188 2256 8192
rect 2192 8132 2196 8188
rect 2196 8132 2252 8188
rect 2252 8132 2256 8188
rect 2192 8128 2256 8132
rect 6952 8188 7016 8192
rect 6952 8132 6956 8188
rect 6956 8132 7012 8188
rect 7012 8132 7016 8188
rect 6952 8128 7016 8132
rect 7032 8188 7096 8192
rect 7032 8132 7036 8188
rect 7036 8132 7092 8188
rect 7092 8132 7096 8188
rect 7032 8128 7096 8132
rect 7112 8188 7176 8192
rect 7112 8132 7116 8188
rect 7116 8132 7172 8188
rect 7172 8132 7176 8188
rect 7112 8128 7176 8132
rect 7192 8188 7256 8192
rect 7192 8132 7196 8188
rect 7196 8132 7252 8188
rect 7252 8132 7256 8188
rect 7192 8128 7256 8132
rect 11952 8188 12016 8192
rect 11952 8132 11956 8188
rect 11956 8132 12012 8188
rect 12012 8132 12016 8188
rect 11952 8128 12016 8132
rect 12032 8188 12096 8192
rect 12032 8132 12036 8188
rect 12036 8132 12092 8188
rect 12092 8132 12096 8188
rect 12032 8128 12096 8132
rect 12112 8188 12176 8192
rect 12112 8132 12116 8188
rect 12116 8132 12172 8188
rect 12172 8132 12176 8188
rect 12112 8128 12176 8132
rect 12192 8188 12256 8192
rect 12192 8132 12196 8188
rect 12196 8132 12252 8188
rect 12252 8132 12256 8188
rect 12192 8128 12256 8132
rect 16952 8188 17016 8192
rect 16952 8132 16956 8188
rect 16956 8132 17012 8188
rect 17012 8132 17016 8188
rect 16952 8128 17016 8132
rect 17032 8188 17096 8192
rect 17032 8132 17036 8188
rect 17036 8132 17092 8188
rect 17092 8132 17096 8188
rect 17032 8128 17096 8132
rect 17112 8188 17176 8192
rect 17112 8132 17116 8188
rect 17116 8132 17172 8188
rect 17172 8132 17176 8188
rect 17112 8128 17176 8132
rect 17192 8188 17256 8192
rect 17192 8132 17196 8188
rect 17196 8132 17252 8188
rect 17252 8132 17256 8188
rect 17192 8128 17256 8132
rect 21952 8188 22016 8192
rect 21952 8132 21956 8188
rect 21956 8132 22012 8188
rect 22012 8132 22016 8188
rect 21952 8128 22016 8132
rect 22032 8188 22096 8192
rect 22032 8132 22036 8188
rect 22036 8132 22092 8188
rect 22092 8132 22096 8188
rect 22032 8128 22096 8132
rect 22112 8188 22176 8192
rect 22112 8132 22116 8188
rect 22116 8132 22172 8188
rect 22172 8132 22176 8188
rect 22112 8128 22176 8132
rect 22192 8188 22256 8192
rect 22192 8132 22196 8188
rect 22196 8132 22252 8188
rect 22252 8132 22256 8188
rect 22192 8128 22256 8132
rect 26952 8188 27016 8192
rect 26952 8132 26956 8188
rect 26956 8132 27012 8188
rect 27012 8132 27016 8188
rect 26952 8128 27016 8132
rect 27032 8188 27096 8192
rect 27032 8132 27036 8188
rect 27036 8132 27092 8188
rect 27092 8132 27096 8188
rect 27032 8128 27096 8132
rect 27112 8188 27176 8192
rect 27112 8132 27116 8188
rect 27116 8132 27172 8188
rect 27172 8132 27176 8188
rect 27112 8128 27176 8132
rect 27192 8188 27256 8192
rect 27192 8132 27196 8188
rect 27196 8132 27252 8188
rect 27252 8132 27256 8188
rect 27192 8128 27256 8132
rect 31952 8188 32016 8192
rect 31952 8132 31956 8188
rect 31956 8132 32012 8188
rect 32012 8132 32016 8188
rect 31952 8128 32016 8132
rect 32032 8188 32096 8192
rect 32032 8132 32036 8188
rect 32036 8132 32092 8188
rect 32092 8132 32096 8188
rect 32032 8128 32096 8132
rect 32112 8188 32176 8192
rect 32112 8132 32116 8188
rect 32116 8132 32172 8188
rect 32172 8132 32176 8188
rect 32112 8128 32176 8132
rect 32192 8188 32256 8192
rect 32192 8132 32196 8188
rect 32196 8132 32252 8188
rect 32252 8132 32256 8188
rect 32192 8128 32256 8132
rect 36952 8188 37016 8192
rect 36952 8132 36956 8188
rect 36956 8132 37012 8188
rect 37012 8132 37016 8188
rect 36952 8128 37016 8132
rect 37032 8188 37096 8192
rect 37032 8132 37036 8188
rect 37036 8132 37092 8188
rect 37092 8132 37096 8188
rect 37032 8128 37096 8132
rect 37112 8188 37176 8192
rect 37112 8132 37116 8188
rect 37116 8132 37172 8188
rect 37172 8132 37176 8188
rect 37112 8128 37176 8132
rect 37192 8188 37256 8192
rect 37192 8132 37196 8188
rect 37196 8132 37252 8188
rect 37252 8132 37256 8188
rect 37192 8128 37256 8132
rect 2612 7644 2676 7648
rect 2612 7588 2616 7644
rect 2616 7588 2672 7644
rect 2672 7588 2676 7644
rect 2612 7584 2676 7588
rect 2692 7644 2756 7648
rect 2692 7588 2696 7644
rect 2696 7588 2752 7644
rect 2752 7588 2756 7644
rect 2692 7584 2756 7588
rect 2772 7644 2836 7648
rect 2772 7588 2776 7644
rect 2776 7588 2832 7644
rect 2832 7588 2836 7644
rect 2772 7584 2836 7588
rect 2852 7644 2916 7648
rect 2852 7588 2856 7644
rect 2856 7588 2912 7644
rect 2912 7588 2916 7644
rect 2852 7584 2916 7588
rect 7612 7644 7676 7648
rect 7612 7588 7616 7644
rect 7616 7588 7672 7644
rect 7672 7588 7676 7644
rect 7612 7584 7676 7588
rect 7692 7644 7756 7648
rect 7692 7588 7696 7644
rect 7696 7588 7752 7644
rect 7752 7588 7756 7644
rect 7692 7584 7756 7588
rect 7772 7644 7836 7648
rect 7772 7588 7776 7644
rect 7776 7588 7832 7644
rect 7832 7588 7836 7644
rect 7772 7584 7836 7588
rect 7852 7644 7916 7648
rect 7852 7588 7856 7644
rect 7856 7588 7912 7644
rect 7912 7588 7916 7644
rect 7852 7584 7916 7588
rect 12612 7644 12676 7648
rect 12612 7588 12616 7644
rect 12616 7588 12672 7644
rect 12672 7588 12676 7644
rect 12612 7584 12676 7588
rect 12692 7644 12756 7648
rect 12692 7588 12696 7644
rect 12696 7588 12752 7644
rect 12752 7588 12756 7644
rect 12692 7584 12756 7588
rect 12772 7644 12836 7648
rect 12772 7588 12776 7644
rect 12776 7588 12832 7644
rect 12832 7588 12836 7644
rect 12772 7584 12836 7588
rect 12852 7644 12916 7648
rect 12852 7588 12856 7644
rect 12856 7588 12912 7644
rect 12912 7588 12916 7644
rect 12852 7584 12916 7588
rect 17612 7644 17676 7648
rect 17612 7588 17616 7644
rect 17616 7588 17672 7644
rect 17672 7588 17676 7644
rect 17612 7584 17676 7588
rect 17692 7644 17756 7648
rect 17692 7588 17696 7644
rect 17696 7588 17752 7644
rect 17752 7588 17756 7644
rect 17692 7584 17756 7588
rect 17772 7644 17836 7648
rect 17772 7588 17776 7644
rect 17776 7588 17832 7644
rect 17832 7588 17836 7644
rect 17772 7584 17836 7588
rect 17852 7644 17916 7648
rect 17852 7588 17856 7644
rect 17856 7588 17912 7644
rect 17912 7588 17916 7644
rect 17852 7584 17916 7588
rect 22612 7644 22676 7648
rect 22612 7588 22616 7644
rect 22616 7588 22672 7644
rect 22672 7588 22676 7644
rect 22612 7584 22676 7588
rect 22692 7644 22756 7648
rect 22692 7588 22696 7644
rect 22696 7588 22752 7644
rect 22752 7588 22756 7644
rect 22692 7584 22756 7588
rect 22772 7644 22836 7648
rect 22772 7588 22776 7644
rect 22776 7588 22832 7644
rect 22832 7588 22836 7644
rect 22772 7584 22836 7588
rect 22852 7644 22916 7648
rect 22852 7588 22856 7644
rect 22856 7588 22912 7644
rect 22912 7588 22916 7644
rect 22852 7584 22916 7588
rect 27612 7644 27676 7648
rect 27612 7588 27616 7644
rect 27616 7588 27672 7644
rect 27672 7588 27676 7644
rect 27612 7584 27676 7588
rect 27692 7644 27756 7648
rect 27692 7588 27696 7644
rect 27696 7588 27752 7644
rect 27752 7588 27756 7644
rect 27692 7584 27756 7588
rect 27772 7644 27836 7648
rect 27772 7588 27776 7644
rect 27776 7588 27832 7644
rect 27832 7588 27836 7644
rect 27772 7584 27836 7588
rect 27852 7644 27916 7648
rect 27852 7588 27856 7644
rect 27856 7588 27912 7644
rect 27912 7588 27916 7644
rect 27852 7584 27916 7588
rect 32612 7644 32676 7648
rect 32612 7588 32616 7644
rect 32616 7588 32672 7644
rect 32672 7588 32676 7644
rect 32612 7584 32676 7588
rect 32692 7644 32756 7648
rect 32692 7588 32696 7644
rect 32696 7588 32752 7644
rect 32752 7588 32756 7644
rect 32692 7584 32756 7588
rect 32772 7644 32836 7648
rect 32772 7588 32776 7644
rect 32776 7588 32832 7644
rect 32832 7588 32836 7644
rect 32772 7584 32836 7588
rect 32852 7644 32916 7648
rect 32852 7588 32856 7644
rect 32856 7588 32912 7644
rect 32912 7588 32916 7644
rect 32852 7584 32916 7588
rect 37612 7644 37676 7648
rect 37612 7588 37616 7644
rect 37616 7588 37672 7644
rect 37672 7588 37676 7644
rect 37612 7584 37676 7588
rect 37692 7644 37756 7648
rect 37692 7588 37696 7644
rect 37696 7588 37752 7644
rect 37752 7588 37756 7644
rect 37692 7584 37756 7588
rect 37772 7644 37836 7648
rect 37772 7588 37776 7644
rect 37776 7588 37832 7644
rect 37832 7588 37836 7644
rect 37772 7584 37836 7588
rect 37852 7644 37916 7648
rect 37852 7588 37856 7644
rect 37856 7588 37912 7644
rect 37912 7588 37916 7644
rect 37852 7584 37916 7588
rect 1952 7100 2016 7104
rect 1952 7044 1956 7100
rect 1956 7044 2012 7100
rect 2012 7044 2016 7100
rect 1952 7040 2016 7044
rect 2032 7100 2096 7104
rect 2032 7044 2036 7100
rect 2036 7044 2092 7100
rect 2092 7044 2096 7100
rect 2032 7040 2096 7044
rect 2112 7100 2176 7104
rect 2112 7044 2116 7100
rect 2116 7044 2172 7100
rect 2172 7044 2176 7100
rect 2112 7040 2176 7044
rect 2192 7100 2256 7104
rect 2192 7044 2196 7100
rect 2196 7044 2252 7100
rect 2252 7044 2256 7100
rect 2192 7040 2256 7044
rect 6952 7100 7016 7104
rect 6952 7044 6956 7100
rect 6956 7044 7012 7100
rect 7012 7044 7016 7100
rect 6952 7040 7016 7044
rect 7032 7100 7096 7104
rect 7032 7044 7036 7100
rect 7036 7044 7092 7100
rect 7092 7044 7096 7100
rect 7032 7040 7096 7044
rect 7112 7100 7176 7104
rect 7112 7044 7116 7100
rect 7116 7044 7172 7100
rect 7172 7044 7176 7100
rect 7112 7040 7176 7044
rect 7192 7100 7256 7104
rect 7192 7044 7196 7100
rect 7196 7044 7252 7100
rect 7252 7044 7256 7100
rect 7192 7040 7256 7044
rect 11952 7100 12016 7104
rect 11952 7044 11956 7100
rect 11956 7044 12012 7100
rect 12012 7044 12016 7100
rect 11952 7040 12016 7044
rect 12032 7100 12096 7104
rect 12032 7044 12036 7100
rect 12036 7044 12092 7100
rect 12092 7044 12096 7100
rect 12032 7040 12096 7044
rect 12112 7100 12176 7104
rect 12112 7044 12116 7100
rect 12116 7044 12172 7100
rect 12172 7044 12176 7100
rect 12112 7040 12176 7044
rect 12192 7100 12256 7104
rect 12192 7044 12196 7100
rect 12196 7044 12252 7100
rect 12252 7044 12256 7100
rect 12192 7040 12256 7044
rect 16952 7100 17016 7104
rect 16952 7044 16956 7100
rect 16956 7044 17012 7100
rect 17012 7044 17016 7100
rect 16952 7040 17016 7044
rect 17032 7100 17096 7104
rect 17032 7044 17036 7100
rect 17036 7044 17092 7100
rect 17092 7044 17096 7100
rect 17032 7040 17096 7044
rect 17112 7100 17176 7104
rect 17112 7044 17116 7100
rect 17116 7044 17172 7100
rect 17172 7044 17176 7100
rect 17112 7040 17176 7044
rect 17192 7100 17256 7104
rect 17192 7044 17196 7100
rect 17196 7044 17252 7100
rect 17252 7044 17256 7100
rect 17192 7040 17256 7044
rect 21952 7100 22016 7104
rect 21952 7044 21956 7100
rect 21956 7044 22012 7100
rect 22012 7044 22016 7100
rect 21952 7040 22016 7044
rect 22032 7100 22096 7104
rect 22032 7044 22036 7100
rect 22036 7044 22092 7100
rect 22092 7044 22096 7100
rect 22032 7040 22096 7044
rect 22112 7100 22176 7104
rect 22112 7044 22116 7100
rect 22116 7044 22172 7100
rect 22172 7044 22176 7100
rect 22112 7040 22176 7044
rect 22192 7100 22256 7104
rect 22192 7044 22196 7100
rect 22196 7044 22252 7100
rect 22252 7044 22256 7100
rect 22192 7040 22256 7044
rect 26952 7100 27016 7104
rect 26952 7044 26956 7100
rect 26956 7044 27012 7100
rect 27012 7044 27016 7100
rect 26952 7040 27016 7044
rect 27032 7100 27096 7104
rect 27032 7044 27036 7100
rect 27036 7044 27092 7100
rect 27092 7044 27096 7100
rect 27032 7040 27096 7044
rect 27112 7100 27176 7104
rect 27112 7044 27116 7100
rect 27116 7044 27172 7100
rect 27172 7044 27176 7100
rect 27112 7040 27176 7044
rect 27192 7100 27256 7104
rect 27192 7044 27196 7100
rect 27196 7044 27252 7100
rect 27252 7044 27256 7100
rect 27192 7040 27256 7044
rect 31952 7100 32016 7104
rect 31952 7044 31956 7100
rect 31956 7044 32012 7100
rect 32012 7044 32016 7100
rect 31952 7040 32016 7044
rect 32032 7100 32096 7104
rect 32032 7044 32036 7100
rect 32036 7044 32092 7100
rect 32092 7044 32096 7100
rect 32032 7040 32096 7044
rect 32112 7100 32176 7104
rect 32112 7044 32116 7100
rect 32116 7044 32172 7100
rect 32172 7044 32176 7100
rect 32112 7040 32176 7044
rect 32192 7100 32256 7104
rect 32192 7044 32196 7100
rect 32196 7044 32252 7100
rect 32252 7044 32256 7100
rect 32192 7040 32256 7044
rect 36952 7100 37016 7104
rect 36952 7044 36956 7100
rect 36956 7044 37012 7100
rect 37012 7044 37016 7100
rect 36952 7040 37016 7044
rect 37032 7100 37096 7104
rect 37032 7044 37036 7100
rect 37036 7044 37092 7100
rect 37092 7044 37096 7100
rect 37032 7040 37096 7044
rect 37112 7100 37176 7104
rect 37112 7044 37116 7100
rect 37116 7044 37172 7100
rect 37172 7044 37176 7100
rect 37112 7040 37176 7044
rect 37192 7100 37256 7104
rect 37192 7044 37196 7100
rect 37196 7044 37252 7100
rect 37252 7044 37256 7100
rect 37192 7040 37256 7044
rect 2612 6556 2676 6560
rect 2612 6500 2616 6556
rect 2616 6500 2672 6556
rect 2672 6500 2676 6556
rect 2612 6496 2676 6500
rect 2692 6556 2756 6560
rect 2692 6500 2696 6556
rect 2696 6500 2752 6556
rect 2752 6500 2756 6556
rect 2692 6496 2756 6500
rect 2772 6556 2836 6560
rect 2772 6500 2776 6556
rect 2776 6500 2832 6556
rect 2832 6500 2836 6556
rect 2772 6496 2836 6500
rect 2852 6556 2916 6560
rect 2852 6500 2856 6556
rect 2856 6500 2912 6556
rect 2912 6500 2916 6556
rect 2852 6496 2916 6500
rect 7612 6556 7676 6560
rect 7612 6500 7616 6556
rect 7616 6500 7672 6556
rect 7672 6500 7676 6556
rect 7612 6496 7676 6500
rect 7692 6556 7756 6560
rect 7692 6500 7696 6556
rect 7696 6500 7752 6556
rect 7752 6500 7756 6556
rect 7692 6496 7756 6500
rect 7772 6556 7836 6560
rect 7772 6500 7776 6556
rect 7776 6500 7832 6556
rect 7832 6500 7836 6556
rect 7772 6496 7836 6500
rect 7852 6556 7916 6560
rect 7852 6500 7856 6556
rect 7856 6500 7912 6556
rect 7912 6500 7916 6556
rect 7852 6496 7916 6500
rect 12612 6556 12676 6560
rect 12612 6500 12616 6556
rect 12616 6500 12672 6556
rect 12672 6500 12676 6556
rect 12612 6496 12676 6500
rect 12692 6556 12756 6560
rect 12692 6500 12696 6556
rect 12696 6500 12752 6556
rect 12752 6500 12756 6556
rect 12692 6496 12756 6500
rect 12772 6556 12836 6560
rect 12772 6500 12776 6556
rect 12776 6500 12832 6556
rect 12832 6500 12836 6556
rect 12772 6496 12836 6500
rect 12852 6556 12916 6560
rect 12852 6500 12856 6556
rect 12856 6500 12912 6556
rect 12912 6500 12916 6556
rect 12852 6496 12916 6500
rect 17612 6556 17676 6560
rect 17612 6500 17616 6556
rect 17616 6500 17672 6556
rect 17672 6500 17676 6556
rect 17612 6496 17676 6500
rect 17692 6556 17756 6560
rect 17692 6500 17696 6556
rect 17696 6500 17752 6556
rect 17752 6500 17756 6556
rect 17692 6496 17756 6500
rect 17772 6556 17836 6560
rect 17772 6500 17776 6556
rect 17776 6500 17832 6556
rect 17832 6500 17836 6556
rect 17772 6496 17836 6500
rect 17852 6556 17916 6560
rect 17852 6500 17856 6556
rect 17856 6500 17912 6556
rect 17912 6500 17916 6556
rect 17852 6496 17916 6500
rect 22612 6556 22676 6560
rect 22612 6500 22616 6556
rect 22616 6500 22672 6556
rect 22672 6500 22676 6556
rect 22612 6496 22676 6500
rect 22692 6556 22756 6560
rect 22692 6500 22696 6556
rect 22696 6500 22752 6556
rect 22752 6500 22756 6556
rect 22692 6496 22756 6500
rect 22772 6556 22836 6560
rect 22772 6500 22776 6556
rect 22776 6500 22832 6556
rect 22832 6500 22836 6556
rect 22772 6496 22836 6500
rect 22852 6556 22916 6560
rect 22852 6500 22856 6556
rect 22856 6500 22912 6556
rect 22912 6500 22916 6556
rect 22852 6496 22916 6500
rect 27612 6556 27676 6560
rect 27612 6500 27616 6556
rect 27616 6500 27672 6556
rect 27672 6500 27676 6556
rect 27612 6496 27676 6500
rect 27692 6556 27756 6560
rect 27692 6500 27696 6556
rect 27696 6500 27752 6556
rect 27752 6500 27756 6556
rect 27692 6496 27756 6500
rect 27772 6556 27836 6560
rect 27772 6500 27776 6556
rect 27776 6500 27832 6556
rect 27832 6500 27836 6556
rect 27772 6496 27836 6500
rect 27852 6556 27916 6560
rect 27852 6500 27856 6556
rect 27856 6500 27912 6556
rect 27912 6500 27916 6556
rect 27852 6496 27916 6500
rect 32612 6556 32676 6560
rect 32612 6500 32616 6556
rect 32616 6500 32672 6556
rect 32672 6500 32676 6556
rect 32612 6496 32676 6500
rect 32692 6556 32756 6560
rect 32692 6500 32696 6556
rect 32696 6500 32752 6556
rect 32752 6500 32756 6556
rect 32692 6496 32756 6500
rect 32772 6556 32836 6560
rect 32772 6500 32776 6556
rect 32776 6500 32832 6556
rect 32832 6500 32836 6556
rect 32772 6496 32836 6500
rect 32852 6556 32916 6560
rect 32852 6500 32856 6556
rect 32856 6500 32912 6556
rect 32912 6500 32916 6556
rect 32852 6496 32916 6500
rect 37612 6556 37676 6560
rect 37612 6500 37616 6556
rect 37616 6500 37672 6556
rect 37672 6500 37676 6556
rect 37612 6496 37676 6500
rect 37692 6556 37756 6560
rect 37692 6500 37696 6556
rect 37696 6500 37752 6556
rect 37752 6500 37756 6556
rect 37692 6496 37756 6500
rect 37772 6556 37836 6560
rect 37772 6500 37776 6556
rect 37776 6500 37832 6556
rect 37832 6500 37836 6556
rect 37772 6496 37836 6500
rect 37852 6556 37916 6560
rect 37852 6500 37856 6556
rect 37856 6500 37912 6556
rect 37912 6500 37916 6556
rect 37852 6496 37916 6500
rect 1952 6012 2016 6016
rect 1952 5956 1956 6012
rect 1956 5956 2012 6012
rect 2012 5956 2016 6012
rect 1952 5952 2016 5956
rect 2032 6012 2096 6016
rect 2032 5956 2036 6012
rect 2036 5956 2092 6012
rect 2092 5956 2096 6012
rect 2032 5952 2096 5956
rect 2112 6012 2176 6016
rect 2112 5956 2116 6012
rect 2116 5956 2172 6012
rect 2172 5956 2176 6012
rect 2112 5952 2176 5956
rect 2192 6012 2256 6016
rect 2192 5956 2196 6012
rect 2196 5956 2252 6012
rect 2252 5956 2256 6012
rect 2192 5952 2256 5956
rect 6952 6012 7016 6016
rect 6952 5956 6956 6012
rect 6956 5956 7012 6012
rect 7012 5956 7016 6012
rect 6952 5952 7016 5956
rect 7032 6012 7096 6016
rect 7032 5956 7036 6012
rect 7036 5956 7092 6012
rect 7092 5956 7096 6012
rect 7032 5952 7096 5956
rect 7112 6012 7176 6016
rect 7112 5956 7116 6012
rect 7116 5956 7172 6012
rect 7172 5956 7176 6012
rect 7112 5952 7176 5956
rect 7192 6012 7256 6016
rect 7192 5956 7196 6012
rect 7196 5956 7252 6012
rect 7252 5956 7256 6012
rect 7192 5952 7256 5956
rect 11952 6012 12016 6016
rect 11952 5956 11956 6012
rect 11956 5956 12012 6012
rect 12012 5956 12016 6012
rect 11952 5952 12016 5956
rect 12032 6012 12096 6016
rect 12032 5956 12036 6012
rect 12036 5956 12092 6012
rect 12092 5956 12096 6012
rect 12032 5952 12096 5956
rect 12112 6012 12176 6016
rect 12112 5956 12116 6012
rect 12116 5956 12172 6012
rect 12172 5956 12176 6012
rect 12112 5952 12176 5956
rect 12192 6012 12256 6016
rect 12192 5956 12196 6012
rect 12196 5956 12252 6012
rect 12252 5956 12256 6012
rect 12192 5952 12256 5956
rect 16952 6012 17016 6016
rect 16952 5956 16956 6012
rect 16956 5956 17012 6012
rect 17012 5956 17016 6012
rect 16952 5952 17016 5956
rect 17032 6012 17096 6016
rect 17032 5956 17036 6012
rect 17036 5956 17092 6012
rect 17092 5956 17096 6012
rect 17032 5952 17096 5956
rect 17112 6012 17176 6016
rect 17112 5956 17116 6012
rect 17116 5956 17172 6012
rect 17172 5956 17176 6012
rect 17112 5952 17176 5956
rect 17192 6012 17256 6016
rect 17192 5956 17196 6012
rect 17196 5956 17252 6012
rect 17252 5956 17256 6012
rect 17192 5952 17256 5956
rect 21952 6012 22016 6016
rect 21952 5956 21956 6012
rect 21956 5956 22012 6012
rect 22012 5956 22016 6012
rect 21952 5952 22016 5956
rect 22032 6012 22096 6016
rect 22032 5956 22036 6012
rect 22036 5956 22092 6012
rect 22092 5956 22096 6012
rect 22032 5952 22096 5956
rect 22112 6012 22176 6016
rect 22112 5956 22116 6012
rect 22116 5956 22172 6012
rect 22172 5956 22176 6012
rect 22112 5952 22176 5956
rect 22192 6012 22256 6016
rect 22192 5956 22196 6012
rect 22196 5956 22252 6012
rect 22252 5956 22256 6012
rect 22192 5952 22256 5956
rect 26952 6012 27016 6016
rect 26952 5956 26956 6012
rect 26956 5956 27012 6012
rect 27012 5956 27016 6012
rect 26952 5952 27016 5956
rect 27032 6012 27096 6016
rect 27032 5956 27036 6012
rect 27036 5956 27092 6012
rect 27092 5956 27096 6012
rect 27032 5952 27096 5956
rect 27112 6012 27176 6016
rect 27112 5956 27116 6012
rect 27116 5956 27172 6012
rect 27172 5956 27176 6012
rect 27112 5952 27176 5956
rect 27192 6012 27256 6016
rect 27192 5956 27196 6012
rect 27196 5956 27252 6012
rect 27252 5956 27256 6012
rect 27192 5952 27256 5956
rect 31952 6012 32016 6016
rect 31952 5956 31956 6012
rect 31956 5956 32012 6012
rect 32012 5956 32016 6012
rect 31952 5952 32016 5956
rect 32032 6012 32096 6016
rect 32032 5956 32036 6012
rect 32036 5956 32092 6012
rect 32092 5956 32096 6012
rect 32032 5952 32096 5956
rect 32112 6012 32176 6016
rect 32112 5956 32116 6012
rect 32116 5956 32172 6012
rect 32172 5956 32176 6012
rect 32112 5952 32176 5956
rect 32192 6012 32256 6016
rect 32192 5956 32196 6012
rect 32196 5956 32252 6012
rect 32252 5956 32256 6012
rect 32192 5952 32256 5956
rect 36952 6012 37016 6016
rect 36952 5956 36956 6012
rect 36956 5956 37012 6012
rect 37012 5956 37016 6012
rect 36952 5952 37016 5956
rect 37032 6012 37096 6016
rect 37032 5956 37036 6012
rect 37036 5956 37092 6012
rect 37092 5956 37096 6012
rect 37032 5952 37096 5956
rect 37112 6012 37176 6016
rect 37112 5956 37116 6012
rect 37116 5956 37172 6012
rect 37172 5956 37176 6012
rect 37112 5952 37176 5956
rect 37192 6012 37256 6016
rect 37192 5956 37196 6012
rect 37196 5956 37252 6012
rect 37252 5956 37256 6012
rect 37192 5952 37256 5956
rect 2612 5468 2676 5472
rect 2612 5412 2616 5468
rect 2616 5412 2672 5468
rect 2672 5412 2676 5468
rect 2612 5408 2676 5412
rect 2692 5468 2756 5472
rect 2692 5412 2696 5468
rect 2696 5412 2752 5468
rect 2752 5412 2756 5468
rect 2692 5408 2756 5412
rect 2772 5468 2836 5472
rect 2772 5412 2776 5468
rect 2776 5412 2832 5468
rect 2832 5412 2836 5468
rect 2772 5408 2836 5412
rect 2852 5468 2916 5472
rect 2852 5412 2856 5468
rect 2856 5412 2912 5468
rect 2912 5412 2916 5468
rect 2852 5408 2916 5412
rect 7612 5468 7676 5472
rect 7612 5412 7616 5468
rect 7616 5412 7672 5468
rect 7672 5412 7676 5468
rect 7612 5408 7676 5412
rect 7692 5468 7756 5472
rect 7692 5412 7696 5468
rect 7696 5412 7752 5468
rect 7752 5412 7756 5468
rect 7692 5408 7756 5412
rect 7772 5468 7836 5472
rect 7772 5412 7776 5468
rect 7776 5412 7832 5468
rect 7832 5412 7836 5468
rect 7772 5408 7836 5412
rect 7852 5468 7916 5472
rect 7852 5412 7856 5468
rect 7856 5412 7912 5468
rect 7912 5412 7916 5468
rect 7852 5408 7916 5412
rect 12612 5468 12676 5472
rect 12612 5412 12616 5468
rect 12616 5412 12672 5468
rect 12672 5412 12676 5468
rect 12612 5408 12676 5412
rect 12692 5468 12756 5472
rect 12692 5412 12696 5468
rect 12696 5412 12752 5468
rect 12752 5412 12756 5468
rect 12692 5408 12756 5412
rect 12772 5468 12836 5472
rect 12772 5412 12776 5468
rect 12776 5412 12832 5468
rect 12832 5412 12836 5468
rect 12772 5408 12836 5412
rect 12852 5468 12916 5472
rect 12852 5412 12856 5468
rect 12856 5412 12912 5468
rect 12912 5412 12916 5468
rect 12852 5408 12916 5412
rect 17612 5468 17676 5472
rect 17612 5412 17616 5468
rect 17616 5412 17672 5468
rect 17672 5412 17676 5468
rect 17612 5408 17676 5412
rect 17692 5468 17756 5472
rect 17692 5412 17696 5468
rect 17696 5412 17752 5468
rect 17752 5412 17756 5468
rect 17692 5408 17756 5412
rect 17772 5468 17836 5472
rect 17772 5412 17776 5468
rect 17776 5412 17832 5468
rect 17832 5412 17836 5468
rect 17772 5408 17836 5412
rect 17852 5468 17916 5472
rect 17852 5412 17856 5468
rect 17856 5412 17912 5468
rect 17912 5412 17916 5468
rect 17852 5408 17916 5412
rect 22612 5468 22676 5472
rect 22612 5412 22616 5468
rect 22616 5412 22672 5468
rect 22672 5412 22676 5468
rect 22612 5408 22676 5412
rect 22692 5468 22756 5472
rect 22692 5412 22696 5468
rect 22696 5412 22752 5468
rect 22752 5412 22756 5468
rect 22692 5408 22756 5412
rect 22772 5468 22836 5472
rect 22772 5412 22776 5468
rect 22776 5412 22832 5468
rect 22832 5412 22836 5468
rect 22772 5408 22836 5412
rect 22852 5468 22916 5472
rect 22852 5412 22856 5468
rect 22856 5412 22912 5468
rect 22912 5412 22916 5468
rect 22852 5408 22916 5412
rect 27612 5468 27676 5472
rect 27612 5412 27616 5468
rect 27616 5412 27672 5468
rect 27672 5412 27676 5468
rect 27612 5408 27676 5412
rect 27692 5468 27756 5472
rect 27692 5412 27696 5468
rect 27696 5412 27752 5468
rect 27752 5412 27756 5468
rect 27692 5408 27756 5412
rect 27772 5468 27836 5472
rect 27772 5412 27776 5468
rect 27776 5412 27832 5468
rect 27832 5412 27836 5468
rect 27772 5408 27836 5412
rect 27852 5468 27916 5472
rect 27852 5412 27856 5468
rect 27856 5412 27912 5468
rect 27912 5412 27916 5468
rect 27852 5408 27916 5412
rect 32612 5468 32676 5472
rect 32612 5412 32616 5468
rect 32616 5412 32672 5468
rect 32672 5412 32676 5468
rect 32612 5408 32676 5412
rect 32692 5468 32756 5472
rect 32692 5412 32696 5468
rect 32696 5412 32752 5468
rect 32752 5412 32756 5468
rect 32692 5408 32756 5412
rect 32772 5468 32836 5472
rect 32772 5412 32776 5468
rect 32776 5412 32832 5468
rect 32832 5412 32836 5468
rect 32772 5408 32836 5412
rect 32852 5468 32916 5472
rect 32852 5412 32856 5468
rect 32856 5412 32912 5468
rect 32912 5412 32916 5468
rect 32852 5408 32916 5412
rect 37612 5468 37676 5472
rect 37612 5412 37616 5468
rect 37616 5412 37672 5468
rect 37672 5412 37676 5468
rect 37612 5408 37676 5412
rect 37692 5468 37756 5472
rect 37692 5412 37696 5468
rect 37696 5412 37752 5468
rect 37752 5412 37756 5468
rect 37692 5408 37756 5412
rect 37772 5468 37836 5472
rect 37772 5412 37776 5468
rect 37776 5412 37832 5468
rect 37832 5412 37836 5468
rect 37772 5408 37836 5412
rect 37852 5468 37916 5472
rect 37852 5412 37856 5468
rect 37856 5412 37912 5468
rect 37912 5412 37916 5468
rect 37852 5408 37916 5412
rect 1952 4924 2016 4928
rect 1952 4868 1956 4924
rect 1956 4868 2012 4924
rect 2012 4868 2016 4924
rect 1952 4864 2016 4868
rect 2032 4924 2096 4928
rect 2032 4868 2036 4924
rect 2036 4868 2092 4924
rect 2092 4868 2096 4924
rect 2032 4864 2096 4868
rect 2112 4924 2176 4928
rect 2112 4868 2116 4924
rect 2116 4868 2172 4924
rect 2172 4868 2176 4924
rect 2112 4864 2176 4868
rect 2192 4924 2256 4928
rect 2192 4868 2196 4924
rect 2196 4868 2252 4924
rect 2252 4868 2256 4924
rect 2192 4864 2256 4868
rect 6952 4924 7016 4928
rect 6952 4868 6956 4924
rect 6956 4868 7012 4924
rect 7012 4868 7016 4924
rect 6952 4864 7016 4868
rect 7032 4924 7096 4928
rect 7032 4868 7036 4924
rect 7036 4868 7092 4924
rect 7092 4868 7096 4924
rect 7032 4864 7096 4868
rect 7112 4924 7176 4928
rect 7112 4868 7116 4924
rect 7116 4868 7172 4924
rect 7172 4868 7176 4924
rect 7112 4864 7176 4868
rect 7192 4924 7256 4928
rect 7192 4868 7196 4924
rect 7196 4868 7252 4924
rect 7252 4868 7256 4924
rect 7192 4864 7256 4868
rect 11952 4924 12016 4928
rect 11952 4868 11956 4924
rect 11956 4868 12012 4924
rect 12012 4868 12016 4924
rect 11952 4864 12016 4868
rect 12032 4924 12096 4928
rect 12032 4868 12036 4924
rect 12036 4868 12092 4924
rect 12092 4868 12096 4924
rect 12032 4864 12096 4868
rect 12112 4924 12176 4928
rect 12112 4868 12116 4924
rect 12116 4868 12172 4924
rect 12172 4868 12176 4924
rect 12112 4864 12176 4868
rect 12192 4924 12256 4928
rect 12192 4868 12196 4924
rect 12196 4868 12252 4924
rect 12252 4868 12256 4924
rect 12192 4864 12256 4868
rect 16952 4924 17016 4928
rect 16952 4868 16956 4924
rect 16956 4868 17012 4924
rect 17012 4868 17016 4924
rect 16952 4864 17016 4868
rect 17032 4924 17096 4928
rect 17032 4868 17036 4924
rect 17036 4868 17092 4924
rect 17092 4868 17096 4924
rect 17032 4864 17096 4868
rect 17112 4924 17176 4928
rect 17112 4868 17116 4924
rect 17116 4868 17172 4924
rect 17172 4868 17176 4924
rect 17112 4864 17176 4868
rect 17192 4924 17256 4928
rect 17192 4868 17196 4924
rect 17196 4868 17252 4924
rect 17252 4868 17256 4924
rect 17192 4864 17256 4868
rect 21952 4924 22016 4928
rect 21952 4868 21956 4924
rect 21956 4868 22012 4924
rect 22012 4868 22016 4924
rect 21952 4864 22016 4868
rect 22032 4924 22096 4928
rect 22032 4868 22036 4924
rect 22036 4868 22092 4924
rect 22092 4868 22096 4924
rect 22032 4864 22096 4868
rect 22112 4924 22176 4928
rect 22112 4868 22116 4924
rect 22116 4868 22172 4924
rect 22172 4868 22176 4924
rect 22112 4864 22176 4868
rect 22192 4924 22256 4928
rect 22192 4868 22196 4924
rect 22196 4868 22252 4924
rect 22252 4868 22256 4924
rect 22192 4864 22256 4868
rect 26952 4924 27016 4928
rect 26952 4868 26956 4924
rect 26956 4868 27012 4924
rect 27012 4868 27016 4924
rect 26952 4864 27016 4868
rect 27032 4924 27096 4928
rect 27032 4868 27036 4924
rect 27036 4868 27092 4924
rect 27092 4868 27096 4924
rect 27032 4864 27096 4868
rect 27112 4924 27176 4928
rect 27112 4868 27116 4924
rect 27116 4868 27172 4924
rect 27172 4868 27176 4924
rect 27112 4864 27176 4868
rect 27192 4924 27256 4928
rect 27192 4868 27196 4924
rect 27196 4868 27252 4924
rect 27252 4868 27256 4924
rect 27192 4864 27256 4868
rect 31952 4924 32016 4928
rect 31952 4868 31956 4924
rect 31956 4868 32012 4924
rect 32012 4868 32016 4924
rect 31952 4864 32016 4868
rect 32032 4924 32096 4928
rect 32032 4868 32036 4924
rect 32036 4868 32092 4924
rect 32092 4868 32096 4924
rect 32032 4864 32096 4868
rect 32112 4924 32176 4928
rect 32112 4868 32116 4924
rect 32116 4868 32172 4924
rect 32172 4868 32176 4924
rect 32112 4864 32176 4868
rect 32192 4924 32256 4928
rect 32192 4868 32196 4924
rect 32196 4868 32252 4924
rect 32252 4868 32256 4924
rect 32192 4864 32256 4868
rect 36952 4924 37016 4928
rect 36952 4868 36956 4924
rect 36956 4868 37012 4924
rect 37012 4868 37016 4924
rect 36952 4864 37016 4868
rect 37032 4924 37096 4928
rect 37032 4868 37036 4924
rect 37036 4868 37092 4924
rect 37092 4868 37096 4924
rect 37032 4864 37096 4868
rect 37112 4924 37176 4928
rect 37112 4868 37116 4924
rect 37116 4868 37172 4924
rect 37172 4868 37176 4924
rect 37112 4864 37176 4868
rect 37192 4924 37256 4928
rect 37192 4868 37196 4924
rect 37196 4868 37252 4924
rect 37252 4868 37256 4924
rect 37192 4864 37256 4868
rect 2612 4380 2676 4384
rect 2612 4324 2616 4380
rect 2616 4324 2672 4380
rect 2672 4324 2676 4380
rect 2612 4320 2676 4324
rect 2692 4380 2756 4384
rect 2692 4324 2696 4380
rect 2696 4324 2752 4380
rect 2752 4324 2756 4380
rect 2692 4320 2756 4324
rect 2772 4380 2836 4384
rect 2772 4324 2776 4380
rect 2776 4324 2832 4380
rect 2832 4324 2836 4380
rect 2772 4320 2836 4324
rect 2852 4380 2916 4384
rect 2852 4324 2856 4380
rect 2856 4324 2912 4380
rect 2912 4324 2916 4380
rect 2852 4320 2916 4324
rect 7612 4380 7676 4384
rect 7612 4324 7616 4380
rect 7616 4324 7672 4380
rect 7672 4324 7676 4380
rect 7612 4320 7676 4324
rect 7692 4380 7756 4384
rect 7692 4324 7696 4380
rect 7696 4324 7752 4380
rect 7752 4324 7756 4380
rect 7692 4320 7756 4324
rect 7772 4380 7836 4384
rect 7772 4324 7776 4380
rect 7776 4324 7832 4380
rect 7832 4324 7836 4380
rect 7772 4320 7836 4324
rect 7852 4380 7916 4384
rect 7852 4324 7856 4380
rect 7856 4324 7912 4380
rect 7912 4324 7916 4380
rect 7852 4320 7916 4324
rect 12612 4380 12676 4384
rect 12612 4324 12616 4380
rect 12616 4324 12672 4380
rect 12672 4324 12676 4380
rect 12612 4320 12676 4324
rect 12692 4380 12756 4384
rect 12692 4324 12696 4380
rect 12696 4324 12752 4380
rect 12752 4324 12756 4380
rect 12692 4320 12756 4324
rect 12772 4380 12836 4384
rect 12772 4324 12776 4380
rect 12776 4324 12832 4380
rect 12832 4324 12836 4380
rect 12772 4320 12836 4324
rect 12852 4380 12916 4384
rect 12852 4324 12856 4380
rect 12856 4324 12912 4380
rect 12912 4324 12916 4380
rect 12852 4320 12916 4324
rect 17612 4380 17676 4384
rect 17612 4324 17616 4380
rect 17616 4324 17672 4380
rect 17672 4324 17676 4380
rect 17612 4320 17676 4324
rect 17692 4380 17756 4384
rect 17692 4324 17696 4380
rect 17696 4324 17752 4380
rect 17752 4324 17756 4380
rect 17692 4320 17756 4324
rect 17772 4380 17836 4384
rect 17772 4324 17776 4380
rect 17776 4324 17832 4380
rect 17832 4324 17836 4380
rect 17772 4320 17836 4324
rect 17852 4380 17916 4384
rect 17852 4324 17856 4380
rect 17856 4324 17912 4380
rect 17912 4324 17916 4380
rect 17852 4320 17916 4324
rect 22612 4380 22676 4384
rect 22612 4324 22616 4380
rect 22616 4324 22672 4380
rect 22672 4324 22676 4380
rect 22612 4320 22676 4324
rect 22692 4380 22756 4384
rect 22692 4324 22696 4380
rect 22696 4324 22752 4380
rect 22752 4324 22756 4380
rect 22692 4320 22756 4324
rect 22772 4380 22836 4384
rect 22772 4324 22776 4380
rect 22776 4324 22832 4380
rect 22832 4324 22836 4380
rect 22772 4320 22836 4324
rect 22852 4380 22916 4384
rect 22852 4324 22856 4380
rect 22856 4324 22912 4380
rect 22912 4324 22916 4380
rect 22852 4320 22916 4324
rect 27612 4380 27676 4384
rect 27612 4324 27616 4380
rect 27616 4324 27672 4380
rect 27672 4324 27676 4380
rect 27612 4320 27676 4324
rect 27692 4380 27756 4384
rect 27692 4324 27696 4380
rect 27696 4324 27752 4380
rect 27752 4324 27756 4380
rect 27692 4320 27756 4324
rect 27772 4380 27836 4384
rect 27772 4324 27776 4380
rect 27776 4324 27832 4380
rect 27832 4324 27836 4380
rect 27772 4320 27836 4324
rect 27852 4380 27916 4384
rect 27852 4324 27856 4380
rect 27856 4324 27912 4380
rect 27912 4324 27916 4380
rect 27852 4320 27916 4324
rect 32612 4380 32676 4384
rect 32612 4324 32616 4380
rect 32616 4324 32672 4380
rect 32672 4324 32676 4380
rect 32612 4320 32676 4324
rect 32692 4380 32756 4384
rect 32692 4324 32696 4380
rect 32696 4324 32752 4380
rect 32752 4324 32756 4380
rect 32692 4320 32756 4324
rect 32772 4380 32836 4384
rect 32772 4324 32776 4380
rect 32776 4324 32832 4380
rect 32832 4324 32836 4380
rect 32772 4320 32836 4324
rect 32852 4380 32916 4384
rect 32852 4324 32856 4380
rect 32856 4324 32912 4380
rect 32912 4324 32916 4380
rect 32852 4320 32916 4324
rect 37612 4380 37676 4384
rect 37612 4324 37616 4380
rect 37616 4324 37672 4380
rect 37672 4324 37676 4380
rect 37612 4320 37676 4324
rect 37692 4380 37756 4384
rect 37692 4324 37696 4380
rect 37696 4324 37752 4380
rect 37752 4324 37756 4380
rect 37692 4320 37756 4324
rect 37772 4380 37836 4384
rect 37772 4324 37776 4380
rect 37776 4324 37832 4380
rect 37832 4324 37836 4380
rect 37772 4320 37836 4324
rect 37852 4380 37916 4384
rect 37852 4324 37856 4380
rect 37856 4324 37912 4380
rect 37912 4324 37916 4380
rect 37852 4320 37916 4324
rect 1952 3836 2016 3840
rect 1952 3780 1956 3836
rect 1956 3780 2012 3836
rect 2012 3780 2016 3836
rect 1952 3776 2016 3780
rect 2032 3836 2096 3840
rect 2032 3780 2036 3836
rect 2036 3780 2092 3836
rect 2092 3780 2096 3836
rect 2032 3776 2096 3780
rect 2112 3836 2176 3840
rect 2112 3780 2116 3836
rect 2116 3780 2172 3836
rect 2172 3780 2176 3836
rect 2112 3776 2176 3780
rect 2192 3836 2256 3840
rect 2192 3780 2196 3836
rect 2196 3780 2252 3836
rect 2252 3780 2256 3836
rect 2192 3776 2256 3780
rect 6952 3836 7016 3840
rect 6952 3780 6956 3836
rect 6956 3780 7012 3836
rect 7012 3780 7016 3836
rect 6952 3776 7016 3780
rect 7032 3836 7096 3840
rect 7032 3780 7036 3836
rect 7036 3780 7092 3836
rect 7092 3780 7096 3836
rect 7032 3776 7096 3780
rect 7112 3836 7176 3840
rect 7112 3780 7116 3836
rect 7116 3780 7172 3836
rect 7172 3780 7176 3836
rect 7112 3776 7176 3780
rect 7192 3836 7256 3840
rect 7192 3780 7196 3836
rect 7196 3780 7252 3836
rect 7252 3780 7256 3836
rect 7192 3776 7256 3780
rect 11952 3836 12016 3840
rect 11952 3780 11956 3836
rect 11956 3780 12012 3836
rect 12012 3780 12016 3836
rect 11952 3776 12016 3780
rect 12032 3836 12096 3840
rect 12032 3780 12036 3836
rect 12036 3780 12092 3836
rect 12092 3780 12096 3836
rect 12032 3776 12096 3780
rect 12112 3836 12176 3840
rect 12112 3780 12116 3836
rect 12116 3780 12172 3836
rect 12172 3780 12176 3836
rect 12112 3776 12176 3780
rect 12192 3836 12256 3840
rect 12192 3780 12196 3836
rect 12196 3780 12252 3836
rect 12252 3780 12256 3836
rect 12192 3776 12256 3780
rect 16952 3836 17016 3840
rect 16952 3780 16956 3836
rect 16956 3780 17012 3836
rect 17012 3780 17016 3836
rect 16952 3776 17016 3780
rect 17032 3836 17096 3840
rect 17032 3780 17036 3836
rect 17036 3780 17092 3836
rect 17092 3780 17096 3836
rect 17032 3776 17096 3780
rect 17112 3836 17176 3840
rect 17112 3780 17116 3836
rect 17116 3780 17172 3836
rect 17172 3780 17176 3836
rect 17112 3776 17176 3780
rect 17192 3836 17256 3840
rect 17192 3780 17196 3836
rect 17196 3780 17252 3836
rect 17252 3780 17256 3836
rect 17192 3776 17256 3780
rect 21952 3836 22016 3840
rect 21952 3780 21956 3836
rect 21956 3780 22012 3836
rect 22012 3780 22016 3836
rect 21952 3776 22016 3780
rect 22032 3836 22096 3840
rect 22032 3780 22036 3836
rect 22036 3780 22092 3836
rect 22092 3780 22096 3836
rect 22032 3776 22096 3780
rect 22112 3836 22176 3840
rect 22112 3780 22116 3836
rect 22116 3780 22172 3836
rect 22172 3780 22176 3836
rect 22112 3776 22176 3780
rect 22192 3836 22256 3840
rect 22192 3780 22196 3836
rect 22196 3780 22252 3836
rect 22252 3780 22256 3836
rect 22192 3776 22256 3780
rect 26952 3836 27016 3840
rect 26952 3780 26956 3836
rect 26956 3780 27012 3836
rect 27012 3780 27016 3836
rect 26952 3776 27016 3780
rect 27032 3836 27096 3840
rect 27032 3780 27036 3836
rect 27036 3780 27092 3836
rect 27092 3780 27096 3836
rect 27032 3776 27096 3780
rect 27112 3836 27176 3840
rect 27112 3780 27116 3836
rect 27116 3780 27172 3836
rect 27172 3780 27176 3836
rect 27112 3776 27176 3780
rect 27192 3836 27256 3840
rect 27192 3780 27196 3836
rect 27196 3780 27252 3836
rect 27252 3780 27256 3836
rect 27192 3776 27256 3780
rect 31952 3836 32016 3840
rect 31952 3780 31956 3836
rect 31956 3780 32012 3836
rect 32012 3780 32016 3836
rect 31952 3776 32016 3780
rect 32032 3836 32096 3840
rect 32032 3780 32036 3836
rect 32036 3780 32092 3836
rect 32092 3780 32096 3836
rect 32032 3776 32096 3780
rect 32112 3836 32176 3840
rect 32112 3780 32116 3836
rect 32116 3780 32172 3836
rect 32172 3780 32176 3836
rect 32112 3776 32176 3780
rect 32192 3836 32256 3840
rect 32192 3780 32196 3836
rect 32196 3780 32252 3836
rect 32252 3780 32256 3836
rect 32192 3776 32256 3780
rect 36952 3836 37016 3840
rect 36952 3780 36956 3836
rect 36956 3780 37012 3836
rect 37012 3780 37016 3836
rect 36952 3776 37016 3780
rect 37032 3836 37096 3840
rect 37032 3780 37036 3836
rect 37036 3780 37092 3836
rect 37092 3780 37096 3836
rect 37032 3776 37096 3780
rect 37112 3836 37176 3840
rect 37112 3780 37116 3836
rect 37116 3780 37172 3836
rect 37172 3780 37176 3836
rect 37112 3776 37176 3780
rect 37192 3836 37256 3840
rect 37192 3780 37196 3836
rect 37196 3780 37252 3836
rect 37252 3780 37256 3836
rect 37192 3776 37256 3780
rect 2612 3292 2676 3296
rect 2612 3236 2616 3292
rect 2616 3236 2672 3292
rect 2672 3236 2676 3292
rect 2612 3232 2676 3236
rect 2692 3292 2756 3296
rect 2692 3236 2696 3292
rect 2696 3236 2752 3292
rect 2752 3236 2756 3292
rect 2692 3232 2756 3236
rect 2772 3292 2836 3296
rect 2772 3236 2776 3292
rect 2776 3236 2832 3292
rect 2832 3236 2836 3292
rect 2772 3232 2836 3236
rect 2852 3292 2916 3296
rect 2852 3236 2856 3292
rect 2856 3236 2912 3292
rect 2912 3236 2916 3292
rect 2852 3232 2916 3236
rect 7612 3292 7676 3296
rect 7612 3236 7616 3292
rect 7616 3236 7672 3292
rect 7672 3236 7676 3292
rect 7612 3232 7676 3236
rect 7692 3292 7756 3296
rect 7692 3236 7696 3292
rect 7696 3236 7752 3292
rect 7752 3236 7756 3292
rect 7692 3232 7756 3236
rect 7772 3292 7836 3296
rect 7772 3236 7776 3292
rect 7776 3236 7832 3292
rect 7832 3236 7836 3292
rect 7772 3232 7836 3236
rect 7852 3292 7916 3296
rect 7852 3236 7856 3292
rect 7856 3236 7912 3292
rect 7912 3236 7916 3292
rect 7852 3232 7916 3236
rect 12612 3292 12676 3296
rect 12612 3236 12616 3292
rect 12616 3236 12672 3292
rect 12672 3236 12676 3292
rect 12612 3232 12676 3236
rect 12692 3292 12756 3296
rect 12692 3236 12696 3292
rect 12696 3236 12752 3292
rect 12752 3236 12756 3292
rect 12692 3232 12756 3236
rect 12772 3292 12836 3296
rect 12772 3236 12776 3292
rect 12776 3236 12832 3292
rect 12832 3236 12836 3292
rect 12772 3232 12836 3236
rect 12852 3292 12916 3296
rect 12852 3236 12856 3292
rect 12856 3236 12912 3292
rect 12912 3236 12916 3292
rect 12852 3232 12916 3236
rect 17612 3292 17676 3296
rect 17612 3236 17616 3292
rect 17616 3236 17672 3292
rect 17672 3236 17676 3292
rect 17612 3232 17676 3236
rect 17692 3292 17756 3296
rect 17692 3236 17696 3292
rect 17696 3236 17752 3292
rect 17752 3236 17756 3292
rect 17692 3232 17756 3236
rect 17772 3292 17836 3296
rect 17772 3236 17776 3292
rect 17776 3236 17832 3292
rect 17832 3236 17836 3292
rect 17772 3232 17836 3236
rect 17852 3292 17916 3296
rect 17852 3236 17856 3292
rect 17856 3236 17912 3292
rect 17912 3236 17916 3292
rect 17852 3232 17916 3236
rect 22612 3292 22676 3296
rect 22612 3236 22616 3292
rect 22616 3236 22672 3292
rect 22672 3236 22676 3292
rect 22612 3232 22676 3236
rect 22692 3292 22756 3296
rect 22692 3236 22696 3292
rect 22696 3236 22752 3292
rect 22752 3236 22756 3292
rect 22692 3232 22756 3236
rect 22772 3292 22836 3296
rect 22772 3236 22776 3292
rect 22776 3236 22832 3292
rect 22832 3236 22836 3292
rect 22772 3232 22836 3236
rect 22852 3292 22916 3296
rect 22852 3236 22856 3292
rect 22856 3236 22912 3292
rect 22912 3236 22916 3292
rect 22852 3232 22916 3236
rect 27612 3292 27676 3296
rect 27612 3236 27616 3292
rect 27616 3236 27672 3292
rect 27672 3236 27676 3292
rect 27612 3232 27676 3236
rect 27692 3292 27756 3296
rect 27692 3236 27696 3292
rect 27696 3236 27752 3292
rect 27752 3236 27756 3292
rect 27692 3232 27756 3236
rect 27772 3292 27836 3296
rect 27772 3236 27776 3292
rect 27776 3236 27832 3292
rect 27832 3236 27836 3292
rect 27772 3232 27836 3236
rect 27852 3292 27916 3296
rect 27852 3236 27856 3292
rect 27856 3236 27912 3292
rect 27912 3236 27916 3292
rect 27852 3232 27916 3236
rect 32612 3292 32676 3296
rect 32612 3236 32616 3292
rect 32616 3236 32672 3292
rect 32672 3236 32676 3292
rect 32612 3232 32676 3236
rect 32692 3292 32756 3296
rect 32692 3236 32696 3292
rect 32696 3236 32752 3292
rect 32752 3236 32756 3292
rect 32692 3232 32756 3236
rect 32772 3292 32836 3296
rect 32772 3236 32776 3292
rect 32776 3236 32832 3292
rect 32832 3236 32836 3292
rect 32772 3232 32836 3236
rect 32852 3292 32916 3296
rect 32852 3236 32856 3292
rect 32856 3236 32912 3292
rect 32912 3236 32916 3292
rect 32852 3232 32916 3236
rect 37612 3292 37676 3296
rect 37612 3236 37616 3292
rect 37616 3236 37672 3292
rect 37672 3236 37676 3292
rect 37612 3232 37676 3236
rect 37692 3292 37756 3296
rect 37692 3236 37696 3292
rect 37696 3236 37752 3292
rect 37752 3236 37756 3292
rect 37692 3232 37756 3236
rect 37772 3292 37836 3296
rect 37772 3236 37776 3292
rect 37776 3236 37832 3292
rect 37832 3236 37836 3292
rect 37772 3232 37836 3236
rect 37852 3292 37916 3296
rect 37852 3236 37856 3292
rect 37856 3236 37912 3292
rect 37912 3236 37916 3292
rect 37852 3232 37916 3236
rect 1952 2748 2016 2752
rect 1952 2692 1956 2748
rect 1956 2692 2012 2748
rect 2012 2692 2016 2748
rect 1952 2688 2016 2692
rect 2032 2748 2096 2752
rect 2032 2692 2036 2748
rect 2036 2692 2092 2748
rect 2092 2692 2096 2748
rect 2032 2688 2096 2692
rect 2112 2748 2176 2752
rect 2112 2692 2116 2748
rect 2116 2692 2172 2748
rect 2172 2692 2176 2748
rect 2112 2688 2176 2692
rect 2192 2748 2256 2752
rect 2192 2692 2196 2748
rect 2196 2692 2252 2748
rect 2252 2692 2256 2748
rect 2192 2688 2256 2692
rect 6952 2748 7016 2752
rect 6952 2692 6956 2748
rect 6956 2692 7012 2748
rect 7012 2692 7016 2748
rect 6952 2688 7016 2692
rect 7032 2748 7096 2752
rect 7032 2692 7036 2748
rect 7036 2692 7092 2748
rect 7092 2692 7096 2748
rect 7032 2688 7096 2692
rect 7112 2748 7176 2752
rect 7112 2692 7116 2748
rect 7116 2692 7172 2748
rect 7172 2692 7176 2748
rect 7112 2688 7176 2692
rect 7192 2748 7256 2752
rect 7192 2692 7196 2748
rect 7196 2692 7252 2748
rect 7252 2692 7256 2748
rect 7192 2688 7256 2692
rect 11952 2748 12016 2752
rect 11952 2692 11956 2748
rect 11956 2692 12012 2748
rect 12012 2692 12016 2748
rect 11952 2688 12016 2692
rect 12032 2748 12096 2752
rect 12032 2692 12036 2748
rect 12036 2692 12092 2748
rect 12092 2692 12096 2748
rect 12032 2688 12096 2692
rect 12112 2748 12176 2752
rect 12112 2692 12116 2748
rect 12116 2692 12172 2748
rect 12172 2692 12176 2748
rect 12112 2688 12176 2692
rect 12192 2748 12256 2752
rect 12192 2692 12196 2748
rect 12196 2692 12252 2748
rect 12252 2692 12256 2748
rect 12192 2688 12256 2692
rect 16952 2748 17016 2752
rect 16952 2692 16956 2748
rect 16956 2692 17012 2748
rect 17012 2692 17016 2748
rect 16952 2688 17016 2692
rect 17032 2748 17096 2752
rect 17032 2692 17036 2748
rect 17036 2692 17092 2748
rect 17092 2692 17096 2748
rect 17032 2688 17096 2692
rect 17112 2748 17176 2752
rect 17112 2692 17116 2748
rect 17116 2692 17172 2748
rect 17172 2692 17176 2748
rect 17112 2688 17176 2692
rect 17192 2748 17256 2752
rect 17192 2692 17196 2748
rect 17196 2692 17252 2748
rect 17252 2692 17256 2748
rect 17192 2688 17256 2692
rect 21952 2748 22016 2752
rect 21952 2692 21956 2748
rect 21956 2692 22012 2748
rect 22012 2692 22016 2748
rect 21952 2688 22016 2692
rect 22032 2748 22096 2752
rect 22032 2692 22036 2748
rect 22036 2692 22092 2748
rect 22092 2692 22096 2748
rect 22032 2688 22096 2692
rect 22112 2748 22176 2752
rect 22112 2692 22116 2748
rect 22116 2692 22172 2748
rect 22172 2692 22176 2748
rect 22112 2688 22176 2692
rect 22192 2748 22256 2752
rect 22192 2692 22196 2748
rect 22196 2692 22252 2748
rect 22252 2692 22256 2748
rect 22192 2688 22256 2692
rect 26952 2748 27016 2752
rect 26952 2692 26956 2748
rect 26956 2692 27012 2748
rect 27012 2692 27016 2748
rect 26952 2688 27016 2692
rect 27032 2748 27096 2752
rect 27032 2692 27036 2748
rect 27036 2692 27092 2748
rect 27092 2692 27096 2748
rect 27032 2688 27096 2692
rect 27112 2748 27176 2752
rect 27112 2692 27116 2748
rect 27116 2692 27172 2748
rect 27172 2692 27176 2748
rect 27112 2688 27176 2692
rect 27192 2748 27256 2752
rect 27192 2692 27196 2748
rect 27196 2692 27252 2748
rect 27252 2692 27256 2748
rect 27192 2688 27256 2692
rect 31952 2748 32016 2752
rect 31952 2692 31956 2748
rect 31956 2692 32012 2748
rect 32012 2692 32016 2748
rect 31952 2688 32016 2692
rect 32032 2748 32096 2752
rect 32032 2692 32036 2748
rect 32036 2692 32092 2748
rect 32092 2692 32096 2748
rect 32032 2688 32096 2692
rect 32112 2748 32176 2752
rect 32112 2692 32116 2748
rect 32116 2692 32172 2748
rect 32172 2692 32176 2748
rect 32112 2688 32176 2692
rect 32192 2748 32256 2752
rect 32192 2692 32196 2748
rect 32196 2692 32252 2748
rect 32252 2692 32256 2748
rect 32192 2688 32256 2692
rect 36952 2748 37016 2752
rect 36952 2692 36956 2748
rect 36956 2692 37012 2748
rect 37012 2692 37016 2748
rect 36952 2688 37016 2692
rect 37032 2748 37096 2752
rect 37032 2692 37036 2748
rect 37036 2692 37092 2748
rect 37092 2692 37096 2748
rect 37032 2688 37096 2692
rect 37112 2748 37176 2752
rect 37112 2692 37116 2748
rect 37116 2692 37172 2748
rect 37172 2692 37176 2748
rect 37112 2688 37176 2692
rect 37192 2748 37256 2752
rect 37192 2692 37196 2748
rect 37196 2692 37252 2748
rect 37252 2692 37256 2748
rect 37192 2688 37256 2692
rect 16436 2348 16500 2412
rect 2612 2204 2676 2208
rect 2612 2148 2616 2204
rect 2616 2148 2672 2204
rect 2672 2148 2676 2204
rect 2612 2144 2676 2148
rect 2692 2204 2756 2208
rect 2692 2148 2696 2204
rect 2696 2148 2752 2204
rect 2752 2148 2756 2204
rect 2692 2144 2756 2148
rect 2772 2204 2836 2208
rect 2772 2148 2776 2204
rect 2776 2148 2832 2204
rect 2832 2148 2836 2204
rect 2772 2144 2836 2148
rect 2852 2204 2916 2208
rect 2852 2148 2856 2204
rect 2856 2148 2912 2204
rect 2912 2148 2916 2204
rect 2852 2144 2916 2148
rect 7612 2204 7676 2208
rect 7612 2148 7616 2204
rect 7616 2148 7672 2204
rect 7672 2148 7676 2204
rect 7612 2144 7676 2148
rect 7692 2204 7756 2208
rect 7692 2148 7696 2204
rect 7696 2148 7752 2204
rect 7752 2148 7756 2204
rect 7692 2144 7756 2148
rect 7772 2204 7836 2208
rect 7772 2148 7776 2204
rect 7776 2148 7832 2204
rect 7832 2148 7836 2204
rect 7772 2144 7836 2148
rect 7852 2204 7916 2208
rect 7852 2148 7856 2204
rect 7856 2148 7912 2204
rect 7912 2148 7916 2204
rect 7852 2144 7916 2148
rect 12612 2204 12676 2208
rect 12612 2148 12616 2204
rect 12616 2148 12672 2204
rect 12672 2148 12676 2204
rect 12612 2144 12676 2148
rect 12692 2204 12756 2208
rect 12692 2148 12696 2204
rect 12696 2148 12752 2204
rect 12752 2148 12756 2204
rect 12692 2144 12756 2148
rect 12772 2204 12836 2208
rect 12772 2148 12776 2204
rect 12776 2148 12832 2204
rect 12832 2148 12836 2204
rect 12772 2144 12836 2148
rect 12852 2204 12916 2208
rect 12852 2148 12856 2204
rect 12856 2148 12912 2204
rect 12912 2148 12916 2204
rect 12852 2144 12916 2148
rect 17612 2204 17676 2208
rect 17612 2148 17616 2204
rect 17616 2148 17672 2204
rect 17672 2148 17676 2204
rect 17612 2144 17676 2148
rect 17692 2204 17756 2208
rect 17692 2148 17696 2204
rect 17696 2148 17752 2204
rect 17752 2148 17756 2204
rect 17692 2144 17756 2148
rect 17772 2204 17836 2208
rect 17772 2148 17776 2204
rect 17776 2148 17832 2204
rect 17832 2148 17836 2204
rect 17772 2144 17836 2148
rect 17852 2204 17916 2208
rect 17852 2148 17856 2204
rect 17856 2148 17912 2204
rect 17912 2148 17916 2204
rect 17852 2144 17916 2148
rect 22612 2204 22676 2208
rect 22612 2148 22616 2204
rect 22616 2148 22672 2204
rect 22672 2148 22676 2204
rect 22612 2144 22676 2148
rect 22692 2204 22756 2208
rect 22692 2148 22696 2204
rect 22696 2148 22752 2204
rect 22752 2148 22756 2204
rect 22692 2144 22756 2148
rect 22772 2204 22836 2208
rect 22772 2148 22776 2204
rect 22776 2148 22832 2204
rect 22832 2148 22836 2204
rect 22772 2144 22836 2148
rect 22852 2204 22916 2208
rect 22852 2148 22856 2204
rect 22856 2148 22912 2204
rect 22912 2148 22916 2204
rect 22852 2144 22916 2148
rect 27612 2204 27676 2208
rect 27612 2148 27616 2204
rect 27616 2148 27672 2204
rect 27672 2148 27676 2204
rect 27612 2144 27676 2148
rect 27692 2204 27756 2208
rect 27692 2148 27696 2204
rect 27696 2148 27752 2204
rect 27752 2148 27756 2204
rect 27692 2144 27756 2148
rect 27772 2204 27836 2208
rect 27772 2148 27776 2204
rect 27776 2148 27832 2204
rect 27832 2148 27836 2204
rect 27772 2144 27836 2148
rect 27852 2204 27916 2208
rect 27852 2148 27856 2204
rect 27856 2148 27912 2204
rect 27912 2148 27916 2204
rect 27852 2144 27916 2148
rect 32612 2204 32676 2208
rect 32612 2148 32616 2204
rect 32616 2148 32672 2204
rect 32672 2148 32676 2204
rect 32612 2144 32676 2148
rect 32692 2204 32756 2208
rect 32692 2148 32696 2204
rect 32696 2148 32752 2204
rect 32752 2148 32756 2204
rect 32692 2144 32756 2148
rect 32772 2204 32836 2208
rect 32772 2148 32776 2204
rect 32776 2148 32832 2204
rect 32832 2148 32836 2204
rect 32772 2144 32836 2148
rect 32852 2204 32916 2208
rect 32852 2148 32856 2204
rect 32856 2148 32912 2204
rect 32912 2148 32916 2204
rect 32852 2144 32916 2148
rect 37612 2204 37676 2208
rect 37612 2148 37616 2204
rect 37616 2148 37672 2204
rect 37672 2148 37676 2204
rect 37612 2144 37676 2148
rect 37692 2204 37756 2208
rect 37692 2148 37696 2204
rect 37696 2148 37752 2204
rect 37752 2148 37756 2204
rect 37692 2144 37756 2148
rect 37772 2204 37836 2208
rect 37772 2148 37776 2204
rect 37776 2148 37832 2204
rect 37832 2148 37836 2204
rect 37772 2144 37836 2148
rect 37852 2204 37916 2208
rect 37852 2148 37856 2204
rect 37856 2148 37912 2204
rect 37912 2148 37916 2204
rect 37852 2144 37916 2148
<< metal4 >>
rect 1944 69120 2264 69680
rect 1944 69056 1952 69120
rect 2016 69056 2032 69120
rect 2096 69056 2112 69120
rect 2176 69056 2192 69120
rect 2256 69056 2264 69120
rect 1944 68294 2264 69056
rect 1944 68058 1986 68294
rect 2222 68058 2264 68294
rect 1944 68032 2264 68058
rect 1944 67968 1952 68032
rect 2016 67968 2032 68032
rect 2096 67968 2112 68032
rect 2176 67968 2192 68032
rect 2256 67968 2264 68032
rect 1944 66944 2264 67968
rect 1944 66880 1952 66944
rect 2016 66880 2032 66944
rect 2096 66880 2112 66944
rect 2176 66880 2192 66944
rect 2256 66880 2264 66944
rect 1944 65856 2264 66880
rect 1944 65792 1952 65856
rect 2016 65792 2032 65856
rect 2096 65792 2112 65856
rect 2176 65792 2192 65856
rect 2256 65792 2264 65856
rect 1944 64768 2264 65792
rect 1944 64704 1952 64768
rect 2016 64704 2032 64768
rect 2096 64704 2112 64768
rect 2176 64704 2192 64768
rect 2256 64704 2264 64768
rect 1944 63680 2264 64704
rect 1944 63616 1952 63680
rect 2016 63616 2032 63680
rect 2096 63616 2112 63680
rect 2176 63616 2192 63680
rect 2256 63616 2264 63680
rect 1944 63294 2264 63616
rect 1944 63058 1986 63294
rect 2222 63058 2264 63294
rect 1944 62592 2264 63058
rect 1944 62528 1952 62592
rect 2016 62528 2032 62592
rect 2096 62528 2112 62592
rect 2176 62528 2192 62592
rect 2256 62528 2264 62592
rect 1944 61504 2264 62528
rect 1944 61440 1952 61504
rect 2016 61440 2032 61504
rect 2096 61440 2112 61504
rect 2176 61440 2192 61504
rect 2256 61440 2264 61504
rect 1944 60416 2264 61440
rect 1944 60352 1952 60416
rect 2016 60352 2032 60416
rect 2096 60352 2112 60416
rect 2176 60352 2192 60416
rect 2256 60352 2264 60416
rect 1944 59328 2264 60352
rect 1944 59264 1952 59328
rect 2016 59264 2032 59328
rect 2096 59264 2112 59328
rect 2176 59264 2192 59328
rect 2256 59264 2264 59328
rect 1944 58294 2264 59264
rect 1944 58240 1986 58294
rect 2222 58240 2264 58294
rect 1944 58176 1952 58240
rect 2256 58176 2264 58240
rect 1944 58058 1986 58176
rect 2222 58058 2264 58176
rect 1944 57152 2264 58058
rect 1944 57088 1952 57152
rect 2016 57088 2032 57152
rect 2096 57088 2112 57152
rect 2176 57088 2192 57152
rect 2256 57088 2264 57152
rect 1944 56064 2264 57088
rect 1944 56000 1952 56064
rect 2016 56000 2032 56064
rect 2096 56000 2112 56064
rect 2176 56000 2192 56064
rect 2256 56000 2264 56064
rect 1944 54976 2264 56000
rect 1944 54912 1952 54976
rect 2016 54912 2032 54976
rect 2096 54912 2112 54976
rect 2176 54912 2192 54976
rect 2256 54912 2264 54976
rect 1944 53888 2264 54912
rect 1944 53824 1952 53888
rect 2016 53824 2032 53888
rect 2096 53824 2112 53888
rect 2176 53824 2192 53888
rect 2256 53824 2264 53888
rect 1944 53294 2264 53824
rect 1944 53058 1986 53294
rect 2222 53058 2264 53294
rect 1944 52800 2264 53058
rect 1944 52736 1952 52800
rect 2016 52736 2032 52800
rect 2096 52736 2112 52800
rect 2176 52736 2192 52800
rect 2256 52736 2264 52800
rect 1944 51712 2264 52736
rect 1944 51648 1952 51712
rect 2016 51648 2032 51712
rect 2096 51648 2112 51712
rect 2176 51648 2192 51712
rect 2256 51648 2264 51712
rect 1944 50624 2264 51648
rect 1944 50560 1952 50624
rect 2016 50560 2032 50624
rect 2096 50560 2112 50624
rect 2176 50560 2192 50624
rect 2256 50560 2264 50624
rect 1944 49536 2264 50560
rect 1944 49472 1952 49536
rect 2016 49472 2032 49536
rect 2096 49472 2112 49536
rect 2176 49472 2192 49536
rect 2256 49472 2264 49536
rect 1944 48448 2264 49472
rect 1944 48384 1952 48448
rect 2016 48384 2032 48448
rect 2096 48384 2112 48448
rect 2176 48384 2192 48448
rect 2256 48384 2264 48448
rect 1944 48294 2264 48384
rect 1944 48058 1986 48294
rect 2222 48058 2264 48294
rect 1944 47360 2264 48058
rect 1944 47296 1952 47360
rect 2016 47296 2032 47360
rect 2096 47296 2112 47360
rect 2176 47296 2192 47360
rect 2256 47296 2264 47360
rect 1944 46272 2264 47296
rect 1944 46208 1952 46272
rect 2016 46208 2032 46272
rect 2096 46208 2112 46272
rect 2176 46208 2192 46272
rect 2256 46208 2264 46272
rect 1944 45184 2264 46208
rect 1944 45120 1952 45184
rect 2016 45120 2032 45184
rect 2096 45120 2112 45184
rect 2176 45120 2192 45184
rect 2256 45120 2264 45184
rect 1944 44096 2264 45120
rect 1944 44032 1952 44096
rect 2016 44032 2032 44096
rect 2096 44032 2112 44096
rect 2176 44032 2192 44096
rect 2256 44032 2264 44096
rect 1944 43294 2264 44032
rect 1944 43058 1986 43294
rect 2222 43058 2264 43294
rect 1944 43008 2264 43058
rect 1944 42944 1952 43008
rect 2016 42944 2032 43008
rect 2096 42944 2112 43008
rect 2176 42944 2192 43008
rect 2256 42944 2264 43008
rect 1944 41920 2264 42944
rect 1944 41856 1952 41920
rect 2016 41856 2032 41920
rect 2096 41856 2112 41920
rect 2176 41856 2192 41920
rect 2256 41856 2264 41920
rect 1944 40832 2264 41856
rect 1944 40768 1952 40832
rect 2016 40768 2032 40832
rect 2096 40768 2112 40832
rect 2176 40768 2192 40832
rect 2256 40768 2264 40832
rect 1944 39744 2264 40768
rect 1944 39680 1952 39744
rect 2016 39680 2032 39744
rect 2096 39680 2112 39744
rect 2176 39680 2192 39744
rect 2256 39680 2264 39744
rect 1944 38656 2264 39680
rect 1944 38592 1952 38656
rect 2016 38592 2032 38656
rect 2096 38592 2112 38656
rect 2176 38592 2192 38656
rect 2256 38592 2264 38656
rect 1944 38294 2264 38592
rect 1944 38058 1986 38294
rect 2222 38058 2264 38294
rect 1944 37568 2264 38058
rect 1944 37504 1952 37568
rect 2016 37504 2032 37568
rect 2096 37504 2112 37568
rect 2176 37504 2192 37568
rect 2256 37504 2264 37568
rect 1944 36480 2264 37504
rect 1944 36416 1952 36480
rect 2016 36416 2032 36480
rect 2096 36416 2112 36480
rect 2176 36416 2192 36480
rect 2256 36416 2264 36480
rect 1944 35392 2264 36416
rect 1944 35328 1952 35392
rect 2016 35328 2032 35392
rect 2096 35328 2112 35392
rect 2176 35328 2192 35392
rect 2256 35328 2264 35392
rect 1944 34304 2264 35328
rect 1944 34240 1952 34304
rect 2016 34240 2032 34304
rect 2096 34240 2112 34304
rect 2176 34240 2192 34304
rect 2256 34240 2264 34304
rect 1944 33294 2264 34240
rect 1944 33216 1986 33294
rect 2222 33216 2264 33294
rect 1944 33152 1952 33216
rect 2256 33152 2264 33216
rect 1944 33058 1986 33152
rect 2222 33058 2264 33152
rect 1944 32128 2264 33058
rect 1944 32064 1952 32128
rect 2016 32064 2032 32128
rect 2096 32064 2112 32128
rect 2176 32064 2192 32128
rect 2256 32064 2264 32128
rect 1944 31040 2264 32064
rect 1944 30976 1952 31040
rect 2016 30976 2032 31040
rect 2096 30976 2112 31040
rect 2176 30976 2192 31040
rect 2256 30976 2264 31040
rect 1944 29952 2264 30976
rect 1944 29888 1952 29952
rect 2016 29888 2032 29952
rect 2096 29888 2112 29952
rect 2176 29888 2192 29952
rect 2256 29888 2264 29952
rect 1944 28864 2264 29888
rect 1944 28800 1952 28864
rect 2016 28800 2032 28864
rect 2096 28800 2112 28864
rect 2176 28800 2192 28864
rect 2256 28800 2264 28864
rect 1944 28294 2264 28800
rect 1944 28058 1986 28294
rect 2222 28058 2264 28294
rect 1944 27776 2264 28058
rect 1944 27712 1952 27776
rect 2016 27712 2032 27776
rect 2096 27712 2112 27776
rect 2176 27712 2192 27776
rect 2256 27712 2264 27776
rect 1944 26688 2264 27712
rect 1944 26624 1952 26688
rect 2016 26624 2032 26688
rect 2096 26624 2112 26688
rect 2176 26624 2192 26688
rect 2256 26624 2264 26688
rect 1944 25600 2264 26624
rect 1944 25536 1952 25600
rect 2016 25536 2032 25600
rect 2096 25536 2112 25600
rect 2176 25536 2192 25600
rect 2256 25536 2264 25600
rect 1944 24512 2264 25536
rect 1944 24448 1952 24512
rect 2016 24448 2032 24512
rect 2096 24448 2112 24512
rect 2176 24448 2192 24512
rect 2256 24448 2264 24512
rect 1944 23424 2264 24448
rect 1944 23360 1952 23424
rect 2016 23360 2032 23424
rect 2096 23360 2112 23424
rect 2176 23360 2192 23424
rect 2256 23360 2264 23424
rect 1944 23294 2264 23360
rect 1944 23058 1986 23294
rect 2222 23058 2264 23294
rect 1944 22336 2264 23058
rect 1944 22272 1952 22336
rect 2016 22272 2032 22336
rect 2096 22272 2112 22336
rect 2176 22272 2192 22336
rect 2256 22272 2264 22336
rect 1944 21248 2264 22272
rect 1944 21184 1952 21248
rect 2016 21184 2032 21248
rect 2096 21184 2112 21248
rect 2176 21184 2192 21248
rect 2256 21184 2264 21248
rect 1944 20160 2264 21184
rect 1944 20096 1952 20160
rect 2016 20096 2032 20160
rect 2096 20096 2112 20160
rect 2176 20096 2192 20160
rect 2256 20096 2264 20160
rect 1944 19072 2264 20096
rect 1944 19008 1952 19072
rect 2016 19008 2032 19072
rect 2096 19008 2112 19072
rect 2176 19008 2192 19072
rect 2256 19008 2264 19072
rect 1944 18294 2264 19008
rect 1944 18058 1986 18294
rect 2222 18058 2264 18294
rect 1944 17984 2264 18058
rect 1944 17920 1952 17984
rect 2016 17920 2032 17984
rect 2096 17920 2112 17984
rect 2176 17920 2192 17984
rect 2256 17920 2264 17984
rect 1944 16896 2264 17920
rect 1944 16832 1952 16896
rect 2016 16832 2032 16896
rect 2096 16832 2112 16896
rect 2176 16832 2192 16896
rect 2256 16832 2264 16896
rect 1944 15808 2264 16832
rect 1944 15744 1952 15808
rect 2016 15744 2032 15808
rect 2096 15744 2112 15808
rect 2176 15744 2192 15808
rect 2256 15744 2264 15808
rect 1944 14720 2264 15744
rect 1944 14656 1952 14720
rect 2016 14656 2032 14720
rect 2096 14656 2112 14720
rect 2176 14656 2192 14720
rect 2256 14656 2264 14720
rect 1944 13632 2264 14656
rect 1944 13568 1952 13632
rect 2016 13568 2032 13632
rect 2096 13568 2112 13632
rect 2176 13568 2192 13632
rect 2256 13568 2264 13632
rect 1944 13294 2264 13568
rect 1944 13058 1986 13294
rect 2222 13058 2264 13294
rect 1944 12544 2264 13058
rect 1944 12480 1952 12544
rect 2016 12480 2032 12544
rect 2096 12480 2112 12544
rect 2176 12480 2192 12544
rect 2256 12480 2264 12544
rect 1944 11456 2264 12480
rect 1944 11392 1952 11456
rect 2016 11392 2032 11456
rect 2096 11392 2112 11456
rect 2176 11392 2192 11456
rect 2256 11392 2264 11456
rect 1944 10368 2264 11392
rect 1944 10304 1952 10368
rect 2016 10304 2032 10368
rect 2096 10304 2112 10368
rect 2176 10304 2192 10368
rect 2256 10304 2264 10368
rect 1944 9280 2264 10304
rect 1944 9216 1952 9280
rect 2016 9216 2032 9280
rect 2096 9216 2112 9280
rect 2176 9216 2192 9280
rect 2256 9216 2264 9280
rect 1944 8294 2264 9216
rect 1944 8192 1986 8294
rect 2222 8192 2264 8294
rect 1944 8128 1952 8192
rect 2256 8128 2264 8192
rect 1944 8058 1986 8128
rect 2222 8058 2264 8128
rect 1944 7104 2264 8058
rect 1944 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2264 7104
rect 1944 6016 2264 7040
rect 1944 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2264 6016
rect 1944 4928 2264 5952
rect 1944 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2264 4928
rect 1944 3840 2264 4864
rect 1944 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2264 3840
rect 1944 3294 2264 3776
rect 1944 3058 1986 3294
rect 2222 3058 2264 3294
rect 1944 2752 2264 3058
rect 1944 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2264 2752
rect 1944 2128 2264 2688
rect 2604 69664 2924 69680
rect 2604 69600 2612 69664
rect 2676 69600 2692 69664
rect 2756 69600 2772 69664
rect 2836 69600 2852 69664
rect 2916 69600 2924 69664
rect 2604 68954 2924 69600
rect 2604 68718 2646 68954
rect 2882 68718 2924 68954
rect 2604 68576 2924 68718
rect 2604 68512 2612 68576
rect 2676 68512 2692 68576
rect 2756 68512 2772 68576
rect 2836 68512 2852 68576
rect 2916 68512 2924 68576
rect 2604 67488 2924 68512
rect 6944 69120 7264 69680
rect 6944 69056 6952 69120
rect 7016 69056 7032 69120
rect 7096 69056 7112 69120
rect 7176 69056 7192 69120
rect 7256 69056 7264 69120
rect 6944 68294 7264 69056
rect 6944 68058 6986 68294
rect 7222 68058 7264 68294
rect 6944 68032 7264 68058
rect 6944 67968 6952 68032
rect 7016 67968 7032 68032
rect 7096 67968 7112 68032
rect 7176 67968 7192 68032
rect 7256 67968 7264 68032
rect 3371 67692 3437 67693
rect 3371 67628 3372 67692
rect 3436 67628 3437 67692
rect 3371 67627 3437 67628
rect 2604 67424 2612 67488
rect 2676 67424 2692 67488
rect 2756 67424 2772 67488
rect 2836 67424 2852 67488
rect 2916 67424 2924 67488
rect 2604 66400 2924 67424
rect 2604 66336 2612 66400
rect 2676 66336 2692 66400
rect 2756 66336 2772 66400
rect 2836 66336 2852 66400
rect 2916 66336 2924 66400
rect 2604 65312 2924 66336
rect 2604 65248 2612 65312
rect 2676 65248 2692 65312
rect 2756 65248 2772 65312
rect 2836 65248 2852 65312
rect 2916 65248 2924 65312
rect 2604 64224 2924 65248
rect 2604 64160 2612 64224
rect 2676 64160 2692 64224
rect 2756 64160 2772 64224
rect 2836 64160 2852 64224
rect 2916 64160 2924 64224
rect 2604 63954 2924 64160
rect 2604 63718 2646 63954
rect 2882 63718 2924 63954
rect 2604 63136 2924 63718
rect 2604 63072 2612 63136
rect 2676 63072 2692 63136
rect 2756 63072 2772 63136
rect 2836 63072 2852 63136
rect 2916 63072 2924 63136
rect 2604 62048 2924 63072
rect 2604 61984 2612 62048
rect 2676 61984 2692 62048
rect 2756 61984 2772 62048
rect 2836 61984 2852 62048
rect 2916 61984 2924 62048
rect 2604 60960 2924 61984
rect 2604 60896 2612 60960
rect 2676 60896 2692 60960
rect 2756 60896 2772 60960
rect 2836 60896 2852 60960
rect 2916 60896 2924 60960
rect 2604 59872 2924 60896
rect 2604 59808 2612 59872
rect 2676 59808 2692 59872
rect 2756 59808 2772 59872
rect 2836 59808 2852 59872
rect 2916 59808 2924 59872
rect 2604 58954 2924 59808
rect 2604 58784 2646 58954
rect 2882 58784 2924 58954
rect 2604 58720 2612 58784
rect 2916 58720 2924 58784
rect 2604 58718 2646 58720
rect 2882 58718 2924 58720
rect 2604 57696 2924 58718
rect 2604 57632 2612 57696
rect 2676 57632 2692 57696
rect 2756 57632 2772 57696
rect 2836 57632 2852 57696
rect 2916 57632 2924 57696
rect 2604 56608 2924 57632
rect 2604 56544 2612 56608
rect 2676 56544 2692 56608
rect 2756 56544 2772 56608
rect 2836 56544 2852 56608
rect 2916 56544 2924 56608
rect 2604 55520 2924 56544
rect 2604 55456 2612 55520
rect 2676 55456 2692 55520
rect 2756 55456 2772 55520
rect 2836 55456 2852 55520
rect 2916 55456 2924 55520
rect 2604 54432 2924 55456
rect 2604 54368 2612 54432
rect 2676 54368 2692 54432
rect 2756 54368 2772 54432
rect 2836 54368 2852 54432
rect 2916 54368 2924 54432
rect 2604 53954 2924 54368
rect 2604 53718 2646 53954
rect 2882 53718 2924 53954
rect 2604 53344 2924 53718
rect 2604 53280 2612 53344
rect 2676 53280 2692 53344
rect 2756 53280 2772 53344
rect 2836 53280 2852 53344
rect 2916 53280 2924 53344
rect 2604 52256 2924 53280
rect 2604 52192 2612 52256
rect 2676 52192 2692 52256
rect 2756 52192 2772 52256
rect 2836 52192 2852 52256
rect 2916 52192 2924 52256
rect 2604 51168 2924 52192
rect 2604 51104 2612 51168
rect 2676 51104 2692 51168
rect 2756 51104 2772 51168
rect 2836 51104 2852 51168
rect 2916 51104 2924 51168
rect 2604 50080 2924 51104
rect 2604 50016 2612 50080
rect 2676 50016 2692 50080
rect 2756 50016 2772 50080
rect 2836 50016 2852 50080
rect 2916 50016 2924 50080
rect 2604 48992 2924 50016
rect 2604 48928 2612 48992
rect 2676 48954 2692 48992
rect 2756 48954 2772 48992
rect 2836 48954 2852 48992
rect 2916 48928 2924 48992
rect 2604 48718 2646 48928
rect 2882 48718 2924 48928
rect 2604 47904 2924 48718
rect 2604 47840 2612 47904
rect 2676 47840 2692 47904
rect 2756 47840 2772 47904
rect 2836 47840 2852 47904
rect 2916 47840 2924 47904
rect 2604 46816 2924 47840
rect 2604 46752 2612 46816
rect 2676 46752 2692 46816
rect 2756 46752 2772 46816
rect 2836 46752 2852 46816
rect 2916 46752 2924 46816
rect 2604 45728 2924 46752
rect 2604 45664 2612 45728
rect 2676 45664 2692 45728
rect 2756 45664 2772 45728
rect 2836 45664 2852 45728
rect 2916 45664 2924 45728
rect 2604 44640 2924 45664
rect 2604 44576 2612 44640
rect 2676 44576 2692 44640
rect 2756 44576 2772 44640
rect 2836 44576 2852 44640
rect 2916 44576 2924 44640
rect 2604 43954 2924 44576
rect 2604 43718 2646 43954
rect 2882 43718 2924 43954
rect 2604 43552 2924 43718
rect 2604 43488 2612 43552
rect 2676 43488 2692 43552
rect 2756 43488 2772 43552
rect 2836 43488 2852 43552
rect 2916 43488 2924 43552
rect 2604 42464 2924 43488
rect 2604 42400 2612 42464
rect 2676 42400 2692 42464
rect 2756 42400 2772 42464
rect 2836 42400 2852 42464
rect 2916 42400 2924 42464
rect 2604 41376 2924 42400
rect 2604 41312 2612 41376
rect 2676 41312 2692 41376
rect 2756 41312 2772 41376
rect 2836 41312 2852 41376
rect 2916 41312 2924 41376
rect 2604 40288 2924 41312
rect 2604 40224 2612 40288
rect 2676 40224 2692 40288
rect 2756 40224 2772 40288
rect 2836 40224 2852 40288
rect 2916 40224 2924 40288
rect 2604 39200 2924 40224
rect 2604 39136 2612 39200
rect 2676 39136 2692 39200
rect 2756 39136 2772 39200
rect 2836 39136 2852 39200
rect 2916 39136 2924 39200
rect 2604 38954 2924 39136
rect 2604 38718 2646 38954
rect 2882 38718 2924 38954
rect 2604 38112 2924 38718
rect 2604 38048 2612 38112
rect 2676 38048 2692 38112
rect 2756 38048 2772 38112
rect 2836 38048 2852 38112
rect 2916 38048 2924 38112
rect 2604 37024 2924 38048
rect 2604 36960 2612 37024
rect 2676 36960 2692 37024
rect 2756 36960 2772 37024
rect 2836 36960 2852 37024
rect 2916 36960 2924 37024
rect 2604 35936 2924 36960
rect 2604 35872 2612 35936
rect 2676 35872 2692 35936
rect 2756 35872 2772 35936
rect 2836 35872 2852 35936
rect 2916 35872 2924 35936
rect 2604 34848 2924 35872
rect 2604 34784 2612 34848
rect 2676 34784 2692 34848
rect 2756 34784 2772 34848
rect 2836 34784 2852 34848
rect 2916 34784 2924 34848
rect 2604 33954 2924 34784
rect 2604 33760 2646 33954
rect 2882 33760 2924 33954
rect 2604 33696 2612 33760
rect 2676 33696 2692 33718
rect 2756 33696 2772 33718
rect 2836 33696 2852 33718
rect 2916 33696 2924 33760
rect 2604 32672 2924 33696
rect 2604 32608 2612 32672
rect 2676 32608 2692 32672
rect 2756 32608 2772 32672
rect 2836 32608 2852 32672
rect 2916 32608 2924 32672
rect 2604 31584 2924 32608
rect 2604 31520 2612 31584
rect 2676 31520 2692 31584
rect 2756 31520 2772 31584
rect 2836 31520 2852 31584
rect 2916 31520 2924 31584
rect 2604 30496 2924 31520
rect 2604 30432 2612 30496
rect 2676 30432 2692 30496
rect 2756 30432 2772 30496
rect 2836 30432 2852 30496
rect 2916 30432 2924 30496
rect 2604 29408 2924 30432
rect 2604 29344 2612 29408
rect 2676 29344 2692 29408
rect 2756 29344 2772 29408
rect 2836 29344 2852 29408
rect 2916 29344 2924 29408
rect 2604 28954 2924 29344
rect 2604 28718 2646 28954
rect 2882 28718 2924 28954
rect 2604 28320 2924 28718
rect 2604 28256 2612 28320
rect 2676 28256 2692 28320
rect 2756 28256 2772 28320
rect 2836 28256 2852 28320
rect 2916 28256 2924 28320
rect 2604 27232 2924 28256
rect 2604 27168 2612 27232
rect 2676 27168 2692 27232
rect 2756 27168 2772 27232
rect 2836 27168 2852 27232
rect 2916 27168 2924 27232
rect 2604 26144 2924 27168
rect 2604 26080 2612 26144
rect 2676 26080 2692 26144
rect 2756 26080 2772 26144
rect 2836 26080 2852 26144
rect 2916 26080 2924 26144
rect 2604 25056 2924 26080
rect 2604 24992 2612 25056
rect 2676 24992 2692 25056
rect 2756 24992 2772 25056
rect 2836 24992 2852 25056
rect 2916 24992 2924 25056
rect 2604 23968 2924 24992
rect 2604 23904 2612 23968
rect 2676 23954 2692 23968
rect 2756 23954 2772 23968
rect 2836 23954 2852 23968
rect 2916 23904 2924 23968
rect 2604 23718 2646 23904
rect 2882 23718 2924 23904
rect 2604 22880 2924 23718
rect 2604 22816 2612 22880
rect 2676 22816 2692 22880
rect 2756 22816 2772 22880
rect 2836 22816 2852 22880
rect 2916 22816 2924 22880
rect 2604 21792 2924 22816
rect 2604 21728 2612 21792
rect 2676 21728 2692 21792
rect 2756 21728 2772 21792
rect 2836 21728 2852 21792
rect 2916 21728 2924 21792
rect 2604 20704 2924 21728
rect 2604 20640 2612 20704
rect 2676 20640 2692 20704
rect 2756 20640 2772 20704
rect 2836 20640 2852 20704
rect 2916 20640 2924 20704
rect 2604 19616 2924 20640
rect 2604 19552 2612 19616
rect 2676 19552 2692 19616
rect 2756 19552 2772 19616
rect 2836 19552 2852 19616
rect 2916 19552 2924 19616
rect 2604 18954 2924 19552
rect 2604 18718 2646 18954
rect 2882 18718 2924 18954
rect 2604 18528 2924 18718
rect 2604 18464 2612 18528
rect 2676 18464 2692 18528
rect 2756 18464 2772 18528
rect 2836 18464 2852 18528
rect 2916 18464 2924 18528
rect 2604 17440 2924 18464
rect 2604 17376 2612 17440
rect 2676 17376 2692 17440
rect 2756 17376 2772 17440
rect 2836 17376 2852 17440
rect 2916 17376 2924 17440
rect 2604 16352 2924 17376
rect 2604 16288 2612 16352
rect 2676 16288 2692 16352
rect 2756 16288 2772 16352
rect 2836 16288 2852 16352
rect 2916 16288 2924 16352
rect 2604 15264 2924 16288
rect 2604 15200 2612 15264
rect 2676 15200 2692 15264
rect 2756 15200 2772 15264
rect 2836 15200 2852 15264
rect 2916 15200 2924 15264
rect 2604 14176 2924 15200
rect 2604 14112 2612 14176
rect 2676 14112 2692 14176
rect 2756 14112 2772 14176
rect 2836 14112 2852 14176
rect 2916 14112 2924 14176
rect 2604 13954 2924 14112
rect 2604 13718 2646 13954
rect 2882 13718 2924 13954
rect 2604 13088 2924 13718
rect 2604 13024 2612 13088
rect 2676 13024 2692 13088
rect 2756 13024 2772 13088
rect 2836 13024 2852 13088
rect 2916 13024 2924 13088
rect 2604 12000 2924 13024
rect 2604 11936 2612 12000
rect 2676 11936 2692 12000
rect 2756 11936 2772 12000
rect 2836 11936 2852 12000
rect 2916 11936 2924 12000
rect 2604 10912 2924 11936
rect 3374 11117 3434 67627
rect 6944 66944 7264 67968
rect 6944 66880 6952 66944
rect 7016 66880 7032 66944
rect 7096 66880 7112 66944
rect 7176 66880 7192 66944
rect 7256 66880 7264 66944
rect 6944 65856 7264 66880
rect 6944 65792 6952 65856
rect 7016 65792 7032 65856
rect 7096 65792 7112 65856
rect 7176 65792 7192 65856
rect 7256 65792 7264 65856
rect 6944 64768 7264 65792
rect 6944 64704 6952 64768
rect 7016 64704 7032 64768
rect 7096 64704 7112 64768
rect 7176 64704 7192 64768
rect 7256 64704 7264 64768
rect 6944 63680 7264 64704
rect 6944 63616 6952 63680
rect 7016 63616 7032 63680
rect 7096 63616 7112 63680
rect 7176 63616 7192 63680
rect 7256 63616 7264 63680
rect 6944 63294 7264 63616
rect 6944 63058 6986 63294
rect 7222 63058 7264 63294
rect 6944 62592 7264 63058
rect 6944 62528 6952 62592
rect 7016 62528 7032 62592
rect 7096 62528 7112 62592
rect 7176 62528 7192 62592
rect 7256 62528 7264 62592
rect 6944 61504 7264 62528
rect 6944 61440 6952 61504
rect 7016 61440 7032 61504
rect 7096 61440 7112 61504
rect 7176 61440 7192 61504
rect 7256 61440 7264 61504
rect 6944 60416 7264 61440
rect 6944 60352 6952 60416
rect 7016 60352 7032 60416
rect 7096 60352 7112 60416
rect 7176 60352 7192 60416
rect 7256 60352 7264 60416
rect 6944 59328 7264 60352
rect 6944 59264 6952 59328
rect 7016 59264 7032 59328
rect 7096 59264 7112 59328
rect 7176 59264 7192 59328
rect 7256 59264 7264 59328
rect 6944 58294 7264 59264
rect 6944 58240 6986 58294
rect 7222 58240 7264 58294
rect 6944 58176 6952 58240
rect 7256 58176 7264 58240
rect 6944 58058 6986 58176
rect 7222 58058 7264 58176
rect 6944 57152 7264 58058
rect 6944 57088 6952 57152
rect 7016 57088 7032 57152
rect 7096 57088 7112 57152
rect 7176 57088 7192 57152
rect 7256 57088 7264 57152
rect 6944 56064 7264 57088
rect 6944 56000 6952 56064
rect 7016 56000 7032 56064
rect 7096 56000 7112 56064
rect 7176 56000 7192 56064
rect 7256 56000 7264 56064
rect 6944 54976 7264 56000
rect 6944 54912 6952 54976
rect 7016 54912 7032 54976
rect 7096 54912 7112 54976
rect 7176 54912 7192 54976
rect 7256 54912 7264 54976
rect 6944 53888 7264 54912
rect 6944 53824 6952 53888
rect 7016 53824 7032 53888
rect 7096 53824 7112 53888
rect 7176 53824 7192 53888
rect 7256 53824 7264 53888
rect 6944 53294 7264 53824
rect 6944 53058 6986 53294
rect 7222 53058 7264 53294
rect 6944 52800 7264 53058
rect 6944 52736 6952 52800
rect 7016 52736 7032 52800
rect 7096 52736 7112 52800
rect 7176 52736 7192 52800
rect 7256 52736 7264 52800
rect 6944 51712 7264 52736
rect 6944 51648 6952 51712
rect 7016 51648 7032 51712
rect 7096 51648 7112 51712
rect 7176 51648 7192 51712
rect 7256 51648 7264 51712
rect 6944 50624 7264 51648
rect 6944 50560 6952 50624
rect 7016 50560 7032 50624
rect 7096 50560 7112 50624
rect 7176 50560 7192 50624
rect 7256 50560 7264 50624
rect 6944 49536 7264 50560
rect 6944 49472 6952 49536
rect 7016 49472 7032 49536
rect 7096 49472 7112 49536
rect 7176 49472 7192 49536
rect 7256 49472 7264 49536
rect 6944 48448 7264 49472
rect 6944 48384 6952 48448
rect 7016 48384 7032 48448
rect 7096 48384 7112 48448
rect 7176 48384 7192 48448
rect 7256 48384 7264 48448
rect 6944 48294 7264 48384
rect 6944 48058 6986 48294
rect 7222 48058 7264 48294
rect 6944 47360 7264 48058
rect 6944 47296 6952 47360
rect 7016 47296 7032 47360
rect 7096 47296 7112 47360
rect 7176 47296 7192 47360
rect 7256 47296 7264 47360
rect 6944 46272 7264 47296
rect 6944 46208 6952 46272
rect 7016 46208 7032 46272
rect 7096 46208 7112 46272
rect 7176 46208 7192 46272
rect 7256 46208 7264 46272
rect 6944 45184 7264 46208
rect 6944 45120 6952 45184
rect 7016 45120 7032 45184
rect 7096 45120 7112 45184
rect 7176 45120 7192 45184
rect 7256 45120 7264 45184
rect 6944 44096 7264 45120
rect 6944 44032 6952 44096
rect 7016 44032 7032 44096
rect 7096 44032 7112 44096
rect 7176 44032 7192 44096
rect 7256 44032 7264 44096
rect 6944 43294 7264 44032
rect 6944 43058 6986 43294
rect 7222 43058 7264 43294
rect 6944 43008 7264 43058
rect 6944 42944 6952 43008
rect 7016 42944 7032 43008
rect 7096 42944 7112 43008
rect 7176 42944 7192 43008
rect 7256 42944 7264 43008
rect 6944 41920 7264 42944
rect 6944 41856 6952 41920
rect 7016 41856 7032 41920
rect 7096 41856 7112 41920
rect 7176 41856 7192 41920
rect 7256 41856 7264 41920
rect 6944 40832 7264 41856
rect 6944 40768 6952 40832
rect 7016 40768 7032 40832
rect 7096 40768 7112 40832
rect 7176 40768 7192 40832
rect 7256 40768 7264 40832
rect 6944 39744 7264 40768
rect 6944 39680 6952 39744
rect 7016 39680 7032 39744
rect 7096 39680 7112 39744
rect 7176 39680 7192 39744
rect 7256 39680 7264 39744
rect 6944 38656 7264 39680
rect 6944 38592 6952 38656
rect 7016 38592 7032 38656
rect 7096 38592 7112 38656
rect 7176 38592 7192 38656
rect 7256 38592 7264 38656
rect 6944 38294 7264 38592
rect 6944 38058 6986 38294
rect 7222 38058 7264 38294
rect 6944 37568 7264 38058
rect 6944 37504 6952 37568
rect 7016 37504 7032 37568
rect 7096 37504 7112 37568
rect 7176 37504 7192 37568
rect 7256 37504 7264 37568
rect 6944 36480 7264 37504
rect 6944 36416 6952 36480
rect 7016 36416 7032 36480
rect 7096 36416 7112 36480
rect 7176 36416 7192 36480
rect 7256 36416 7264 36480
rect 6944 35392 7264 36416
rect 6944 35328 6952 35392
rect 7016 35328 7032 35392
rect 7096 35328 7112 35392
rect 7176 35328 7192 35392
rect 7256 35328 7264 35392
rect 6944 34304 7264 35328
rect 6944 34240 6952 34304
rect 7016 34240 7032 34304
rect 7096 34240 7112 34304
rect 7176 34240 7192 34304
rect 7256 34240 7264 34304
rect 6944 33294 7264 34240
rect 6944 33216 6986 33294
rect 7222 33216 7264 33294
rect 6944 33152 6952 33216
rect 7256 33152 7264 33216
rect 6944 33058 6986 33152
rect 7222 33058 7264 33152
rect 6944 32128 7264 33058
rect 6944 32064 6952 32128
rect 7016 32064 7032 32128
rect 7096 32064 7112 32128
rect 7176 32064 7192 32128
rect 7256 32064 7264 32128
rect 6944 31040 7264 32064
rect 6944 30976 6952 31040
rect 7016 30976 7032 31040
rect 7096 30976 7112 31040
rect 7176 30976 7192 31040
rect 7256 30976 7264 31040
rect 6944 29952 7264 30976
rect 6944 29888 6952 29952
rect 7016 29888 7032 29952
rect 7096 29888 7112 29952
rect 7176 29888 7192 29952
rect 7256 29888 7264 29952
rect 6944 28864 7264 29888
rect 6944 28800 6952 28864
rect 7016 28800 7032 28864
rect 7096 28800 7112 28864
rect 7176 28800 7192 28864
rect 7256 28800 7264 28864
rect 6944 28294 7264 28800
rect 6944 28058 6986 28294
rect 7222 28058 7264 28294
rect 6944 27776 7264 28058
rect 6944 27712 6952 27776
rect 7016 27712 7032 27776
rect 7096 27712 7112 27776
rect 7176 27712 7192 27776
rect 7256 27712 7264 27776
rect 6944 26688 7264 27712
rect 6944 26624 6952 26688
rect 7016 26624 7032 26688
rect 7096 26624 7112 26688
rect 7176 26624 7192 26688
rect 7256 26624 7264 26688
rect 6944 25600 7264 26624
rect 6944 25536 6952 25600
rect 7016 25536 7032 25600
rect 7096 25536 7112 25600
rect 7176 25536 7192 25600
rect 7256 25536 7264 25600
rect 6944 24512 7264 25536
rect 6944 24448 6952 24512
rect 7016 24448 7032 24512
rect 7096 24448 7112 24512
rect 7176 24448 7192 24512
rect 7256 24448 7264 24512
rect 6944 23424 7264 24448
rect 6944 23360 6952 23424
rect 7016 23360 7032 23424
rect 7096 23360 7112 23424
rect 7176 23360 7192 23424
rect 7256 23360 7264 23424
rect 6944 23294 7264 23360
rect 6944 23058 6986 23294
rect 7222 23058 7264 23294
rect 6944 22336 7264 23058
rect 6944 22272 6952 22336
rect 7016 22272 7032 22336
rect 7096 22272 7112 22336
rect 7176 22272 7192 22336
rect 7256 22272 7264 22336
rect 6944 21248 7264 22272
rect 6944 21184 6952 21248
rect 7016 21184 7032 21248
rect 7096 21184 7112 21248
rect 7176 21184 7192 21248
rect 7256 21184 7264 21248
rect 6944 20160 7264 21184
rect 6944 20096 6952 20160
rect 7016 20096 7032 20160
rect 7096 20096 7112 20160
rect 7176 20096 7192 20160
rect 7256 20096 7264 20160
rect 6944 19072 7264 20096
rect 6944 19008 6952 19072
rect 7016 19008 7032 19072
rect 7096 19008 7112 19072
rect 7176 19008 7192 19072
rect 7256 19008 7264 19072
rect 6944 18294 7264 19008
rect 6944 18058 6986 18294
rect 7222 18058 7264 18294
rect 6944 17984 7264 18058
rect 6944 17920 6952 17984
rect 7016 17920 7032 17984
rect 7096 17920 7112 17984
rect 7176 17920 7192 17984
rect 7256 17920 7264 17984
rect 6944 16896 7264 17920
rect 6944 16832 6952 16896
rect 7016 16832 7032 16896
rect 7096 16832 7112 16896
rect 7176 16832 7192 16896
rect 7256 16832 7264 16896
rect 6944 15808 7264 16832
rect 6944 15744 6952 15808
rect 7016 15744 7032 15808
rect 7096 15744 7112 15808
rect 7176 15744 7192 15808
rect 7256 15744 7264 15808
rect 6944 14720 7264 15744
rect 6944 14656 6952 14720
rect 7016 14656 7032 14720
rect 7096 14656 7112 14720
rect 7176 14656 7192 14720
rect 7256 14656 7264 14720
rect 6944 13632 7264 14656
rect 6944 13568 6952 13632
rect 7016 13568 7032 13632
rect 7096 13568 7112 13632
rect 7176 13568 7192 13632
rect 7256 13568 7264 13632
rect 6944 13294 7264 13568
rect 6944 13058 6986 13294
rect 7222 13058 7264 13294
rect 6944 12544 7264 13058
rect 6944 12480 6952 12544
rect 7016 12480 7032 12544
rect 7096 12480 7112 12544
rect 7176 12480 7192 12544
rect 7256 12480 7264 12544
rect 6944 11456 7264 12480
rect 6944 11392 6952 11456
rect 7016 11392 7032 11456
rect 7096 11392 7112 11456
rect 7176 11392 7192 11456
rect 7256 11392 7264 11456
rect 3371 11116 3437 11117
rect 3371 11052 3372 11116
rect 3436 11052 3437 11116
rect 3371 11051 3437 11052
rect 2604 10848 2612 10912
rect 2676 10848 2692 10912
rect 2756 10848 2772 10912
rect 2836 10848 2852 10912
rect 2916 10848 2924 10912
rect 2604 9824 2924 10848
rect 2604 9760 2612 9824
rect 2676 9760 2692 9824
rect 2756 9760 2772 9824
rect 2836 9760 2852 9824
rect 2916 9760 2924 9824
rect 2604 8954 2924 9760
rect 2604 8736 2646 8954
rect 2882 8736 2924 8954
rect 2604 8672 2612 8736
rect 2676 8672 2692 8718
rect 2756 8672 2772 8718
rect 2836 8672 2852 8718
rect 2916 8672 2924 8736
rect 2604 7648 2924 8672
rect 2604 7584 2612 7648
rect 2676 7584 2692 7648
rect 2756 7584 2772 7648
rect 2836 7584 2852 7648
rect 2916 7584 2924 7648
rect 2604 6560 2924 7584
rect 2604 6496 2612 6560
rect 2676 6496 2692 6560
rect 2756 6496 2772 6560
rect 2836 6496 2852 6560
rect 2916 6496 2924 6560
rect 2604 5472 2924 6496
rect 2604 5408 2612 5472
rect 2676 5408 2692 5472
rect 2756 5408 2772 5472
rect 2836 5408 2852 5472
rect 2916 5408 2924 5472
rect 2604 4384 2924 5408
rect 2604 4320 2612 4384
rect 2676 4320 2692 4384
rect 2756 4320 2772 4384
rect 2836 4320 2852 4384
rect 2916 4320 2924 4384
rect 2604 3954 2924 4320
rect 2604 3718 2646 3954
rect 2882 3718 2924 3954
rect 2604 3296 2924 3718
rect 2604 3232 2612 3296
rect 2676 3232 2692 3296
rect 2756 3232 2772 3296
rect 2836 3232 2852 3296
rect 2916 3232 2924 3296
rect 2604 2208 2924 3232
rect 2604 2144 2612 2208
rect 2676 2144 2692 2208
rect 2756 2144 2772 2208
rect 2836 2144 2852 2208
rect 2916 2144 2924 2208
rect 2604 2128 2924 2144
rect 6944 10368 7264 11392
rect 6944 10304 6952 10368
rect 7016 10304 7032 10368
rect 7096 10304 7112 10368
rect 7176 10304 7192 10368
rect 7256 10304 7264 10368
rect 6944 9280 7264 10304
rect 6944 9216 6952 9280
rect 7016 9216 7032 9280
rect 7096 9216 7112 9280
rect 7176 9216 7192 9280
rect 7256 9216 7264 9280
rect 6944 8294 7264 9216
rect 6944 8192 6986 8294
rect 7222 8192 7264 8294
rect 6944 8128 6952 8192
rect 7256 8128 7264 8192
rect 6944 8058 6986 8128
rect 7222 8058 7264 8128
rect 6944 7104 7264 8058
rect 6944 7040 6952 7104
rect 7016 7040 7032 7104
rect 7096 7040 7112 7104
rect 7176 7040 7192 7104
rect 7256 7040 7264 7104
rect 6944 6016 7264 7040
rect 6944 5952 6952 6016
rect 7016 5952 7032 6016
rect 7096 5952 7112 6016
rect 7176 5952 7192 6016
rect 7256 5952 7264 6016
rect 6944 4928 7264 5952
rect 6944 4864 6952 4928
rect 7016 4864 7032 4928
rect 7096 4864 7112 4928
rect 7176 4864 7192 4928
rect 7256 4864 7264 4928
rect 6944 3840 7264 4864
rect 6944 3776 6952 3840
rect 7016 3776 7032 3840
rect 7096 3776 7112 3840
rect 7176 3776 7192 3840
rect 7256 3776 7264 3840
rect 6944 3294 7264 3776
rect 6944 3058 6986 3294
rect 7222 3058 7264 3294
rect 6944 2752 7264 3058
rect 6944 2688 6952 2752
rect 7016 2688 7032 2752
rect 7096 2688 7112 2752
rect 7176 2688 7192 2752
rect 7256 2688 7264 2752
rect 6944 2128 7264 2688
rect 7604 69664 7924 69680
rect 7604 69600 7612 69664
rect 7676 69600 7692 69664
rect 7756 69600 7772 69664
rect 7836 69600 7852 69664
rect 7916 69600 7924 69664
rect 7604 68954 7924 69600
rect 7604 68718 7646 68954
rect 7882 68718 7924 68954
rect 7604 68576 7924 68718
rect 7604 68512 7612 68576
rect 7676 68512 7692 68576
rect 7756 68512 7772 68576
rect 7836 68512 7852 68576
rect 7916 68512 7924 68576
rect 7604 67488 7924 68512
rect 7604 67424 7612 67488
rect 7676 67424 7692 67488
rect 7756 67424 7772 67488
rect 7836 67424 7852 67488
rect 7916 67424 7924 67488
rect 7604 66400 7924 67424
rect 7604 66336 7612 66400
rect 7676 66336 7692 66400
rect 7756 66336 7772 66400
rect 7836 66336 7852 66400
rect 7916 66336 7924 66400
rect 7604 65312 7924 66336
rect 7604 65248 7612 65312
rect 7676 65248 7692 65312
rect 7756 65248 7772 65312
rect 7836 65248 7852 65312
rect 7916 65248 7924 65312
rect 7604 64224 7924 65248
rect 7604 64160 7612 64224
rect 7676 64160 7692 64224
rect 7756 64160 7772 64224
rect 7836 64160 7852 64224
rect 7916 64160 7924 64224
rect 7604 63954 7924 64160
rect 7604 63718 7646 63954
rect 7882 63718 7924 63954
rect 7604 63136 7924 63718
rect 7604 63072 7612 63136
rect 7676 63072 7692 63136
rect 7756 63072 7772 63136
rect 7836 63072 7852 63136
rect 7916 63072 7924 63136
rect 7604 62048 7924 63072
rect 7604 61984 7612 62048
rect 7676 61984 7692 62048
rect 7756 61984 7772 62048
rect 7836 61984 7852 62048
rect 7916 61984 7924 62048
rect 7604 60960 7924 61984
rect 7604 60896 7612 60960
rect 7676 60896 7692 60960
rect 7756 60896 7772 60960
rect 7836 60896 7852 60960
rect 7916 60896 7924 60960
rect 7604 59872 7924 60896
rect 7604 59808 7612 59872
rect 7676 59808 7692 59872
rect 7756 59808 7772 59872
rect 7836 59808 7852 59872
rect 7916 59808 7924 59872
rect 7604 58954 7924 59808
rect 7604 58784 7646 58954
rect 7882 58784 7924 58954
rect 7604 58720 7612 58784
rect 7916 58720 7924 58784
rect 7604 58718 7646 58720
rect 7882 58718 7924 58720
rect 7604 57696 7924 58718
rect 7604 57632 7612 57696
rect 7676 57632 7692 57696
rect 7756 57632 7772 57696
rect 7836 57632 7852 57696
rect 7916 57632 7924 57696
rect 7604 56608 7924 57632
rect 7604 56544 7612 56608
rect 7676 56544 7692 56608
rect 7756 56544 7772 56608
rect 7836 56544 7852 56608
rect 7916 56544 7924 56608
rect 7604 55520 7924 56544
rect 7604 55456 7612 55520
rect 7676 55456 7692 55520
rect 7756 55456 7772 55520
rect 7836 55456 7852 55520
rect 7916 55456 7924 55520
rect 7604 54432 7924 55456
rect 7604 54368 7612 54432
rect 7676 54368 7692 54432
rect 7756 54368 7772 54432
rect 7836 54368 7852 54432
rect 7916 54368 7924 54432
rect 7604 53954 7924 54368
rect 7604 53718 7646 53954
rect 7882 53718 7924 53954
rect 7604 53344 7924 53718
rect 7604 53280 7612 53344
rect 7676 53280 7692 53344
rect 7756 53280 7772 53344
rect 7836 53280 7852 53344
rect 7916 53280 7924 53344
rect 7604 52256 7924 53280
rect 7604 52192 7612 52256
rect 7676 52192 7692 52256
rect 7756 52192 7772 52256
rect 7836 52192 7852 52256
rect 7916 52192 7924 52256
rect 7604 51168 7924 52192
rect 7604 51104 7612 51168
rect 7676 51104 7692 51168
rect 7756 51104 7772 51168
rect 7836 51104 7852 51168
rect 7916 51104 7924 51168
rect 7604 50080 7924 51104
rect 7604 50016 7612 50080
rect 7676 50016 7692 50080
rect 7756 50016 7772 50080
rect 7836 50016 7852 50080
rect 7916 50016 7924 50080
rect 7604 48992 7924 50016
rect 7604 48928 7612 48992
rect 7676 48954 7692 48992
rect 7756 48954 7772 48992
rect 7836 48954 7852 48992
rect 7916 48928 7924 48992
rect 7604 48718 7646 48928
rect 7882 48718 7924 48928
rect 7604 47904 7924 48718
rect 7604 47840 7612 47904
rect 7676 47840 7692 47904
rect 7756 47840 7772 47904
rect 7836 47840 7852 47904
rect 7916 47840 7924 47904
rect 7604 46816 7924 47840
rect 7604 46752 7612 46816
rect 7676 46752 7692 46816
rect 7756 46752 7772 46816
rect 7836 46752 7852 46816
rect 7916 46752 7924 46816
rect 7604 45728 7924 46752
rect 7604 45664 7612 45728
rect 7676 45664 7692 45728
rect 7756 45664 7772 45728
rect 7836 45664 7852 45728
rect 7916 45664 7924 45728
rect 7604 44640 7924 45664
rect 7604 44576 7612 44640
rect 7676 44576 7692 44640
rect 7756 44576 7772 44640
rect 7836 44576 7852 44640
rect 7916 44576 7924 44640
rect 7604 43954 7924 44576
rect 7604 43718 7646 43954
rect 7882 43718 7924 43954
rect 7604 43552 7924 43718
rect 7604 43488 7612 43552
rect 7676 43488 7692 43552
rect 7756 43488 7772 43552
rect 7836 43488 7852 43552
rect 7916 43488 7924 43552
rect 7604 42464 7924 43488
rect 7604 42400 7612 42464
rect 7676 42400 7692 42464
rect 7756 42400 7772 42464
rect 7836 42400 7852 42464
rect 7916 42400 7924 42464
rect 7604 41376 7924 42400
rect 7604 41312 7612 41376
rect 7676 41312 7692 41376
rect 7756 41312 7772 41376
rect 7836 41312 7852 41376
rect 7916 41312 7924 41376
rect 7604 40288 7924 41312
rect 7604 40224 7612 40288
rect 7676 40224 7692 40288
rect 7756 40224 7772 40288
rect 7836 40224 7852 40288
rect 7916 40224 7924 40288
rect 7604 39200 7924 40224
rect 7604 39136 7612 39200
rect 7676 39136 7692 39200
rect 7756 39136 7772 39200
rect 7836 39136 7852 39200
rect 7916 39136 7924 39200
rect 7604 38954 7924 39136
rect 7604 38718 7646 38954
rect 7882 38718 7924 38954
rect 7604 38112 7924 38718
rect 7604 38048 7612 38112
rect 7676 38048 7692 38112
rect 7756 38048 7772 38112
rect 7836 38048 7852 38112
rect 7916 38048 7924 38112
rect 7604 37024 7924 38048
rect 7604 36960 7612 37024
rect 7676 36960 7692 37024
rect 7756 36960 7772 37024
rect 7836 36960 7852 37024
rect 7916 36960 7924 37024
rect 7604 35936 7924 36960
rect 7604 35872 7612 35936
rect 7676 35872 7692 35936
rect 7756 35872 7772 35936
rect 7836 35872 7852 35936
rect 7916 35872 7924 35936
rect 7604 34848 7924 35872
rect 7604 34784 7612 34848
rect 7676 34784 7692 34848
rect 7756 34784 7772 34848
rect 7836 34784 7852 34848
rect 7916 34784 7924 34848
rect 7604 33954 7924 34784
rect 7604 33760 7646 33954
rect 7882 33760 7924 33954
rect 7604 33696 7612 33760
rect 7676 33696 7692 33718
rect 7756 33696 7772 33718
rect 7836 33696 7852 33718
rect 7916 33696 7924 33760
rect 7604 32672 7924 33696
rect 7604 32608 7612 32672
rect 7676 32608 7692 32672
rect 7756 32608 7772 32672
rect 7836 32608 7852 32672
rect 7916 32608 7924 32672
rect 7604 31584 7924 32608
rect 7604 31520 7612 31584
rect 7676 31520 7692 31584
rect 7756 31520 7772 31584
rect 7836 31520 7852 31584
rect 7916 31520 7924 31584
rect 7604 30496 7924 31520
rect 7604 30432 7612 30496
rect 7676 30432 7692 30496
rect 7756 30432 7772 30496
rect 7836 30432 7852 30496
rect 7916 30432 7924 30496
rect 7604 29408 7924 30432
rect 7604 29344 7612 29408
rect 7676 29344 7692 29408
rect 7756 29344 7772 29408
rect 7836 29344 7852 29408
rect 7916 29344 7924 29408
rect 7604 28954 7924 29344
rect 7604 28718 7646 28954
rect 7882 28718 7924 28954
rect 7604 28320 7924 28718
rect 7604 28256 7612 28320
rect 7676 28256 7692 28320
rect 7756 28256 7772 28320
rect 7836 28256 7852 28320
rect 7916 28256 7924 28320
rect 7604 27232 7924 28256
rect 7604 27168 7612 27232
rect 7676 27168 7692 27232
rect 7756 27168 7772 27232
rect 7836 27168 7852 27232
rect 7916 27168 7924 27232
rect 7604 26144 7924 27168
rect 7604 26080 7612 26144
rect 7676 26080 7692 26144
rect 7756 26080 7772 26144
rect 7836 26080 7852 26144
rect 7916 26080 7924 26144
rect 7604 25056 7924 26080
rect 7604 24992 7612 25056
rect 7676 24992 7692 25056
rect 7756 24992 7772 25056
rect 7836 24992 7852 25056
rect 7916 24992 7924 25056
rect 7604 23968 7924 24992
rect 7604 23904 7612 23968
rect 7676 23954 7692 23968
rect 7756 23954 7772 23968
rect 7836 23954 7852 23968
rect 7916 23904 7924 23968
rect 7604 23718 7646 23904
rect 7882 23718 7924 23904
rect 7604 22880 7924 23718
rect 7604 22816 7612 22880
rect 7676 22816 7692 22880
rect 7756 22816 7772 22880
rect 7836 22816 7852 22880
rect 7916 22816 7924 22880
rect 7604 21792 7924 22816
rect 7604 21728 7612 21792
rect 7676 21728 7692 21792
rect 7756 21728 7772 21792
rect 7836 21728 7852 21792
rect 7916 21728 7924 21792
rect 7604 20704 7924 21728
rect 7604 20640 7612 20704
rect 7676 20640 7692 20704
rect 7756 20640 7772 20704
rect 7836 20640 7852 20704
rect 7916 20640 7924 20704
rect 7604 19616 7924 20640
rect 7604 19552 7612 19616
rect 7676 19552 7692 19616
rect 7756 19552 7772 19616
rect 7836 19552 7852 19616
rect 7916 19552 7924 19616
rect 7604 18954 7924 19552
rect 7604 18718 7646 18954
rect 7882 18718 7924 18954
rect 7604 18528 7924 18718
rect 7604 18464 7612 18528
rect 7676 18464 7692 18528
rect 7756 18464 7772 18528
rect 7836 18464 7852 18528
rect 7916 18464 7924 18528
rect 7604 17440 7924 18464
rect 7604 17376 7612 17440
rect 7676 17376 7692 17440
rect 7756 17376 7772 17440
rect 7836 17376 7852 17440
rect 7916 17376 7924 17440
rect 7604 16352 7924 17376
rect 7604 16288 7612 16352
rect 7676 16288 7692 16352
rect 7756 16288 7772 16352
rect 7836 16288 7852 16352
rect 7916 16288 7924 16352
rect 7604 15264 7924 16288
rect 7604 15200 7612 15264
rect 7676 15200 7692 15264
rect 7756 15200 7772 15264
rect 7836 15200 7852 15264
rect 7916 15200 7924 15264
rect 7604 14176 7924 15200
rect 7604 14112 7612 14176
rect 7676 14112 7692 14176
rect 7756 14112 7772 14176
rect 7836 14112 7852 14176
rect 7916 14112 7924 14176
rect 7604 13954 7924 14112
rect 7604 13718 7646 13954
rect 7882 13718 7924 13954
rect 7604 13088 7924 13718
rect 7604 13024 7612 13088
rect 7676 13024 7692 13088
rect 7756 13024 7772 13088
rect 7836 13024 7852 13088
rect 7916 13024 7924 13088
rect 7604 12000 7924 13024
rect 7604 11936 7612 12000
rect 7676 11936 7692 12000
rect 7756 11936 7772 12000
rect 7836 11936 7852 12000
rect 7916 11936 7924 12000
rect 7604 10912 7924 11936
rect 7604 10848 7612 10912
rect 7676 10848 7692 10912
rect 7756 10848 7772 10912
rect 7836 10848 7852 10912
rect 7916 10848 7924 10912
rect 7604 9824 7924 10848
rect 7604 9760 7612 9824
rect 7676 9760 7692 9824
rect 7756 9760 7772 9824
rect 7836 9760 7852 9824
rect 7916 9760 7924 9824
rect 7604 8954 7924 9760
rect 7604 8736 7646 8954
rect 7882 8736 7924 8954
rect 7604 8672 7612 8736
rect 7676 8672 7692 8718
rect 7756 8672 7772 8718
rect 7836 8672 7852 8718
rect 7916 8672 7924 8736
rect 7604 7648 7924 8672
rect 7604 7584 7612 7648
rect 7676 7584 7692 7648
rect 7756 7584 7772 7648
rect 7836 7584 7852 7648
rect 7916 7584 7924 7648
rect 7604 6560 7924 7584
rect 7604 6496 7612 6560
rect 7676 6496 7692 6560
rect 7756 6496 7772 6560
rect 7836 6496 7852 6560
rect 7916 6496 7924 6560
rect 7604 5472 7924 6496
rect 7604 5408 7612 5472
rect 7676 5408 7692 5472
rect 7756 5408 7772 5472
rect 7836 5408 7852 5472
rect 7916 5408 7924 5472
rect 7604 4384 7924 5408
rect 7604 4320 7612 4384
rect 7676 4320 7692 4384
rect 7756 4320 7772 4384
rect 7836 4320 7852 4384
rect 7916 4320 7924 4384
rect 7604 3954 7924 4320
rect 7604 3718 7646 3954
rect 7882 3718 7924 3954
rect 7604 3296 7924 3718
rect 7604 3232 7612 3296
rect 7676 3232 7692 3296
rect 7756 3232 7772 3296
rect 7836 3232 7852 3296
rect 7916 3232 7924 3296
rect 7604 2208 7924 3232
rect 7604 2144 7612 2208
rect 7676 2144 7692 2208
rect 7756 2144 7772 2208
rect 7836 2144 7852 2208
rect 7916 2144 7924 2208
rect 7604 2128 7924 2144
rect 11944 69120 12264 69680
rect 11944 69056 11952 69120
rect 12016 69056 12032 69120
rect 12096 69056 12112 69120
rect 12176 69056 12192 69120
rect 12256 69056 12264 69120
rect 11944 68294 12264 69056
rect 11944 68058 11986 68294
rect 12222 68058 12264 68294
rect 11944 68032 12264 68058
rect 11944 67968 11952 68032
rect 12016 67968 12032 68032
rect 12096 67968 12112 68032
rect 12176 67968 12192 68032
rect 12256 67968 12264 68032
rect 11944 66944 12264 67968
rect 11944 66880 11952 66944
rect 12016 66880 12032 66944
rect 12096 66880 12112 66944
rect 12176 66880 12192 66944
rect 12256 66880 12264 66944
rect 11944 65856 12264 66880
rect 11944 65792 11952 65856
rect 12016 65792 12032 65856
rect 12096 65792 12112 65856
rect 12176 65792 12192 65856
rect 12256 65792 12264 65856
rect 11944 64768 12264 65792
rect 11944 64704 11952 64768
rect 12016 64704 12032 64768
rect 12096 64704 12112 64768
rect 12176 64704 12192 64768
rect 12256 64704 12264 64768
rect 11944 63680 12264 64704
rect 11944 63616 11952 63680
rect 12016 63616 12032 63680
rect 12096 63616 12112 63680
rect 12176 63616 12192 63680
rect 12256 63616 12264 63680
rect 11944 63294 12264 63616
rect 11944 63058 11986 63294
rect 12222 63058 12264 63294
rect 11944 62592 12264 63058
rect 11944 62528 11952 62592
rect 12016 62528 12032 62592
rect 12096 62528 12112 62592
rect 12176 62528 12192 62592
rect 12256 62528 12264 62592
rect 11944 61504 12264 62528
rect 11944 61440 11952 61504
rect 12016 61440 12032 61504
rect 12096 61440 12112 61504
rect 12176 61440 12192 61504
rect 12256 61440 12264 61504
rect 11944 60416 12264 61440
rect 11944 60352 11952 60416
rect 12016 60352 12032 60416
rect 12096 60352 12112 60416
rect 12176 60352 12192 60416
rect 12256 60352 12264 60416
rect 11944 59328 12264 60352
rect 11944 59264 11952 59328
rect 12016 59264 12032 59328
rect 12096 59264 12112 59328
rect 12176 59264 12192 59328
rect 12256 59264 12264 59328
rect 11944 58294 12264 59264
rect 11944 58240 11986 58294
rect 12222 58240 12264 58294
rect 11944 58176 11952 58240
rect 12256 58176 12264 58240
rect 11944 58058 11986 58176
rect 12222 58058 12264 58176
rect 11944 57152 12264 58058
rect 11944 57088 11952 57152
rect 12016 57088 12032 57152
rect 12096 57088 12112 57152
rect 12176 57088 12192 57152
rect 12256 57088 12264 57152
rect 11944 56064 12264 57088
rect 11944 56000 11952 56064
rect 12016 56000 12032 56064
rect 12096 56000 12112 56064
rect 12176 56000 12192 56064
rect 12256 56000 12264 56064
rect 11944 54976 12264 56000
rect 11944 54912 11952 54976
rect 12016 54912 12032 54976
rect 12096 54912 12112 54976
rect 12176 54912 12192 54976
rect 12256 54912 12264 54976
rect 11944 53888 12264 54912
rect 11944 53824 11952 53888
rect 12016 53824 12032 53888
rect 12096 53824 12112 53888
rect 12176 53824 12192 53888
rect 12256 53824 12264 53888
rect 11944 53294 12264 53824
rect 11944 53058 11986 53294
rect 12222 53058 12264 53294
rect 11944 52800 12264 53058
rect 11944 52736 11952 52800
rect 12016 52736 12032 52800
rect 12096 52736 12112 52800
rect 12176 52736 12192 52800
rect 12256 52736 12264 52800
rect 11944 51712 12264 52736
rect 11944 51648 11952 51712
rect 12016 51648 12032 51712
rect 12096 51648 12112 51712
rect 12176 51648 12192 51712
rect 12256 51648 12264 51712
rect 11944 50624 12264 51648
rect 11944 50560 11952 50624
rect 12016 50560 12032 50624
rect 12096 50560 12112 50624
rect 12176 50560 12192 50624
rect 12256 50560 12264 50624
rect 11944 49536 12264 50560
rect 11944 49472 11952 49536
rect 12016 49472 12032 49536
rect 12096 49472 12112 49536
rect 12176 49472 12192 49536
rect 12256 49472 12264 49536
rect 11944 48448 12264 49472
rect 11944 48384 11952 48448
rect 12016 48384 12032 48448
rect 12096 48384 12112 48448
rect 12176 48384 12192 48448
rect 12256 48384 12264 48448
rect 11944 48294 12264 48384
rect 11944 48058 11986 48294
rect 12222 48058 12264 48294
rect 11944 47360 12264 48058
rect 11944 47296 11952 47360
rect 12016 47296 12032 47360
rect 12096 47296 12112 47360
rect 12176 47296 12192 47360
rect 12256 47296 12264 47360
rect 11944 46272 12264 47296
rect 11944 46208 11952 46272
rect 12016 46208 12032 46272
rect 12096 46208 12112 46272
rect 12176 46208 12192 46272
rect 12256 46208 12264 46272
rect 11944 45184 12264 46208
rect 11944 45120 11952 45184
rect 12016 45120 12032 45184
rect 12096 45120 12112 45184
rect 12176 45120 12192 45184
rect 12256 45120 12264 45184
rect 11944 44096 12264 45120
rect 11944 44032 11952 44096
rect 12016 44032 12032 44096
rect 12096 44032 12112 44096
rect 12176 44032 12192 44096
rect 12256 44032 12264 44096
rect 11944 43294 12264 44032
rect 11944 43058 11986 43294
rect 12222 43058 12264 43294
rect 11944 43008 12264 43058
rect 11944 42944 11952 43008
rect 12016 42944 12032 43008
rect 12096 42944 12112 43008
rect 12176 42944 12192 43008
rect 12256 42944 12264 43008
rect 11944 41920 12264 42944
rect 11944 41856 11952 41920
rect 12016 41856 12032 41920
rect 12096 41856 12112 41920
rect 12176 41856 12192 41920
rect 12256 41856 12264 41920
rect 11944 40832 12264 41856
rect 11944 40768 11952 40832
rect 12016 40768 12032 40832
rect 12096 40768 12112 40832
rect 12176 40768 12192 40832
rect 12256 40768 12264 40832
rect 11944 39744 12264 40768
rect 11944 39680 11952 39744
rect 12016 39680 12032 39744
rect 12096 39680 12112 39744
rect 12176 39680 12192 39744
rect 12256 39680 12264 39744
rect 11944 38656 12264 39680
rect 11944 38592 11952 38656
rect 12016 38592 12032 38656
rect 12096 38592 12112 38656
rect 12176 38592 12192 38656
rect 12256 38592 12264 38656
rect 11944 38294 12264 38592
rect 11944 38058 11986 38294
rect 12222 38058 12264 38294
rect 11944 37568 12264 38058
rect 11944 37504 11952 37568
rect 12016 37504 12032 37568
rect 12096 37504 12112 37568
rect 12176 37504 12192 37568
rect 12256 37504 12264 37568
rect 11944 36480 12264 37504
rect 11944 36416 11952 36480
rect 12016 36416 12032 36480
rect 12096 36416 12112 36480
rect 12176 36416 12192 36480
rect 12256 36416 12264 36480
rect 11944 35392 12264 36416
rect 11944 35328 11952 35392
rect 12016 35328 12032 35392
rect 12096 35328 12112 35392
rect 12176 35328 12192 35392
rect 12256 35328 12264 35392
rect 11944 34304 12264 35328
rect 11944 34240 11952 34304
rect 12016 34240 12032 34304
rect 12096 34240 12112 34304
rect 12176 34240 12192 34304
rect 12256 34240 12264 34304
rect 11944 33294 12264 34240
rect 11944 33216 11986 33294
rect 12222 33216 12264 33294
rect 11944 33152 11952 33216
rect 12256 33152 12264 33216
rect 11944 33058 11986 33152
rect 12222 33058 12264 33152
rect 11944 32128 12264 33058
rect 11944 32064 11952 32128
rect 12016 32064 12032 32128
rect 12096 32064 12112 32128
rect 12176 32064 12192 32128
rect 12256 32064 12264 32128
rect 11944 31040 12264 32064
rect 11944 30976 11952 31040
rect 12016 30976 12032 31040
rect 12096 30976 12112 31040
rect 12176 30976 12192 31040
rect 12256 30976 12264 31040
rect 11944 29952 12264 30976
rect 11944 29888 11952 29952
rect 12016 29888 12032 29952
rect 12096 29888 12112 29952
rect 12176 29888 12192 29952
rect 12256 29888 12264 29952
rect 11944 28864 12264 29888
rect 11944 28800 11952 28864
rect 12016 28800 12032 28864
rect 12096 28800 12112 28864
rect 12176 28800 12192 28864
rect 12256 28800 12264 28864
rect 11944 28294 12264 28800
rect 11944 28058 11986 28294
rect 12222 28058 12264 28294
rect 11944 27776 12264 28058
rect 11944 27712 11952 27776
rect 12016 27712 12032 27776
rect 12096 27712 12112 27776
rect 12176 27712 12192 27776
rect 12256 27712 12264 27776
rect 11944 26688 12264 27712
rect 11944 26624 11952 26688
rect 12016 26624 12032 26688
rect 12096 26624 12112 26688
rect 12176 26624 12192 26688
rect 12256 26624 12264 26688
rect 11944 25600 12264 26624
rect 11944 25536 11952 25600
rect 12016 25536 12032 25600
rect 12096 25536 12112 25600
rect 12176 25536 12192 25600
rect 12256 25536 12264 25600
rect 11944 24512 12264 25536
rect 11944 24448 11952 24512
rect 12016 24448 12032 24512
rect 12096 24448 12112 24512
rect 12176 24448 12192 24512
rect 12256 24448 12264 24512
rect 11944 23424 12264 24448
rect 11944 23360 11952 23424
rect 12016 23360 12032 23424
rect 12096 23360 12112 23424
rect 12176 23360 12192 23424
rect 12256 23360 12264 23424
rect 11944 23294 12264 23360
rect 11944 23058 11986 23294
rect 12222 23058 12264 23294
rect 11944 22336 12264 23058
rect 11944 22272 11952 22336
rect 12016 22272 12032 22336
rect 12096 22272 12112 22336
rect 12176 22272 12192 22336
rect 12256 22272 12264 22336
rect 11944 21248 12264 22272
rect 11944 21184 11952 21248
rect 12016 21184 12032 21248
rect 12096 21184 12112 21248
rect 12176 21184 12192 21248
rect 12256 21184 12264 21248
rect 11944 20160 12264 21184
rect 11944 20096 11952 20160
rect 12016 20096 12032 20160
rect 12096 20096 12112 20160
rect 12176 20096 12192 20160
rect 12256 20096 12264 20160
rect 11944 19072 12264 20096
rect 11944 19008 11952 19072
rect 12016 19008 12032 19072
rect 12096 19008 12112 19072
rect 12176 19008 12192 19072
rect 12256 19008 12264 19072
rect 11944 18294 12264 19008
rect 11944 18058 11986 18294
rect 12222 18058 12264 18294
rect 11944 17984 12264 18058
rect 11944 17920 11952 17984
rect 12016 17920 12032 17984
rect 12096 17920 12112 17984
rect 12176 17920 12192 17984
rect 12256 17920 12264 17984
rect 11944 16896 12264 17920
rect 11944 16832 11952 16896
rect 12016 16832 12032 16896
rect 12096 16832 12112 16896
rect 12176 16832 12192 16896
rect 12256 16832 12264 16896
rect 11944 15808 12264 16832
rect 11944 15744 11952 15808
rect 12016 15744 12032 15808
rect 12096 15744 12112 15808
rect 12176 15744 12192 15808
rect 12256 15744 12264 15808
rect 11944 14720 12264 15744
rect 11944 14656 11952 14720
rect 12016 14656 12032 14720
rect 12096 14656 12112 14720
rect 12176 14656 12192 14720
rect 12256 14656 12264 14720
rect 11944 13632 12264 14656
rect 11944 13568 11952 13632
rect 12016 13568 12032 13632
rect 12096 13568 12112 13632
rect 12176 13568 12192 13632
rect 12256 13568 12264 13632
rect 11944 13294 12264 13568
rect 11944 13058 11986 13294
rect 12222 13058 12264 13294
rect 11944 12544 12264 13058
rect 11944 12480 11952 12544
rect 12016 12480 12032 12544
rect 12096 12480 12112 12544
rect 12176 12480 12192 12544
rect 12256 12480 12264 12544
rect 11944 11456 12264 12480
rect 11944 11392 11952 11456
rect 12016 11392 12032 11456
rect 12096 11392 12112 11456
rect 12176 11392 12192 11456
rect 12256 11392 12264 11456
rect 11944 10368 12264 11392
rect 11944 10304 11952 10368
rect 12016 10304 12032 10368
rect 12096 10304 12112 10368
rect 12176 10304 12192 10368
rect 12256 10304 12264 10368
rect 11944 9280 12264 10304
rect 11944 9216 11952 9280
rect 12016 9216 12032 9280
rect 12096 9216 12112 9280
rect 12176 9216 12192 9280
rect 12256 9216 12264 9280
rect 11944 8294 12264 9216
rect 11944 8192 11986 8294
rect 12222 8192 12264 8294
rect 11944 8128 11952 8192
rect 12256 8128 12264 8192
rect 11944 8058 11986 8128
rect 12222 8058 12264 8128
rect 11944 7104 12264 8058
rect 11944 7040 11952 7104
rect 12016 7040 12032 7104
rect 12096 7040 12112 7104
rect 12176 7040 12192 7104
rect 12256 7040 12264 7104
rect 11944 6016 12264 7040
rect 11944 5952 11952 6016
rect 12016 5952 12032 6016
rect 12096 5952 12112 6016
rect 12176 5952 12192 6016
rect 12256 5952 12264 6016
rect 11944 4928 12264 5952
rect 11944 4864 11952 4928
rect 12016 4864 12032 4928
rect 12096 4864 12112 4928
rect 12176 4864 12192 4928
rect 12256 4864 12264 4928
rect 11944 3840 12264 4864
rect 11944 3776 11952 3840
rect 12016 3776 12032 3840
rect 12096 3776 12112 3840
rect 12176 3776 12192 3840
rect 12256 3776 12264 3840
rect 11944 3294 12264 3776
rect 11944 3058 11986 3294
rect 12222 3058 12264 3294
rect 11944 2752 12264 3058
rect 11944 2688 11952 2752
rect 12016 2688 12032 2752
rect 12096 2688 12112 2752
rect 12176 2688 12192 2752
rect 12256 2688 12264 2752
rect 11944 2128 12264 2688
rect 12604 69664 12924 69680
rect 12604 69600 12612 69664
rect 12676 69600 12692 69664
rect 12756 69600 12772 69664
rect 12836 69600 12852 69664
rect 12916 69600 12924 69664
rect 12604 68954 12924 69600
rect 12604 68718 12646 68954
rect 12882 68718 12924 68954
rect 12604 68576 12924 68718
rect 12604 68512 12612 68576
rect 12676 68512 12692 68576
rect 12756 68512 12772 68576
rect 12836 68512 12852 68576
rect 12916 68512 12924 68576
rect 12604 67488 12924 68512
rect 16944 69120 17264 69680
rect 16944 69056 16952 69120
rect 17016 69056 17032 69120
rect 17096 69056 17112 69120
rect 17176 69056 17192 69120
rect 17256 69056 17264 69120
rect 16944 68294 17264 69056
rect 16944 68058 16986 68294
rect 17222 68058 17264 68294
rect 16944 68032 17264 68058
rect 16944 67968 16952 68032
rect 17016 67968 17032 68032
rect 17096 67968 17112 68032
rect 17176 67968 17192 68032
rect 17256 67968 17264 68032
rect 14963 67828 15029 67829
rect 14963 67764 14964 67828
rect 15028 67764 15029 67828
rect 14963 67763 15029 67764
rect 12604 67424 12612 67488
rect 12676 67424 12692 67488
rect 12756 67424 12772 67488
rect 12836 67424 12852 67488
rect 12916 67424 12924 67488
rect 12604 66400 12924 67424
rect 12604 66336 12612 66400
rect 12676 66336 12692 66400
rect 12756 66336 12772 66400
rect 12836 66336 12852 66400
rect 12916 66336 12924 66400
rect 12604 65312 12924 66336
rect 12604 65248 12612 65312
rect 12676 65248 12692 65312
rect 12756 65248 12772 65312
rect 12836 65248 12852 65312
rect 12916 65248 12924 65312
rect 12604 64224 12924 65248
rect 12604 64160 12612 64224
rect 12676 64160 12692 64224
rect 12756 64160 12772 64224
rect 12836 64160 12852 64224
rect 12916 64160 12924 64224
rect 12604 63954 12924 64160
rect 12604 63718 12646 63954
rect 12882 63718 12924 63954
rect 12604 63136 12924 63718
rect 12604 63072 12612 63136
rect 12676 63072 12692 63136
rect 12756 63072 12772 63136
rect 12836 63072 12852 63136
rect 12916 63072 12924 63136
rect 12604 62048 12924 63072
rect 12604 61984 12612 62048
rect 12676 61984 12692 62048
rect 12756 61984 12772 62048
rect 12836 61984 12852 62048
rect 12916 61984 12924 62048
rect 12604 60960 12924 61984
rect 12604 60896 12612 60960
rect 12676 60896 12692 60960
rect 12756 60896 12772 60960
rect 12836 60896 12852 60960
rect 12916 60896 12924 60960
rect 12604 59872 12924 60896
rect 12604 59808 12612 59872
rect 12676 59808 12692 59872
rect 12756 59808 12772 59872
rect 12836 59808 12852 59872
rect 12916 59808 12924 59872
rect 12604 58954 12924 59808
rect 12604 58784 12646 58954
rect 12882 58784 12924 58954
rect 12604 58720 12612 58784
rect 12916 58720 12924 58784
rect 12604 58718 12646 58720
rect 12882 58718 12924 58720
rect 12604 57696 12924 58718
rect 12604 57632 12612 57696
rect 12676 57632 12692 57696
rect 12756 57632 12772 57696
rect 12836 57632 12852 57696
rect 12916 57632 12924 57696
rect 12604 56608 12924 57632
rect 12604 56544 12612 56608
rect 12676 56544 12692 56608
rect 12756 56544 12772 56608
rect 12836 56544 12852 56608
rect 12916 56544 12924 56608
rect 12604 55520 12924 56544
rect 12604 55456 12612 55520
rect 12676 55456 12692 55520
rect 12756 55456 12772 55520
rect 12836 55456 12852 55520
rect 12916 55456 12924 55520
rect 12604 54432 12924 55456
rect 12604 54368 12612 54432
rect 12676 54368 12692 54432
rect 12756 54368 12772 54432
rect 12836 54368 12852 54432
rect 12916 54368 12924 54432
rect 12604 53954 12924 54368
rect 12604 53718 12646 53954
rect 12882 53718 12924 53954
rect 12604 53344 12924 53718
rect 12604 53280 12612 53344
rect 12676 53280 12692 53344
rect 12756 53280 12772 53344
rect 12836 53280 12852 53344
rect 12916 53280 12924 53344
rect 12604 52256 12924 53280
rect 12604 52192 12612 52256
rect 12676 52192 12692 52256
rect 12756 52192 12772 52256
rect 12836 52192 12852 52256
rect 12916 52192 12924 52256
rect 12604 51168 12924 52192
rect 12604 51104 12612 51168
rect 12676 51104 12692 51168
rect 12756 51104 12772 51168
rect 12836 51104 12852 51168
rect 12916 51104 12924 51168
rect 12604 50080 12924 51104
rect 12604 50016 12612 50080
rect 12676 50016 12692 50080
rect 12756 50016 12772 50080
rect 12836 50016 12852 50080
rect 12916 50016 12924 50080
rect 12604 48992 12924 50016
rect 12604 48928 12612 48992
rect 12676 48954 12692 48992
rect 12756 48954 12772 48992
rect 12836 48954 12852 48992
rect 12916 48928 12924 48992
rect 12604 48718 12646 48928
rect 12882 48718 12924 48928
rect 12604 47904 12924 48718
rect 12604 47840 12612 47904
rect 12676 47840 12692 47904
rect 12756 47840 12772 47904
rect 12836 47840 12852 47904
rect 12916 47840 12924 47904
rect 12604 46816 12924 47840
rect 12604 46752 12612 46816
rect 12676 46752 12692 46816
rect 12756 46752 12772 46816
rect 12836 46752 12852 46816
rect 12916 46752 12924 46816
rect 12604 45728 12924 46752
rect 12604 45664 12612 45728
rect 12676 45664 12692 45728
rect 12756 45664 12772 45728
rect 12836 45664 12852 45728
rect 12916 45664 12924 45728
rect 12604 44640 12924 45664
rect 12604 44576 12612 44640
rect 12676 44576 12692 44640
rect 12756 44576 12772 44640
rect 12836 44576 12852 44640
rect 12916 44576 12924 44640
rect 12604 43954 12924 44576
rect 12604 43718 12646 43954
rect 12882 43718 12924 43954
rect 12604 43552 12924 43718
rect 12604 43488 12612 43552
rect 12676 43488 12692 43552
rect 12756 43488 12772 43552
rect 12836 43488 12852 43552
rect 12916 43488 12924 43552
rect 12604 42464 12924 43488
rect 12604 42400 12612 42464
rect 12676 42400 12692 42464
rect 12756 42400 12772 42464
rect 12836 42400 12852 42464
rect 12916 42400 12924 42464
rect 12604 41376 12924 42400
rect 12604 41312 12612 41376
rect 12676 41312 12692 41376
rect 12756 41312 12772 41376
rect 12836 41312 12852 41376
rect 12916 41312 12924 41376
rect 12604 40288 12924 41312
rect 12604 40224 12612 40288
rect 12676 40224 12692 40288
rect 12756 40224 12772 40288
rect 12836 40224 12852 40288
rect 12916 40224 12924 40288
rect 12604 39200 12924 40224
rect 12604 39136 12612 39200
rect 12676 39136 12692 39200
rect 12756 39136 12772 39200
rect 12836 39136 12852 39200
rect 12916 39136 12924 39200
rect 12604 38954 12924 39136
rect 12604 38718 12646 38954
rect 12882 38718 12924 38954
rect 12604 38112 12924 38718
rect 12604 38048 12612 38112
rect 12676 38048 12692 38112
rect 12756 38048 12772 38112
rect 12836 38048 12852 38112
rect 12916 38048 12924 38112
rect 12604 37024 12924 38048
rect 12604 36960 12612 37024
rect 12676 36960 12692 37024
rect 12756 36960 12772 37024
rect 12836 36960 12852 37024
rect 12916 36960 12924 37024
rect 12604 35936 12924 36960
rect 12604 35872 12612 35936
rect 12676 35872 12692 35936
rect 12756 35872 12772 35936
rect 12836 35872 12852 35936
rect 12916 35872 12924 35936
rect 12604 34848 12924 35872
rect 12604 34784 12612 34848
rect 12676 34784 12692 34848
rect 12756 34784 12772 34848
rect 12836 34784 12852 34848
rect 12916 34784 12924 34848
rect 12604 33954 12924 34784
rect 12604 33760 12646 33954
rect 12882 33760 12924 33954
rect 12604 33696 12612 33760
rect 12676 33696 12692 33718
rect 12756 33696 12772 33718
rect 12836 33696 12852 33718
rect 12916 33696 12924 33760
rect 12604 32672 12924 33696
rect 12604 32608 12612 32672
rect 12676 32608 12692 32672
rect 12756 32608 12772 32672
rect 12836 32608 12852 32672
rect 12916 32608 12924 32672
rect 12604 31584 12924 32608
rect 12604 31520 12612 31584
rect 12676 31520 12692 31584
rect 12756 31520 12772 31584
rect 12836 31520 12852 31584
rect 12916 31520 12924 31584
rect 12604 30496 12924 31520
rect 12604 30432 12612 30496
rect 12676 30432 12692 30496
rect 12756 30432 12772 30496
rect 12836 30432 12852 30496
rect 12916 30432 12924 30496
rect 12604 29408 12924 30432
rect 12604 29344 12612 29408
rect 12676 29344 12692 29408
rect 12756 29344 12772 29408
rect 12836 29344 12852 29408
rect 12916 29344 12924 29408
rect 12604 28954 12924 29344
rect 12604 28718 12646 28954
rect 12882 28718 12924 28954
rect 12604 28320 12924 28718
rect 12604 28256 12612 28320
rect 12676 28256 12692 28320
rect 12756 28256 12772 28320
rect 12836 28256 12852 28320
rect 12916 28256 12924 28320
rect 12604 27232 12924 28256
rect 12604 27168 12612 27232
rect 12676 27168 12692 27232
rect 12756 27168 12772 27232
rect 12836 27168 12852 27232
rect 12916 27168 12924 27232
rect 12604 26144 12924 27168
rect 12604 26080 12612 26144
rect 12676 26080 12692 26144
rect 12756 26080 12772 26144
rect 12836 26080 12852 26144
rect 12916 26080 12924 26144
rect 12604 25056 12924 26080
rect 12604 24992 12612 25056
rect 12676 24992 12692 25056
rect 12756 24992 12772 25056
rect 12836 24992 12852 25056
rect 12916 24992 12924 25056
rect 12604 23968 12924 24992
rect 12604 23904 12612 23968
rect 12676 23954 12692 23968
rect 12756 23954 12772 23968
rect 12836 23954 12852 23968
rect 12916 23904 12924 23968
rect 12604 23718 12646 23904
rect 12882 23718 12924 23904
rect 12604 22880 12924 23718
rect 12604 22816 12612 22880
rect 12676 22816 12692 22880
rect 12756 22816 12772 22880
rect 12836 22816 12852 22880
rect 12916 22816 12924 22880
rect 12604 21792 12924 22816
rect 14966 22813 15026 67763
rect 16944 66944 17264 67968
rect 16944 66880 16952 66944
rect 17016 66880 17032 66944
rect 17096 66880 17112 66944
rect 17176 66880 17192 66944
rect 17256 66880 17264 66944
rect 16944 65856 17264 66880
rect 16944 65792 16952 65856
rect 17016 65792 17032 65856
rect 17096 65792 17112 65856
rect 17176 65792 17192 65856
rect 17256 65792 17264 65856
rect 16944 64768 17264 65792
rect 16944 64704 16952 64768
rect 17016 64704 17032 64768
rect 17096 64704 17112 64768
rect 17176 64704 17192 64768
rect 17256 64704 17264 64768
rect 16944 63680 17264 64704
rect 16944 63616 16952 63680
rect 17016 63616 17032 63680
rect 17096 63616 17112 63680
rect 17176 63616 17192 63680
rect 17256 63616 17264 63680
rect 16944 63294 17264 63616
rect 16944 63058 16986 63294
rect 17222 63058 17264 63294
rect 16944 62592 17264 63058
rect 16944 62528 16952 62592
rect 17016 62528 17032 62592
rect 17096 62528 17112 62592
rect 17176 62528 17192 62592
rect 17256 62528 17264 62592
rect 16944 61504 17264 62528
rect 16944 61440 16952 61504
rect 17016 61440 17032 61504
rect 17096 61440 17112 61504
rect 17176 61440 17192 61504
rect 17256 61440 17264 61504
rect 16944 60416 17264 61440
rect 16944 60352 16952 60416
rect 17016 60352 17032 60416
rect 17096 60352 17112 60416
rect 17176 60352 17192 60416
rect 17256 60352 17264 60416
rect 16944 59328 17264 60352
rect 16944 59264 16952 59328
rect 17016 59264 17032 59328
rect 17096 59264 17112 59328
rect 17176 59264 17192 59328
rect 17256 59264 17264 59328
rect 16944 58294 17264 59264
rect 16944 58240 16986 58294
rect 17222 58240 17264 58294
rect 16944 58176 16952 58240
rect 17256 58176 17264 58240
rect 16944 58058 16986 58176
rect 17222 58058 17264 58176
rect 16944 57152 17264 58058
rect 16944 57088 16952 57152
rect 17016 57088 17032 57152
rect 17096 57088 17112 57152
rect 17176 57088 17192 57152
rect 17256 57088 17264 57152
rect 16944 56064 17264 57088
rect 16944 56000 16952 56064
rect 17016 56000 17032 56064
rect 17096 56000 17112 56064
rect 17176 56000 17192 56064
rect 17256 56000 17264 56064
rect 16435 55316 16501 55317
rect 16435 55252 16436 55316
rect 16500 55252 16501 55316
rect 16435 55251 16501 55252
rect 14963 22812 15029 22813
rect 14963 22748 14964 22812
rect 15028 22748 15029 22812
rect 14963 22747 15029 22748
rect 12604 21728 12612 21792
rect 12676 21728 12692 21792
rect 12756 21728 12772 21792
rect 12836 21728 12852 21792
rect 12916 21728 12924 21792
rect 12604 20704 12924 21728
rect 12604 20640 12612 20704
rect 12676 20640 12692 20704
rect 12756 20640 12772 20704
rect 12836 20640 12852 20704
rect 12916 20640 12924 20704
rect 12604 19616 12924 20640
rect 12604 19552 12612 19616
rect 12676 19552 12692 19616
rect 12756 19552 12772 19616
rect 12836 19552 12852 19616
rect 12916 19552 12924 19616
rect 12604 18954 12924 19552
rect 12604 18718 12646 18954
rect 12882 18718 12924 18954
rect 12604 18528 12924 18718
rect 12604 18464 12612 18528
rect 12676 18464 12692 18528
rect 12756 18464 12772 18528
rect 12836 18464 12852 18528
rect 12916 18464 12924 18528
rect 12604 17440 12924 18464
rect 12604 17376 12612 17440
rect 12676 17376 12692 17440
rect 12756 17376 12772 17440
rect 12836 17376 12852 17440
rect 12916 17376 12924 17440
rect 12604 16352 12924 17376
rect 12604 16288 12612 16352
rect 12676 16288 12692 16352
rect 12756 16288 12772 16352
rect 12836 16288 12852 16352
rect 12916 16288 12924 16352
rect 12604 15264 12924 16288
rect 12604 15200 12612 15264
rect 12676 15200 12692 15264
rect 12756 15200 12772 15264
rect 12836 15200 12852 15264
rect 12916 15200 12924 15264
rect 12604 14176 12924 15200
rect 12604 14112 12612 14176
rect 12676 14112 12692 14176
rect 12756 14112 12772 14176
rect 12836 14112 12852 14176
rect 12916 14112 12924 14176
rect 12604 13954 12924 14112
rect 12604 13718 12646 13954
rect 12882 13718 12924 13954
rect 12604 13088 12924 13718
rect 12604 13024 12612 13088
rect 12676 13024 12692 13088
rect 12756 13024 12772 13088
rect 12836 13024 12852 13088
rect 12916 13024 12924 13088
rect 12604 12000 12924 13024
rect 12604 11936 12612 12000
rect 12676 11936 12692 12000
rect 12756 11936 12772 12000
rect 12836 11936 12852 12000
rect 12916 11936 12924 12000
rect 12604 10912 12924 11936
rect 12604 10848 12612 10912
rect 12676 10848 12692 10912
rect 12756 10848 12772 10912
rect 12836 10848 12852 10912
rect 12916 10848 12924 10912
rect 12604 9824 12924 10848
rect 12604 9760 12612 9824
rect 12676 9760 12692 9824
rect 12756 9760 12772 9824
rect 12836 9760 12852 9824
rect 12916 9760 12924 9824
rect 12604 8954 12924 9760
rect 12604 8736 12646 8954
rect 12882 8736 12924 8954
rect 12604 8672 12612 8736
rect 12676 8672 12692 8718
rect 12756 8672 12772 8718
rect 12836 8672 12852 8718
rect 12916 8672 12924 8736
rect 12604 7648 12924 8672
rect 12604 7584 12612 7648
rect 12676 7584 12692 7648
rect 12756 7584 12772 7648
rect 12836 7584 12852 7648
rect 12916 7584 12924 7648
rect 12604 6560 12924 7584
rect 12604 6496 12612 6560
rect 12676 6496 12692 6560
rect 12756 6496 12772 6560
rect 12836 6496 12852 6560
rect 12916 6496 12924 6560
rect 12604 5472 12924 6496
rect 12604 5408 12612 5472
rect 12676 5408 12692 5472
rect 12756 5408 12772 5472
rect 12836 5408 12852 5472
rect 12916 5408 12924 5472
rect 12604 4384 12924 5408
rect 12604 4320 12612 4384
rect 12676 4320 12692 4384
rect 12756 4320 12772 4384
rect 12836 4320 12852 4384
rect 12916 4320 12924 4384
rect 12604 3954 12924 4320
rect 12604 3718 12646 3954
rect 12882 3718 12924 3954
rect 12604 3296 12924 3718
rect 12604 3232 12612 3296
rect 12676 3232 12692 3296
rect 12756 3232 12772 3296
rect 12836 3232 12852 3296
rect 12916 3232 12924 3296
rect 12604 2208 12924 3232
rect 16438 2413 16498 55251
rect 16944 54976 17264 56000
rect 16944 54912 16952 54976
rect 17016 54912 17032 54976
rect 17096 54912 17112 54976
rect 17176 54912 17192 54976
rect 17256 54912 17264 54976
rect 16944 53888 17264 54912
rect 16944 53824 16952 53888
rect 17016 53824 17032 53888
rect 17096 53824 17112 53888
rect 17176 53824 17192 53888
rect 17256 53824 17264 53888
rect 16944 53294 17264 53824
rect 16944 53058 16986 53294
rect 17222 53058 17264 53294
rect 16944 52800 17264 53058
rect 16944 52736 16952 52800
rect 17016 52736 17032 52800
rect 17096 52736 17112 52800
rect 17176 52736 17192 52800
rect 17256 52736 17264 52800
rect 16944 51712 17264 52736
rect 16944 51648 16952 51712
rect 17016 51648 17032 51712
rect 17096 51648 17112 51712
rect 17176 51648 17192 51712
rect 17256 51648 17264 51712
rect 16944 50624 17264 51648
rect 16944 50560 16952 50624
rect 17016 50560 17032 50624
rect 17096 50560 17112 50624
rect 17176 50560 17192 50624
rect 17256 50560 17264 50624
rect 16944 49536 17264 50560
rect 16944 49472 16952 49536
rect 17016 49472 17032 49536
rect 17096 49472 17112 49536
rect 17176 49472 17192 49536
rect 17256 49472 17264 49536
rect 16944 48448 17264 49472
rect 16944 48384 16952 48448
rect 17016 48384 17032 48448
rect 17096 48384 17112 48448
rect 17176 48384 17192 48448
rect 17256 48384 17264 48448
rect 16944 48294 17264 48384
rect 16944 48058 16986 48294
rect 17222 48058 17264 48294
rect 16944 47360 17264 48058
rect 16944 47296 16952 47360
rect 17016 47296 17032 47360
rect 17096 47296 17112 47360
rect 17176 47296 17192 47360
rect 17256 47296 17264 47360
rect 16944 46272 17264 47296
rect 16944 46208 16952 46272
rect 17016 46208 17032 46272
rect 17096 46208 17112 46272
rect 17176 46208 17192 46272
rect 17256 46208 17264 46272
rect 16944 45184 17264 46208
rect 16944 45120 16952 45184
rect 17016 45120 17032 45184
rect 17096 45120 17112 45184
rect 17176 45120 17192 45184
rect 17256 45120 17264 45184
rect 16944 44096 17264 45120
rect 16944 44032 16952 44096
rect 17016 44032 17032 44096
rect 17096 44032 17112 44096
rect 17176 44032 17192 44096
rect 17256 44032 17264 44096
rect 16944 43294 17264 44032
rect 16944 43058 16986 43294
rect 17222 43058 17264 43294
rect 16944 43008 17264 43058
rect 16944 42944 16952 43008
rect 17016 42944 17032 43008
rect 17096 42944 17112 43008
rect 17176 42944 17192 43008
rect 17256 42944 17264 43008
rect 16944 41920 17264 42944
rect 16944 41856 16952 41920
rect 17016 41856 17032 41920
rect 17096 41856 17112 41920
rect 17176 41856 17192 41920
rect 17256 41856 17264 41920
rect 16944 40832 17264 41856
rect 16944 40768 16952 40832
rect 17016 40768 17032 40832
rect 17096 40768 17112 40832
rect 17176 40768 17192 40832
rect 17256 40768 17264 40832
rect 16944 39744 17264 40768
rect 16944 39680 16952 39744
rect 17016 39680 17032 39744
rect 17096 39680 17112 39744
rect 17176 39680 17192 39744
rect 17256 39680 17264 39744
rect 16944 38656 17264 39680
rect 16944 38592 16952 38656
rect 17016 38592 17032 38656
rect 17096 38592 17112 38656
rect 17176 38592 17192 38656
rect 17256 38592 17264 38656
rect 16944 38294 17264 38592
rect 16944 38058 16986 38294
rect 17222 38058 17264 38294
rect 16944 37568 17264 38058
rect 16944 37504 16952 37568
rect 17016 37504 17032 37568
rect 17096 37504 17112 37568
rect 17176 37504 17192 37568
rect 17256 37504 17264 37568
rect 16944 36480 17264 37504
rect 16944 36416 16952 36480
rect 17016 36416 17032 36480
rect 17096 36416 17112 36480
rect 17176 36416 17192 36480
rect 17256 36416 17264 36480
rect 16944 35392 17264 36416
rect 16944 35328 16952 35392
rect 17016 35328 17032 35392
rect 17096 35328 17112 35392
rect 17176 35328 17192 35392
rect 17256 35328 17264 35392
rect 16944 34304 17264 35328
rect 16944 34240 16952 34304
rect 17016 34240 17032 34304
rect 17096 34240 17112 34304
rect 17176 34240 17192 34304
rect 17256 34240 17264 34304
rect 16944 33294 17264 34240
rect 16944 33216 16986 33294
rect 17222 33216 17264 33294
rect 16944 33152 16952 33216
rect 17256 33152 17264 33216
rect 16944 33058 16986 33152
rect 17222 33058 17264 33152
rect 16944 32128 17264 33058
rect 16944 32064 16952 32128
rect 17016 32064 17032 32128
rect 17096 32064 17112 32128
rect 17176 32064 17192 32128
rect 17256 32064 17264 32128
rect 16944 31040 17264 32064
rect 16944 30976 16952 31040
rect 17016 30976 17032 31040
rect 17096 30976 17112 31040
rect 17176 30976 17192 31040
rect 17256 30976 17264 31040
rect 16944 29952 17264 30976
rect 16944 29888 16952 29952
rect 17016 29888 17032 29952
rect 17096 29888 17112 29952
rect 17176 29888 17192 29952
rect 17256 29888 17264 29952
rect 16944 28864 17264 29888
rect 16944 28800 16952 28864
rect 17016 28800 17032 28864
rect 17096 28800 17112 28864
rect 17176 28800 17192 28864
rect 17256 28800 17264 28864
rect 16944 28294 17264 28800
rect 16944 28058 16986 28294
rect 17222 28058 17264 28294
rect 16944 27776 17264 28058
rect 16944 27712 16952 27776
rect 17016 27712 17032 27776
rect 17096 27712 17112 27776
rect 17176 27712 17192 27776
rect 17256 27712 17264 27776
rect 16944 26688 17264 27712
rect 16944 26624 16952 26688
rect 17016 26624 17032 26688
rect 17096 26624 17112 26688
rect 17176 26624 17192 26688
rect 17256 26624 17264 26688
rect 16944 25600 17264 26624
rect 16944 25536 16952 25600
rect 17016 25536 17032 25600
rect 17096 25536 17112 25600
rect 17176 25536 17192 25600
rect 17256 25536 17264 25600
rect 16944 24512 17264 25536
rect 16944 24448 16952 24512
rect 17016 24448 17032 24512
rect 17096 24448 17112 24512
rect 17176 24448 17192 24512
rect 17256 24448 17264 24512
rect 16944 23424 17264 24448
rect 16944 23360 16952 23424
rect 17016 23360 17032 23424
rect 17096 23360 17112 23424
rect 17176 23360 17192 23424
rect 17256 23360 17264 23424
rect 16944 23294 17264 23360
rect 16944 23058 16986 23294
rect 17222 23058 17264 23294
rect 16944 22336 17264 23058
rect 16944 22272 16952 22336
rect 17016 22272 17032 22336
rect 17096 22272 17112 22336
rect 17176 22272 17192 22336
rect 17256 22272 17264 22336
rect 16944 21248 17264 22272
rect 16944 21184 16952 21248
rect 17016 21184 17032 21248
rect 17096 21184 17112 21248
rect 17176 21184 17192 21248
rect 17256 21184 17264 21248
rect 16944 20160 17264 21184
rect 16944 20096 16952 20160
rect 17016 20096 17032 20160
rect 17096 20096 17112 20160
rect 17176 20096 17192 20160
rect 17256 20096 17264 20160
rect 16944 19072 17264 20096
rect 16944 19008 16952 19072
rect 17016 19008 17032 19072
rect 17096 19008 17112 19072
rect 17176 19008 17192 19072
rect 17256 19008 17264 19072
rect 16944 18294 17264 19008
rect 16944 18058 16986 18294
rect 17222 18058 17264 18294
rect 16944 17984 17264 18058
rect 16944 17920 16952 17984
rect 17016 17920 17032 17984
rect 17096 17920 17112 17984
rect 17176 17920 17192 17984
rect 17256 17920 17264 17984
rect 16944 16896 17264 17920
rect 16944 16832 16952 16896
rect 17016 16832 17032 16896
rect 17096 16832 17112 16896
rect 17176 16832 17192 16896
rect 17256 16832 17264 16896
rect 16944 15808 17264 16832
rect 16944 15744 16952 15808
rect 17016 15744 17032 15808
rect 17096 15744 17112 15808
rect 17176 15744 17192 15808
rect 17256 15744 17264 15808
rect 16944 14720 17264 15744
rect 16944 14656 16952 14720
rect 17016 14656 17032 14720
rect 17096 14656 17112 14720
rect 17176 14656 17192 14720
rect 17256 14656 17264 14720
rect 16944 13632 17264 14656
rect 16944 13568 16952 13632
rect 17016 13568 17032 13632
rect 17096 13568 17112 13632
rect 17176 13568 17192 13632
rect 17256 13568 17264 13632
rect 16944 13294 17264 13568
rect 16944 13058 16986 13294
rect 17222 13058 17264 13294
rect 16944 12544 17264 13058
rect 16944 12480 16952 12544
rect 17016 12480 17032 12544
rect 17096 12480 17112 12544
rect 17176 12480 17192 12544
rect 17256 12480 17264 12544
rect 16944 11456 17264 12480
rect 16944 11392 16952 11456
rect 17016 11392 17032 11456
rect 17096 11392 17112 11456
rect 17176 11392 17192 11456
rect 17256 11392 17264 11456
rect 16944 10368 17264 11392
rect 16944 10304 16952 10368
rect 17016 10304 17032 10368
rect 17096 10304 17112 10368
rect 17176 10304 17192 10368
rect 17256 10304 17264 10368
rect 16944 9280 17264 10304
rect 16944 9216 16952 9280
rect 17016 9216 17032 9280
rect 17096 9216 17112 9280
rect 17176 9216 17192 9280
rect 17256 9216 17264 9280
rect 16944 8294 17264 9216
rect 16944 8192 16986 8294
rect 17222 8192 17264 8294
rect 16944 8128 16952 8192
rect 17256 8128 17264 8192
rect 16944 8058 16986 8128
rect 17222 8058 17264 8128
rect 16944 7104 17264 8058
rect 16944 7040 16952 7104
rect 17016 7040 17032 7104
rect 17096 7040 17112 7104
rect 17176 7040 17192 7104
rect 17256 7040 17264 7104
rect 16944 6016 17264 7040
rect 16944 5952 16952 6016
rect 17016 5952 17032 6016
rect 17096 5952 17112 6016
rect 17176 5952 17192 6016
rect 17256 5952 17264 6016
rect 16944 4928 17264 5952
rect 16944 4864 16952 4928
rect 17016 4864 17032 4928
rect 17096 4864 17112 4928
rect 17176 4864 17192 4928
rect 17256 4864 17264 4928
rect 16944 3840 17264 4864
rect 16944 3776 16952 3840
rect 17016 3776 17032 3840
rect 17096 3776 17112 3840
rect 17176 3776 17192 3840
rect 17256 3776 17264 3840
rect 16944 3294 17264 3776
rect 16944 3058 16986 3294
rect 17222 3058 17264 3294
rect 16944 2752 17264 3058
rect 16944 2688 16952 2752
rect 17016 2688 17032 2752
rect 17096 2688 17112 2752
rect 17176 2688 17192 2752
rect 17256 2688 17264 2752
rect 16435 2412 16501 2413
rect 16435 2348 16436 2412
rect 16500 2348 16501 2412
rect 16435 2347 16501 2348
rect 12604 2144 12612 2208
rect 12676 2144 12692 2208
rect 12756 2144 12772 2208
rect 12836 2144 12852 2208
rect 12916 2144 12924 2208
rect 12604 2128 12924 2144
rect 16944 2128 17264 2688
rect 17604 69664 17924 69680
rect 17604 69600 17612 69664
rect 17676 69600 17692 69664
rect 17756 69600 17772 69664
rect 17836 69600 17852 69664
rect 17916 69600 17924 69664
rect 17604 68954 17924 69600
rect 17604 68718 17646 68954
rect 17882 68718 17924 68954
rect 17604 68576 17924 68718
rect 17604 68512 17612 68576
rect 17676 68512 17692 68576
rect 17756 68512 17772 68576
rect 17836 68512 17852 68576
rect 17916 68512 17924 68576
rect 17604 67488 17924 68512
rect 17604 67424 17612 67488
rect 17676 67424 17692 67488
rect 17756 67424 17772 67488
rect 17836 67424 17852 67488
rect 17916 67424 17924 67488
rect 17604 66400 17924 67424
rect 17604 66336 17612 66400
rect 17676 66336 17692 66400
rect 17756 66336 17772 66400
rect 17836 66336 17852 66400
rect 17916 66336 17924 66400
rect 17604 65312 17924 66336
rect 17604 65248 17612 65312
rect 17676 65248 17692 65312
rect 17756 65248 17772 65312
rect 17836 65248 17852 65312
rect 17916 65248 17924 65312
rect 17604 64224 17924 65248
rect 17604 64160 17612 64224
rect 17676 64160 17692 64224
rect 17756 64160 17772 64224
rect 17836 64160 17852 64224
rect 17916 64160 17924 64224
rect 17604 63954 17924 64160
rect 17604 63718 17646 63954
rect 17882 63718 17924 63954
rect 17604 63136 17924 63718
rect 21944 69120 22264 69680
rect 21944 69056 21952 69120
rect 22016 69056 22032 69120
rect 22096 69056 22112 69120
rect 22176 69056 22192 69120
rect 22256 69056 22264 69120
rect 21944 68294 22264 69056
rect 21944 68058 21986 68294
rect 22222 68058 22264 68294
rect 21944 68032 22264 68058
rect 21944 67968 21952 68032
rect 22016 67968 22032 68032
rect 22096 67968 22112 68032
rect 22176 67968 22192 68032
rect 22256 67968 22264 68032
rect 21944 66944 22264 67968
rect 21944 66880 21952 66944
rect 22016 66880 22032 66944
rect 22096 66880 22112 66944
rect 22176 66880 22192 66944
rect 22256 66880 22264 66944
rect 21944 65856 22264 66880
rect 21944 65792 21952 65856
rect 22016 65792 22032 65856
rect 22096 65792 22112 65856
rect 22176 65792 22192 65856
rect 22256 65792 22264 65856
rect 21944 64768 22264 65792
rect 21944 64704 21952 64768
rect 22016 64704 22032 64768
rect 22096 64704 22112 64768
rect 22176 64704 22192 64768
rect 22256 64704 22264 64768
rect 21944 63680 22264 64704
rect 21944 63616 21952 63680
rect 22016 63616 22032 63680
rect 22096 63616 22112 63680
rect 22176 63616 22192 63680
rect 22256 63616 22264 63680
rect 20483 63612 20549 63613
rect 20483 63548 20484 63612
rect 20548 63548 20549 63612
rect 20483 63547 20549 63548
rect 21587 63612 21653 63613
rect 21587 63548 21588 63612
rect 21652 63548 21653 63612
rect 21587 63547 21653 63548
rect 17604 63072 17612 63136
rect 17676 63072 17692 63136
rect 17756 63072 17772 63136
rect 17836 63072 17852 63136
rect 17916 63072 17924 63136
rect 17604 62048 17924 63072
rect 17604 61984 17612 62048
rect 17676 61984 17692 62048
rect 17756 61984 17772 62048
rect 17836 61984 17852 62048
rect 17916 61984 17924 62048
rect 17604 60960 17924 61984
rect 17604 60896 17612 60960
rect 17676 60896 17692 60960
rect 17756 60896 17772 60960
rect 17836 60896 17852 60960
rect 17916 60896 17924 60960
rect 17604 59872 17924 60896
rect 17604 59808 17612 59872
rect 17676 59808 17692 59872
rect 17756 59808 17772 59872
rect 17836 59808 17852 59872
rect 17916 59808 17924 59872
rect 17604 58954 17924 59808
rect 17604 58784 17646 58954
rect 17882 58784 17924 58954
rect 17604 58720 17612 58784
rect 17916 58720 17924 58784
rect 17604 58718 17646 58720
rect 17882 58718 17924 58720
rect 17604 57696 17924 58718
rect 17604 57632 17612 57696
rect 17676 57632 17692 57696
rect 17756 57632 17772 57696
rect 17836 57632 17852 57696
rect 17916 57632 17924 57696
rect 17604 56608 17924 57632
rect 18459 56812 18525 56813
rect 18459 56748 18460 56812
rect 18524 56748 18525 56812
rect 18459 56747 18525 56748
rect 17604 56544 17612 56608
rect 17676 56544 17692 56608
rect 17756 56544 17772 56608
rect 17836 56544 17852 56608
rect 17916 56544 17924 56608
rect 17604 55520 17924 56544
rect 17604 55456 17612 55520
rect 17676 55456 17692 55520
rect 17756 55456 17772 55520
rect 17836 55456 17852 55520
rect 17916 55456 17924 55520
rect 17604 54432 17924 55456
rect 17604 54368 17612 54432
rect 17676 54368 17692 54432
rect 17756 54368 17772 54432
rect 17836 54368 17852 54432
rect 17916 54368 17924 54432
rect 17604 53954 17924 54368
rect 17604 53718 17646 53954
rect 17882 53718 17924 53954
rect 17604 53344 17924 53718
rect 17604 53280 17612 53344
rect 17676 53280 17692 53344
rect 17756 53280 17772 53344
rect 17836 53280 17852 53344
rect 17916 53280 17924 53344
rect 17604 52256 17924 53280
rect 17604 52192 17612 52256
rect 17676 52192 17692 52256
rect 17756 52192 17772 52256
rect 17836 52192 17852 52256
rect 17916 52192 17924 52256
rect 17604 51168 17924 52192
rect 17604 51104 17612 51168
rect 17676 51104 17692 51168
rect 17756 51104 17772 51168
rect 17836 51104 17852 51168
rect 17916 51104 17924 51168
rect 17604 50080 17924 51104
rect 17604 50016 17612 50080
rect 17676 50016 17692 50080
rect 17756 50016 17772 50080
rect 17836 50016 17852 50080
rect 17916 50016 17924 50080
rect 17604 48992 17924 50016
rect 17604 48928 17612 48992
rect 17676 48954 17692 48992
rect 17756 48954 17772 48992
rect 17836 48954 17852 48992
rect 17916 48928 17924 48992
rect 17604 48718 17646 48928
rect 17882 48718 17924 48928
rect 17604 47904 17924 48718
rect 17604 47840 17612 47904
rect 17676 47840 17692 47904
rect 17756 47840 17772 47904
rect 17836 47840 17852 47904
rect 17916 47840 17924 47904
rect 17604 46816 17924 47840
rect 17604 46752 17612 46816
rect 17676 46752 17692 46816
rect 17756 46752 17772 46816
rect 17836 46752 17852 46816
rect 17916 46752 17924 46816
rect 17604 45728 17924 46752
rect 17604 45664 17612 45728
rect 17676 45664 17692 45728
rect 17756 45664 17772 45728
rect 17836 45664 17852 45728
rect 17916 45664 17924 45728
rect 17604 44640 17924 45664
rect 17604 44576 17612 44640
rect 17676 44576 17692 44640
rect 17756 44576 17772 44640
rect 17836 44576 17852 44640
rect 17916 44576 17924 44640
rect 17604 43954 17924 44576
rect 17604 43718 17646 43954
rect 17882 43718 17924 43954
rect 17604 43552 17924 43718
rect 17604 43488 17612 43552
rect 17676 43488 17692 43552
rect 17756 43488 17772 43552
rect 17836 43488 17852 43552
rect 17916 43488 17924 43552
rect 17604 42464 17924 43488
rect 17604 42400 17612 42464
rect 17676 42400 17692 42464
rect 17756 42400 17772 42464
rect 17836 42400 17852 42464
rect 17916 42400 17924 42464
rect 17604 41376 17924 42400
rect 17604 41312 17612 41376
rect 17676 41312 17692 41376
rect 17756 41312 17772 41376
rect 17836 41312 17852 41376
rect 17916 41312 17924 41376
rect 17604 40288 17924 41312
rect 17604 40224 17612 40288
rect 17676 40224 17692 40288
rect 17756 40224 17772 40288
rect 17836 40224 17852 40288
rect 17916 40224 17924 40288
rect 17604 39200 17924 40224
rect 17604 39136 17612 39200
rect 17676 39136 17692 39200
rect 17756 39136 17772 39200
rect 17836 39136 17852 39200
rect 17916 39136 17924 39200
rect 17604 38954 17924 39136
rect 17604 38718 17646 38954
rect 17882 38718 17924 38954
rect 17604 38112 17924 38718
rect 17604 38048 17612 38112
rect 17676 38048 17692 38112
rect 17756 38048 17772 38112
rect 17836 38048 17852 38112
rect 17916 38048 17924 38112
rect 17604 37024 17924 38048
rect 17604 36960 17612 37024
rect 17676 36960 17692 37024
rect 17756 36960 17772 37024
rect 17836 36960 17852 37024
rect 17916 36960 17924 37024
rect 17604 35936 17924 36960
rect 17604 35872 17612 35936
rect 17676 35872 17692 35936
rect 17756 35872 17772 35936
rect 17836 35872 17852 35936
rect 17916 35872 17924 35936
rect 17604 34848 17924 35872
rect 17604 34784 17612 34848
rect 17676 34784 17692 34848
rect 17756 34784 17772 34848
rect 17836 34784 17852 34848
rect 17916 34784 17924 34848
rect 17604 33954 17924 34784
rect 17604 33760 17646 33954
rect 17882 33760 17924 33954
rect 17604 33696 17612 33760
rect 17676 33696 17692 33718
rect 17756 33696 17772 33718
rect 17836 33696 17852 33718
rect 17916 33696 17924 33760
rect 17604 32672 17924 33696
rect 17604 32608 17612 32672
rect 17676 32608 17692 32672
rect 17756 32608 17772 32672
rect 17836 32608 17852 32672
rect 17916 32608 17924 32672
rect 17604 31584 17924 32608
rect 17604 31520 17612 31584
rect 17676 31520 17692 31584
rect 17756 31520 17772 31584
rect 17836 31520 17852 31584
rect 17916 31520 17924 31584
rect 17604 30496 17924 31520
rect 17604 30432 17612 30496
rect 17676 30432 17692 30496
rect 17756 30432 17772 30496
rect 17836 30432 17852 30496
rect 17916 30432 17924 30496
rect 17604 29408 17924 30432
rect 17604 29344 17612 29408
rect 17676 29344 17692 29408
rect 17756 29344 17772 29408
rect 17836 29344 17852 29408
rect 17916 29344 17924 29408
rect 17604 28954 17924 29344
rect 17604 28718 17646 28954
rect 17882 28718 17924 28954
rect 17604 28320 17924 28718
rect 17604 28256 17612 28320
rect 17676 28256 17692 28320
rect 17756 28256 17772 28320
rect 17836 28256 17852 28320
rect 17916 28256 17924 28320
rect 17604 27232 17924 28256
rect 17604 27168 17612 27232
rect 17676 27168 17692 27232
rect 17756 27168 17772 27232
rect 17836 27168 17852 27232
rect 17916 27168 17924 27232
rect 17604 26144 17924 27168
rect 18462 26349 18522 56747
rect 18459 26348 18525 26349
rect 18459 26284 18460 26348
rect 18524 26284 18525 26348
rect 18459 26283 18525 26284
rect 17604 26080 17612 26144
rect 17676 26080 17692 26144
rect 17756 26080 17772 26144
rect 17836 26080 17852 26144
rect 17916 26080 17924 26144
rect 17604 25056 17924 26080
rect 17604 24992 17612 25056
rect 17676 24992 17692 25056
rect 17756 24992 17772 25056
rect 17836 24992 17852 25056
rect 17916 24992 17924 25056
rect 17604 23968 17924 24992
rect 17604 23904 17612 23968
rect 17676 23954 17692 23968
rect 17756 23954 17772 23968
rect 17836 23954 17852 23968
rect 17916 23904 17924 23968
rect 17604 23718 17646 23904
rect 17882 23718 17924 23904
rect 17604 22880 17924 23718
rect 17604 22816 17612 22880
rect 17676 22816 17692 22880
rect 17756 22816 17772 22880
rect 17836 22816 17852 22880
rect 17916 22816 17924 22880
rect 17604 21792 17924 22816
rect 17604 21728 17612 21792
rect 17676 21728 17692 21792
rect 17756 21728 17772 21792
rect 17836 21728 17852 21792
rect 17916 21728 17924 21792
rect 17604 20704 17924 21728
rect 17604 20640 17612 20704
rect 17676 20640 17692 20704
rect 17756 20640 17772 20704
rect 17836 20640 17852 20704
rect 17916 20640 17924 20704
rect 17604 19616 17924 20640
rect 17604 19552 17612 19616
rect 17676 19552 17692 19616
rect 17756 19552 17772 19616
rect 17836 19552 17852 19616
rect 17916 19552 17924 19616
rect 17604 18954 17924 19552
rect 17604 18718 17646 18954
rect 17882 18718 17924 18954
rect 17604 18528 17924 18718
rect 17604 18464 17612 18528
rect 17676 18464 17692 18528
rect 17756 18464 17772 18528
rect 17836 18464 17852 18528
rect 17916 18464 17924 18528
rect 17604 17440 17924 18464
rect 17604 17376 17612 17440
rect 17676 17376 17692 17440
rect 17756 17376 17772 17440
rect 17836 17376 17852 17440
rect 17916 17376 17924 17440
rect 17604 16352 17924 17376
rect 17604 16288 17612 16352
rect 17676 16288 17692 16352
rect 17756 16288 17772 16352
rect 17836 16288 17852 16352
rect 17916 16288 17924 16352
rect 17604 15264 17924 16288
rect 17604 15200 17612 15264
rect 17676 15200 17692 15264
rect 17756 15200 17772 15264
rect 17836 15200 17852 15264
rect 17916 15200 17924 15264
rect 17604 14176 17924 15200
rect 17604 14112 17612 14176
rect 17676 14112 17692 14176
rect 17756 14112 17772 14176
rect 17836 14112 17852 14176
rect 17916 14112 17924 14176
rect 17604 13954 17924 14112
rect 17604 13718 17646 13954
rect 17882 13718 17924 13954
rect 17604 13088 17924 13718
rect 17604 13024 17612 13088
rect 17676 13024 17692 13088
rect 17756 13024 17772 13088
rect 17836 13024 17852 13088
rect 17916 13024 17924 13088
rect 17604 12000 17924 13024
rect 20486 12205 20546 63547
rect 21590 13429 21650 63547
rect 21944 63294 22264 63616
rect 21944 63058 21986 63294
rect 22222 63058 22264 63294
rect 21944 62592 22264 63058
rect 21944 62528 21952 62592
rect 22016 62528 22032 62592
rect 22096 62528 22112 62592
rect 22176 62528 22192 62592
rect 22256 62528 22264 62592
rect 21944 61504 22264 62528
rect 21944 61440 21952 61504
rect 22016 61440 22032 61504
rect 22096 61440 22112 61504
rect 22176 61440 22192 61504
rect 22256 61440 22264 61504
rect 21944 60416 22264 61440
rect 21944 60352 21952 60416
rect 22016 60352 22032 60416
rect 22096 60352 22112 60416
rect 22176 60352 22192 60416
rect 22256 60352 22264 60416
rect 21944 59328 22264 60352
rect 21944 59264 21952 59328
rect 22016 59264 22032 59328
rect 22096 59264 22112 59328
rect 22176 59264 22192 59328
rect 22256 59264 22264 59328
rect 21944 58294 22264 59264
rect 21944 58240 21986 58294
rect 22222 58240 22264 58294
rect 21944 58176 21952 58240
rect 22256 58176 22264 58240
rect 21944 58058 21986 58176
rect 22222 58058 22264 58176
rect 21944 57152 22264 58058
rect 21944 57088 21952 57152
rect 22016 57088 22032 57152
rect 22096 57088 22112 57152
rect 22176 57088 22192 57152
rect 22256 57088 22264 57152
rect 21944 56064 22264 57088
rect 21944 56000 21952 56064
rect 22016 56000 22032 56064
rect 22096 56000 22112 56064
rect 22176 56000 22192 56064
rect 22256 56000 22264 56064
rect 21944 54976 22264 56000
rect 21944 54912 21952 54976
rect 22016 54912 22032 54976
rect 22096 54912 22112 54976
rect 22176 54912 22192 54976
rect 22256 54912 22264 54976
rect 21944 53888 22264 54912
rect 21944 53824 21952 53888
rect 22016 53824 22032 53888
rect 22096 53824 22112 53888
rect 22176 53824 22192 53888
rect 22256 53824 22264 53888
rect 21944 53294 22264 53824
rect 21944 53058 21986 53294
rect 22222 53058 22264 53294
rect 21944 52800 22264 53058
rect 21944 52736 21952 52800
rect 22016 52736 22032 52800
rect 22096 52736 22112 52800
rect 22176 52736 22192 52800
rect 22256 52736 22264 52800
rect 21944 51712 22264 52736
rect 21944 51648 21952 51712
rect 22016 51648 22032 51712
rect 22096 51648 22112 51712
rect 22176 51648 22192 51712
rect 22256 51648 22264 51712
rect 21944 50624 22264 51648
rect 21944 50560 21952 50624
rect 22016 50560 22032 50624
rect 22096 50560 22112 50624
rect 22176 50560 22192 50624
rect 22256 50560 22264 50624
rect 21944 49536 22264 50560
rect 21944 49472 21952 49536
rect 22016 49472 22032 49536
rect 22096 49472 22112 49536
rect 22176 49472 22192 49536
rect 22256 49472 22264 49536
rect 21944 48448 22264 49472
rect 21944 48384 21952 48448
rect 22016 48384 22032 48448
rect 22096 48384 22112 48448
rect 22176 48384 22192 48448
rect 22256 48384 22264 48448
rect 21944 48294 22264 48384
rect 21944 48058 21986 48294
rect 22222 48058 22264 48294
rect 21944 47360 22264 48058
rect 21944 47296 21952 47360
rect 22016 47296 22032 47360
rect 22096 47296 22112 47360
rect 22176 47296 22192 47360
rect 22256 47296 22264 47360
rect 21944 46272 22264 47296
rect 21944 46208 21952 46272
rect 22016 46208 22032 46272
rect 22096 46208 22112 46272
rect 22176 46208 22192 46272
rect 22256 46208 22264 46272
rect 21944 45184 22264 46208
rect 21944 45120 21952 45184
rect 22016 45120 22032 45184
rect 22096 45120 22112 45184
rect 22176 45120 22192 45184
rect 22256 45120 22264 45184
rect 21944 44096 22264 45120
rect 21944 44032 21952 44096
rect 22016 44032 22032 44096
rect 22096 44032 22112 44096
rect 22176 44032 22192 44096
rect 22256 44032 22264 44096
rect 21944 43294 22264 44032
rect 21944 43058 21986 43294
rect 22222 43058 22264 43294
rect 21944 43008 22264 43058
rect 21944 42944 21952 43008
rect 22016 42944 22032 43008
rect 22096 42944 22112 43008
rect 22176 42944 22192 43008
rect 22256 42944 22264 43008
rect 21944 41920 22264 42944
rect 21944 41856 21952 41920
rect 22016 41856 22032 41920
rect 22096 41856 22112 41920
rect 22176 41856 22192 41920
rect 22256 41856 22264 41920
rect 21944 40832 22264 41856
rect 21944 40768 21952 40832
rect 22016 40768 22032 40832
rect 22096 40768 22112 40832
rect 22176 40768 22192 40832
rect 22256 40768 22264 40832
rect 21944 39744 22264 40768
rect 21944 39680 21952 39744
rect 22016 39680 22032 39744
rect 22096 39680 22112 39744
rect 22176 39680 22192 39744
rect 22256 39680 22264 39744
rect 21944 38656 22264 39680
rect 21944 38592 21952 38656
rect 22016 38592 22032 38656
rect 22096 38592 22112 38656
rect 22176 38592 22192 38656
rect 22256 38592 22264 38656
rect 21944 38294 22264 38592
rect 21944 38058 21986 38294
rect 22222 38058 22264 38294
rect 21944 37568 22264 38058
rect 21944 37504 21952 37568
rect 22016 37504 22032 37568
rect 22096 37504 22112 37568
rect 22176 37504 22192 37568
rect 22256 37504 22264 37568
rect 21944 36480 22264 37504
rect 21944 36416 21952 36480
rect 22016 36416 22032 36480
rect 22096 36416 22112 36480
rect 22176 36416 22192 36480
rect 22256 36416 22264 36480
rect 21944 35392 22264 36416
rect 21944 35328 21952 35392
rect 22016 35328 22032 35392
rect 22096 35328 22112 35392
rect 22176 35328 22192 35392
rect 22256 35328 22264 35392
rect 21944 34304 22264 35328
rect 21944 34240 21952 34304
rect 22016 34240 22032 34304
rect 22096 34240 22112 34304
rect 22176 34240 22192 34304
rect 22256 34240 22264 34304
rect 21944 33294 22264 34240
rect 21944 33216 21986 33294
rect 22222 33216 22264 33294
rect 21944 33152 21952 33216
rect 22256 33152 22264 33216
rect 21944 33058 21986 33152
rect 22222 33058 22264 33152
rect 21944 32128 22264 33058
rect 21944 32064 21952 32128
rect 22016 32064 22032 32128
rect 22096 32064 22112 32128
rect 22176 32064 22192 32128
rect 22256 32064 22264 32128
rect 21944 31040 22264 32064
rect 21944 30976 21952 31040
rect 22016 30976 22032 31040
rect 22096 30976 22112 31040
rect 22176 30976 22192 31040
rect 22256 30976 22264 31040
rect 21944 29952 22264 30976
rect 21944 29888 21952 29952
rect 22016 29888 22032 29952
rect 22096 29888 22112 29952
rect 22176 29888 22192 29952
rect 22256 29888 22264 29952
rect 21944 28864 22264 29888
rect 21944 28800 21952 28864
rect 22016 28800 22032 28864
rect 22096 28800 22112 28864
rect 22176 28800 22192 28864
rect 22256 28800 22264 28864
rect 21944 28294 22264 28800
rect 21944 28058 21986 28294
rect 22222 28058 22264 28294
rect 21944 27776 22264 28058
rect 21944 27712 21952 27776
rect 22016 27712 22032 27776
rect 22096 27712 22112 27776
rect 22176 27712 22192 27776
rect 22256 27712 22264 27776
rect 21944 26688 22264 27712
rect 21944 26624 21952 26688
rect 22016 26624 22032 26688
rect 22096 26624 22112 26688
rect 22176 26624 22192 26688
rect 22256 26624 22264 26688
rect 21944 25600 22264 26624
rect 21944 25536 21952 25600
rect 22016 25536 22032 25600
rect 22096 25536 22112 25600
rect 22176 25536 22192 25600
rect 22256 25536 22264 25600
rect 21944 24512 22264 25536
rect 21944 24448 21952 24512
rect 22016 24448 22032 24512
rect 22096 24448 22112 24512
rect 22176 24448 22192 24512
rect 22256 24448 22264 24512
rect 21944 23424 22264 24448
rect 21944 23360 21952 23424
rect 22016 23360 22032 23424
rect 22096 23360 22112 23424
rect 22176 23360 22192 23424
rect 22256 23360 22264 23424
rect 21944 23294 22264 23360
rect 21944 23058 21986 23294
rect 22222 23058 22264 23294
rect 21944 22336 22264 23058
rect 21944 22272 21952 22336
rect 22016 22272 22032 22336
rect 22096 22272 22112 22336
rect 22176 22272 22192 22336
rect 22256 22272 22264 22336
rect 21944 21248 22264 22272
rect 21944 21184 21952 21248
rect 22016 21184 22032 21248
rect 22096 21184 22112 21248
rect 22176 21184 22192 21248
rect 22256 21184 22264 21248
rect 21944 20160 22264 21184
rect 21944 20096 21952 20160
rect 22016 20096 22032 20160
rect 22096 20096 22112 20160
rect 22176 20096 22192 20160
rect 22256 20096 22264 20160
rect 21944 19072 22264 20096
rect 21944 19008 21952 19072
rect 22016 19008 22032 19072
rect 22096 19008 22112 19072
rect 22176 19008 22192 19072
rect 22256 19008 22264 19072
rect 21944 18294 22264 19008
rect 21944 18058 21986 18294
rect 22222 18058 22264 18294
rect 21944 17984 22264 18058
rect 21944 17920 21952 17984
rect 22016 17920 22032 17984
rect 22096 17920 22112 17984
rect 22176 17920 22192 17984
rect 22256 17920 22264 17984
rect 21944 16896 22264 17920
rect 21944 16832 21952 16896
rect 22016 16832 22032 16896
rect 22096 16832 22112 16896
rect 22176 16832 22192 16896
rect 22256 16832 22264 16896
rect 21944 15808 22264 16832
rect 21944 15744 21952 15808
rect 22016 15744 22032 15808
rect 22096 15744 22112 15808
rect 22176 15744 22192 15808
rect 22256 15744 22264 15808
rect 21944 14720 22264 15744
rect 21944 14656 21952 14720
rect 22016 14656 22032 14720
rect 22096 14656 22112 14720
rect 22176 14656 22192 14720
rect 22256 14656 22264 14720
rect 21944 13632 22264 14656
rect 21944 13568 21952 13632
rect 22016 13568 22032 13632
rect 22096 13568 22112 13632
rect 22176 13568 22192 13632
rect 22256 13568 22264 13632
rect 21587 13428 21653 13429
rect 21587 13364 21588 13428
rect 21652 13364 21653 13428
rect 21587 13363 21653 13364
rect 21944 13294 22264 13568
rect 21944 13058 21986 13294
rect 22222 13058 22264 13294
rect 21944 12544 22264 13058
rect 21944 12480 21952 12544
rect 22016 12480 22032 12544
rect 22096 12480 22112 12544
rect 22176 12480 22192 12544
rect 22256 12480 22264 12544
rect 20483 12204 20549 12205
rect 20483 12140 20484 12204
rect 20548 12140 20549 12204
rect 20483 12139 20549 12140
rect 17604 11936 17612 12000
rect 17676 11936 17692 12000
rect 17756 11936 17772 12000
rect 17836 11936 17852 12000
rect 17916 11936 17924 12000
rect 17604 10912 17924 11936
rect 17604 10848 17612 10912
rect 17676 10848 17692 10912
rect 17756 10848 17772 10912
rect 17836 10848 17852 10912
rect 17916 10848 17924 10912
rect 17604 9824 17924 10848
rect 17604 9760 17612 9824
rect 17676 9760 17692 9824
rect 17756 9760 17772 9824
rect 17836 9760 17852 9824
rect 17916 9760 17924 9824
rect 17604 8954 17924 9760
rect 17604 8736 17646 8954
rect 17882 8736 17924 8954
rect 17604 8672 17612 8736
rect 17676 8672 17692 8718
rect 17756 8672 17772 8718
rect 17836 8672 17852 8718
rect 17916 8672 17924 8736
rect 17604 7648 17924 8672
rect 17604 7584 17612 7648
rect 17676 7584 17692 7648
rect 17756 7584 17772 7648
rect 17836 7584 17852 7648
rect 17916 7584 17924 7648
rect 17604 6560 17924 7584
rect 17604 6496 17612 6560
rect 17676 6496 17692 6560
rect 17756 6496 17772 6560
rect 17836 6496 17852 6560
rect 17916 6496 17924 6560
rect 17604 5472 17924 6496
rect 17604 5408 17612 5472
rect 17676 5408 17692 5472
rect 17756 5408 17772 5472
rect 17836 5408 17852 5472
rect 17916 5408 17924 5472
rect 17604 4384 17924 5408
rect 17604 4320 17612 4384
rect 17676 4320 17692 4384
rect 17756 4320 17772 4384
rect 17836 4320 17852 4384
rect 17916 4320 17924 4384
rect 17604 3954 17924 4320
rect 17604 3718 17646 3954
rect 17882 3718 17924 3954
rect 17604 3296 17924 3718
rect 17604 3232 17612 3296
rect 17676 3232 17692 3296
rect 17756 3232 17772 3296
rect 17836 3232 17852 3296
rect 17916 3232 17924 3296
rect 17604 2208 17924 3232
rect 17604 2144 17612 2208
rect 17676 2144 17692 2208
rect 17756 2144 17772 2208
rect 17836 2144 17852 2208
rect 17916 2144 17924 2208
rect 17604 2128 17924 2144
rect 21944 11456 22264 12480
rect 21944 11392 21952 11456
rect 22016 11392 22032 11456
rect 22096 11392 22112 11456
rect 22176 11392 22192 11456
rect 22256 11392 22264 11456
rect 21944 10368 22264 11392
rect 21944 10304 21952 10368
rect 22016 10304 22032 10368
rect 22096 10304 22112 10368
rect 22176 10304 22192 10368
rect 22256 10304 22264 10368
rect 21944 9280 22264 10304
rect 21944 9216 21952 9280
rect 22016 9216 22032 9280
rect 22096 9216 22112 9280
rect 22176 9216 22192 9280
rect 22256 9216 22264 9280
rect 21944 8294 22264 9216
rect 21944 8192 21986 8294
rect 22222 8192 22264 8294
rect 21944 8128 21952 8192
rect 22256 8128 22264 8192
rect 21944 8058 21986 8128
rect 22222 8058 22264 8128
rect 21944 7104 22264 8058
rect 21944 7040 21952 7104
rect 22016 7040 22032 7104
rect 22096 7040 22112 7104
rect 22176 7040 22192 7104
rect 22256 7040 22264 7104
rect 21944 6016 22264 7040
rect 21944 5952 21952 6016
rect 22016 5952 22032 6016
rect 22096 5952 22112 6016
rect 22176 5952 22192 6016
rect 22256 5952 22264 6016
rect 21944 4928 22264 5952
rect 21944 4864 21952 4928
rect 22016 4864 22032 4928
rect 22096 4864 22112 4928
rect 22176 4864 22192 4928
rect 22256 4864 22264 4928
rect 21944 3840 22264 4864
rect 21944 3776 21952 3840
rect 22016 3776 22032 3840
rect 22096 3776 22112 3840
rect 22176 3776 22192 3840
rect 22256 3776 22264 3840
rect 21944 3294 22264 3776
rect 21944 3058 21986 3294
rect 22222 3058 22264 3294
rect 21944 2752 22264 3058
rect 21944 2688 21952 2752
rect 22016 2688 22032 2752
rect 22096 2688 22112 2752
rect 22176 2688 22192 2752
rect 22256 2688 22264 2752
rect 21944 2128 22264 2688
rect 22604 69664 22924 69680
rect 22604 69600 22612 69664
rect 22676 69600 22692 69664
rect 22756 69600 22772 69664
rect 22836 69600 22852 69664
rect 22916 69600 22924 69664
rect 22604 68954 22924 69600
rect 22604 68718 22646 68954
rect 22882 68718 22924 68954
rect 22604 68576 22924 68718
rect 22604 68512 22612 68576
rect 22676 68512 22692 68576
rect 22756 68512 22772 68576
rect 22836 68512 22852 68576
rect 22916 68512 22924 68576
rect 22604 67488 22924 68512
rect 22604 67424 22612 67488
rect 22676 67424 22692 67488
rect 22756 67424 22772 67488
rect 22836 67424 22852 67488
rect 22916 67424 22924 67488
rect 22604 66400 22924 67424
rect 22604 66336 22612 66400
rect 22676 66336 22692 66400
rect 22756 66336 22772 66400
rect 22836 66336 22852 66400
rect 22916 66336 22924 66400
rect 22604 65312 22924 66336
rect 26944 69120 27264 69680
rect 26944 69056 26952 69120
rect 27016 69056 27032 69120
rect 27096 69056 27112 69120
rect 27176 69056 27192 69120
rect 27256 69056 27264 69120
rect 26944 68294 27264 69056
rect 26944 68058 26986 68294
rect 27222 68058 27264 68294
rect 26944 68032 27264 68058
rect 26944 67968 26952 68032
rect 27016 67968 27032 68032
rect 27096 67968 27112 68032
rect 27176 67968 27192 68032
rect 27256 67968 27264 68032
rect 26944 66944 27264 67968
rect 26944 66880 26952 66944
rect 27016 66880 27032 66944
rect 27096 66880 27112 66944
rect 27176 66880 27192 66944
rect 27256 66880 27264 66944
rect 26944 65856 27264 66880
rect 26944 65792 26952 65856
rect 27016 65792 27032 65856
rect 27096 65792 27112 65856
rect 27176 65792 27192 65856
rect 27256 65792 27264 65856
rect 23611 65516 23677 65517
rect 23611 65452 23612 65516
rect 23676 65452 23677 65516
rect 23611 65451 23677 65452
rect 22604 65248 22612 65312
rect 22676 65248 22692 65312
rect 22756 65248 22772 65312
rect 22836 65248 22852 65312
rect 22916 65248 22924 65312
rect 22604 64224 22924 65248
rect 22604 64160 22612 64224
rect 22676 64160 22692 64224
rect 22756 64160 22772 64224
rect 22836 64160 22852 64224
rect 22916 64160 22924 64224
rect 22604 63954 22924 64160
rect 22604 63718 22646 63954
rect 22882 63718 22924 63954
rect 22604 63136 22924 63718
rect 22604 63072 22612 63136
rect 22676 63072 22692 63136
rect 22756 63072 22772 63136
rect 22836 63072 22852 63136
rect 22916 63072 22924 63136
rect 22604 62048 22924 63072
rect 22604 61984 22612 62048
rect 22676 61984 22692 62048
rect 22756 61984 22772 62048
rect 22836 61984 22852 62048
rect 22916 61984 22924 62048
rect 22604 60960 22924 61984
rect 22604 60896 22612 60960
rect 22676 60896 22692 60960
rect 22756 60896 22772 60960
rect 22836 60896 22852 60960
rect 22916 60896 22924 60960
rect 22604 59872 22924 60896
rect 22604 59808 22612 59872
rect 22676 59808 22692 59872
rect 22756 59808 22772 59872
rect 22836 59808 22852 59872
rect 22916 59808 22924 59872
rect 22604 58954 22924 59808
rect 22604 58784 22646 58954
rect 22882 58784 22924 58954
rect 22604 58720 22612 58784
rect 22916 58720 22924 58784
rect 22604 58718 22646 58720
rect 22882 58718 22924 58720
rect 22604 57696 22924 58718
rect 22604 57632 22612 57696
rect 22676 57632 22692 57696
rect 22756 57632 22772 57696
rect 22836 57632 22852 57696
rect 22916 57632 22924 57696
rect 22604 56608 22924 57632
rect 22604 56544 22612 56608
rect 22676 56544 22692 56608
rect 22756 56544 22772 56608
rect 22836 56544 22852 56608
rect 22916 56544 22924 56608
rect 22604 55520 22924 56544
rect 22604 55456 22612 55520
rect 22676 55456 22692 55520
rect 22756 55456 22772 55520
rect 22836 55456 22852 55520
rect 22916 55456 22924 55520
rect 22604 54432 22924 55456
rect 22604 54368 22612 54432
rect 22676 54368 22692 54432
rect 22756 54368 22772 54432
rect 22836 54368 22852 54432
rect 22916 54368 22924 54432
rect 22604 53954 22924 54368
rect 22604 53718 22646 53954
rect 22882 53718 22924 53954
rect 22604 53344 22924 53718
rect 22604 53280 22612 53344
rect 22676 53280 22692 53344
rect 22756 53280 22772 53344
rect 22836 53280 22852 53344
rect 22916 53280 22924 53344
rect 22604 52256 22924 53280
rect 22604 52192 22612 52256
rect 22676 52192 22692 52256
rect 22756 52192 22772 52256
rect 22836 52192 22852 52256
rect 22916 52192 22924 52256
rect 22604 51168 22924 52192
rect 22604 51104 22612 51168
rect 22676 51104 22692 51168
rect 22756 51104 22772 51168
rect 22836 51104 22852 51168
rect 22916 51104 22924 51168
rect 22604 50080 22924 51104
rect 22604 50016 22612 50080
rect 22676 50016 22692 50080
rect 22756 50016 22772 50080
rect 22836 50016 22852 50080
rect 22916 50016 22924 50080
rect 22604 48992 22924 50016
rect 22604 48928 22612 48992
rect 22676 48954 22692 48992
rect 22756 48954 22772 48992
rect 22836 48954 22852 48992
rect 22916 48928 22924 48992
rect 22604 48718 22646 48928
rect 22882 48718 22924 48928
rect 22604 47904 22924 48718
rect 22604 47840 22612 47904
rect 22676 47840 22692 47904
rect 22756 47840 22772 47904
rect 22836 47840 22852 47904
rect 22916 47840 22924 47904
rect 22604 46816 22924 47840
rect 22604 46752 22612 46816
rect 22676 46752 22692 46816
rect 22756 46752 22772 46816
rect 22836 46752 22852 46816
rect 22916 46752 22924 46816
rect 22604 45728 22924 46752
rect 22604 45664 22612 45728
rect 22676 45664 22692 45728
rect 22756 45664 22772 45728
rect 22836 45664 22852 45728
rect 22916 45664 22924 45728
rect 22604 44640 22924 45664
rect 22604 44576 22612 44640
rect 22676 44576 22692 44640
rect 22756 44576 22772 44640
rect 22836 44576 22852 44640
rect 22916 44576 22924 44640
rect 22604 43954 22924 44576
rect 22604 43718 22646 43954
rect 22882 43718 22924 43954
rect 22604 43552 22924 43718
rect 22604 43488 22612 43552
rect 22676 43488 22692 43552
rect 22756 43488 22772 43552
rect 22836 43488 22852 43552
rect 22916 43488 22924 43552
rect 22604 42464 22924 43488
rect 22604 42400 22612 42464
rect 22676 42400 22692 42464
rect 22756 42400 22772 42464
rect 22836 42400 22852 42464
rect 22916 42400 22924 42464
rect 22604 41376 22924 42400
rect 22604 41312 22612 41376
rect 22676 41312 22692 41376
rect 22756 41312 22772 41376
rect 22836 41312 22852 41376
rect 22916 41312 22924 41376
rect 22604 40288 22924 41312
rect 23614 40629 23674 65451
rect 26944 64768 27264 65792
rect 26944 64704 26952 64768
rect 27016 64704 27032 64768
rect 27096 64704 27112 64768
rect 27176 64704 27192 64768
rect 27256 64704 27264 64768
rect 26944 63680 27264 64704
rect 26944 63616 26952 63680
rect 27016 63616 27032 63680
rect 27096 63616 27112 63680
rect 27176 63616 27192 63680
rect 27256 63616 27264 63680
rect 26944 63294 27264 63616
rect 26944 63058 26986 63294
rect 27222 63058 27264 63294
rect 24715 62796 24781 62797
rect 24715 62732 24716 62796
rect 24780 62732 24781 62796
rect 24715 62731 24781 62732
rect 23611 40628 23677 40629
rect 23611 40564 23612 40628
rect 23676 40564 23677 40628
rect 23611 40563 23677 40564
rect 22604 40224 22612 40288
rect 22676 40224 22692 40288
rect 22756 40224 22772 40288
rect 22836 40224 22852 40288
rect 22916 40224 22924 40288
rect 22604 39200 22924 40224
rect 22604 39136 22612 39200
rect 22676 39136 22692 39200
rect 22756 39136 22772 39200
rect 22836 39136 22852 39200
rect 22916 39136 22924 39200
rect 22604 38954 22924 39136
rect 22604 38718 22646 38954
rect 22882 38718 22924 38954
rect 22604 38112 22924 38718
rect 23243 38724 23309 38725
rect 23243 38660 23244 38724
rect 23308 38660 23309 38724
rect 23243 38659 23309 38660
rect 22604 38048 22612 38112
rect 22676 38048 22692 38112
rect 22756 38048 22772 38112
rect 22836 38048 22852 38112
rect 22916 38048 22924 38112
rect 22604 37024 22924 38048
rect 22604 36960 22612 37024
rect 22676 36960 22692 37024
rect 22756 36960 22772 37024
rect 22836 36960 22852 37024
rect 22916 36960 22924 37024
rect 22604 35936 22924 36960
rect 22604 35872 22612 35936
rect 22676 35872 22692 35936
rect 22756 35872 22772 35936
rect 22836 35872 22852 35936
rect 22916 35872 22924 35936
rect 22604 34848 22924 35872
rect 22604 34784 22612 34848
rect 22676 34784 22692 34848
rect 22756 34784 22772 34848
rect 22836 34784 22852 34848
rect 22916 34784 22924 34848
rect 22604 33954 22924 34784
rect 22604 33760 22646 33954
rect 22882 33760 22924 33954
rect 22604 33696 22612 33760
rect 22676 33696 22692 33718
rect 22756 33696 22772 33718
rect 22836 33696 22852 33718
rect 22916 33696 22924 33760
rect 22604 32672 22924 33696
rect 22604 32608 22612 32672
rect 22676 32608 22692 32672
rect 22756 32608 22772 32672
rect 22836 32608 22852 32672
rect 22916 32608 22924 32672
rect 22604 31584 22924 32608
rect 22604 31520 22612 31584
rect 22676 31520 22692 31584
rect 22756 31520 22772 31584
rect 22836 31520 22852 31584
rect 22916 31520 22924 31584
rect 22604 30496 22924 31520
rect 23246 31109 23306 38659
rect 24718 38453 24778 62731
rect 26944 62592 27264 63058
rect 26944 62528 26952 62592
rect 27016 62528 27032 62592
rect 27096 62528 27112 62592
rect 27176 62528 27192 62592
rect 27256 62528 27264 62592
rect 25267 61708 25333 61709
rect 25267 61644 25268 61708
rect 25332 61644 25333 61708
rect 25267 61643 25333 61644
rect 24899 59532 24965 59533
rect 24899 59468 24900 59532
rect 24964 59468 24965 59532
rect 24899 59467 24965 59468
rect 24715 38452 24781 38453
rect 24715 38388 24716 38452
rect 24780 38388 24781 38452
rect 24715 38387 24781 38388
rect 23243 31108 23309 31109
rect 23243 31044 23244 31108
rect 23308 31044 23309 31108
rect 23243 31043 23309 31044
rect 22604 30432 22612 30496
rect 22676 30432 22692 30496
rect 22756 30432 22772 30496
rect 22836 30432 22852 30496
rect 22916 30432 22924 30496
rect 22604 29408 22924 30432
rect 22604 29344 22612 29408
rect 22676 29344 22692 29408
rect 22756 29344 22772 29408
rect 22836 29344 22852 29408
rect 22916 29344 22924 29408
rect 22604 28954 22924 29344
rect 22604 28718 22646 28954
rect 22882 28718 22924 28954
rect 22604 28320 22924 28718
rect 22604 28256 22612 28320
rect 22676 28256 22692 28320
rect 22756 28256 22772 28320
rect 22836 28256 22852 28320
rect 22916 28256 22924 28320
rect 22604 27232 22924 28256
rect 22604 27168 22612 27232
rect 22676 27168 22692 27232
rect 22756 27168 22772 27232
rect 22836 27168 22852 27232
rect 22916 27168 22924 27232
rect 22604 26144 22924 27168
rect 22604 26080 22612 26144
rect 22676 26080 22692 26144
rect 22756 26080 22772 26144
rect 22836 26080 22852 26144
rect 22916 26080 22924 26144
rect 22604 25056 22924 26080
rect 22604 24992 22612 25056
rect 22676 24992 22692 25056
rect 22756 24992 22772 25056
rect 22836 24992 22852 25056
rect 22916 24992 22924 25056
rect 22604 23968 22924 24992
rect 22604 23904 22612 23968
rect 22676 23954 22692 23968
rect 22756 23954 22772 23968
rect 22836 23954 22852 23968
rect 22916 23904 22924 23968
rect 22604 23718 22646 23904
rect 22882 23718 22924 23904
rect 22604 22880 22924 23718
rect 22604 22816 22612 22880
rect 22676 22816 22692 22880
rect 22756 22816 22772 22880
rect 22836 22816 22852 22880
rect 22916 22816 22924 22880
rect 22604 21792 22924 22816
rect 22604 21728 22612 21792
rect 22676 21728 22692 21792
rect 22756 21728 22772 21792
rect 22836 21728 22852 21792
rect 22916 21728 22924 21792
rect 22604 20704 22924 21728
rect 22604 20640 22612 20704
rect 22676 20640 22692 20704
rect 22756 20640 22772 20704
rect 22836 20640 22852 20704
rect 22916 20640 22924 20704
rect 22604 19616 22924 20640
rect 22604 19552 22612 19616
rect 22676 19552 22692 19616
rect 22756 19552 22772 19616
rect 22836 19552 22852 19616
rect 22916 19552 22924 19616
rect 22604 18954 22924 19552
rect 22604 18718 22646 18954
rect 22882 18718 22924 18954
rect 22604 18528 22924 18718
rect 22604 18464 22612 18528
rect 22676 18464 22692 18528
rect 22756 18464 22772 18528
rect 22836 18464 22852 18528
rect 22916 18464 22924 18528
rect 22604 17440 22924 18464
rect 22604 17376 22612 17440
rect 22676 17376 22692 17440
rect 22756 17376 22772 17440
rect 22836 17376 22852 17440
rect 22916 17376 22924 17440
rect 22604 16352 22924 17376
rect 22604 16288 22612 16352
rect 22676 16288 22692 16352
rect 22756 16288 22772 16352
rect 22836 16288 22852 16352
rect 22916 16288 22924 16352
rect 22604 15264 22924 16288
rect 22604 15200 22612 15264
rect 22676 15200 22692 15264
rect 22756 15200 22772 15264
rect 22836 15200 22852 15264
rect 22916 15200 22924 15264
rect 22604 14176 22924 15200
rect 24902 15061 24962 59467
rect 25270 38045 25330 61643
rect 26944 61504 27264 62528
rect 26944 61440 26952 61504
rect 27016 61440 27032 61504
rect 27096 61440 27112 61504
rect 27176 61440 27192 61504
rect 27256 61440 27264 61504
rect 26944 60416 27264 61440
rect 26944 60352 26952 60416
rect 27016 60352 27032 60416
rect 27096 60352 27112 60416
rect 27176 60352 27192 60416
rect 27256 60352 27264 60416
rect 26944 59328 27264 60352
rect 26944 59264 26952 59328
rect 27016 59264 27032 59328
rect 27096 59264 27112 59328
rect 27176 59264 27192 59328
rect 27256 59264 27264 59328
rect 26944 58294 27264 59264
rect 26944 58240 26986 58294
rect 27222 58240 27264 58294
rect 26944 58176 26952 58240
rect 27256 58176 27264 58240
rect 26944 58058 26986 58176
rect 27222 58058 27264 58176
rect 26944 57152 27264 58058
rect 26944 57088 26952 57152
rect 27016 57088 27032 57152
rect 27096 57088 27112 57152
rect 27176 57088 27192 57152
rect 27256 57088 27264 57152
rect 26944 56064 27264 57088
rect 26944 56000 26952 56064
rect 27016 56000 27032 56064
rect 27096 56000 27112 56064
rect 27176 56000 27192 56064
rect 27256 56000 27264 56064
rect 26944 54976 27264 56000
rect 26944 54912 26952 54976
rect 27016 54912 27032 54976
rect 27096 54912 27112 54976
rect 27176 54912 27192 54976
rect 27256 54912 27264 54976
rect 26944 53888 27264 54912
rect 26944 53824 26952 53888
rect 27016 53824 27032 53888
rect 27096 53824 27112 53888
rect 27176 53824 27192 53888
rect 27256 53824 27264 53888
rect 26944 53294 27264 53824
rect 26944 53058 26986 53294
rect 27222 53058 27264 53294
rect 26944 52800 27264 53058
rect 26944 52736 26952 52800
rect 27016 52736 27032 52800
rect 27096 52736 27112 52800
rect 27176 52736 27192 52800
rect 27256 52736 27264 52800
rect 26944 51712 27264 52736
rect 26944 51648 26952 51712
rect 27016 51648 27032 51712
rect 27096 51648 27112 51712
rect 27176 51648 27192 51712
rect 27256 51648 27264 51712
rect 26944 50624 27264 51648
rect 26944 50560 26952 50624
rect 27016 50560 27032 50624
rect 27096 50560 27112 50624
rect 27176 50560 27192 50624
rect 27256 50560 27264 50624
rect 26944 49536 27264 50560
rect 26944 49472 26952 49536
rect 27016 49472 27032 49536
rect 27096 49472 27112 49536
rect 27176 49472 27192 49536
rect 27256 49472 27264 49536
rect 26944 48448 27264 49472
rect 26944 48384 26952 48448
rect 27016 48384 27032 48448
rect 27096 48384 27112 48448
rect 27176 48384 27192 48448
rect 27256 48384 27264 48448
rect 26944 48294 27264 48384
rect 26944 48058 26986 48294
rect 27222 48058 27264 48294
rect 26944 47360 27264 48058
rect 26944 47296 26952 47360
rect 27016 47296 27032 47360
rect 27096 47296 27112 47360
rect 27176 47296 27192 47360
rect 27256 47296 27264 47360
rect 26944 46272 27264 47296
rect 26944 46208 26952 46272
rect 27016 46208 27032 46272
rect 27096 46208 27112 46272
rect 27176 46208 27192 46272
rect 27256 46208 27264 46272
rect 26944 45184 27264 46208
rect 26944 45120 26952 45184
rect 27016 45120 27032 45184
rect 27096 45120 27112 45184
rect 27176 45120 27192 45184
rect 27256 45120 27264 45184
rect 26944 44096 27264 45120
rect 26944 44032 26952 44096
rect 27016 44032 27032 44096
rect 27096 44032 27112 44096
rect 27176 44032 27192 44096
rect 27256 44032 27264 44096
rect 26944 43294 27264 44032
rect 26944 43058 26986 43294
rect 27222 43058 27264 43294
rect 26944 43008 27264 43058
rect 26944 42944 26952 43008
rect 27016 42944 27032 43008
rect 27096 42944 27112 43008
rect 27176 42944 27192 43008
rect 27256 42944 27264 43008
rect 26944 41920 27264 42944
rect 26944 41856 26952 41920
rect 27016 41856 27032 41920
rect 27096 41856 27112 41920
rect 27176 41856 27192 41920
rect 27256 41856 27264 41920
rect 26944 40832 27264 41856
rect 26944 40768 26952 40832
rect 27016 40768 27032 40832
rect 27096 40768 27112 40832
rect 27176 40768 27192 40832
rect 27256 40768 27264 40832
rect 26944 39744 27264 40768
rect 26944 39680 26952 39744
rect 27016 39680 27032 39744
rect 27096 39680 27112 39744
rect 27176 39680 27192 39744
rect 27256 39680 27264 39744
rect 26944 38656 27264 39680
rect 26944 38592 26952 38656
rect 27016 38592 27032 38656
rect 27096 38592 27112 38656
rect 27176 38592 27192 38656
rect 27256 38592 27264 38656
rect 26944 38294 27264 38592
rect 26944 38058 26986 38294
rect 27222 38058 27264 38294
rect 25267 38044 25333 38045
rect 25267 37980 25268 38044
rect 25332 37980 25333 38044
rect 25267 37979 25333 37980
rect 26944 37568 27264 38058
rect 26944 37504 26952 37568
rect 27016 37504 27032 37568
rect 27096 37504 27112 37568
rect 27176 37504 27192 37568
rect 27256 37504 27264 37568
rect 26944 36480 27264 37504
rect 26944 36416 26952 36480
rect 27016 36416 27032 36480
rect 27096 36416 27112 36480
rect 27176 36416 27192 36480
rect 27256 36416 27264 36480
rect 26944 35392 27264 36416
rect 26944 35328 26952 35392
rect 27016 35328 27032 35392
rect 27096 35328 27112 35392
rect 27176 35328 27192 35392
rect 27256 35328 27264 35392
rect 26944 34304 27264 35328
rect 26944 34240 26952 34304
rect 27016 34240 27032 34304
rect 27096 34240 27112 34304
rect 27176 34240 27192 34304
rect 27256 34240 27264 34304
rect 26944 33294 27264 34240
rect 26944 33216 26986 33294
rect 27222 33216 27264 33294
rect 26944 33152 26952 33216
rect 27256 33152 27264 33216
rect 26944 33058 26986 33152
rect 27222 33058 27264 33152
rect 26944 32128 27264 33058
rect 26944 32064 26952 32128
rect 27016 32064 27032 32128
rect 27096 32064 27112 32128
rect 27176 32064 27192 32128
rect 27256 32064 27264 32128
rect 26944 31040 27264 32064
rect 26944 30976 26952 31040
rect 27016 30976 27032 31040
rect 27096 30976 27112 31040
rect 27176 30976 27192 31040
rect 27256 30976 27264 31040
rect 26944 29952 27264 30976
rect 26944 29888 26952 29952
rect 27016 29888 27032 29952
rect 27096 29888 27112 29952
rect 27176 29888 27192 29952
rect 27256 29888 27264 29952
rect 26944 28864 27264 29888
rect 26944 28800 26952 28864
rect 27016 28800 27032 28864
rect 27096 28800 27112 28864
rect 27176 28800 27192 28864
rect 27256 28800 27264 28864
rect 26944 28294 27264 28800
rect 26944 28058 26986 28294
rect 27222 28058 27264 28294
rect 26944 27776 27264 28058
rect 26944 27712 26952 27776
rect 27016 27712 27032 27776
rect 27096 27712 27112 27776
rect 27176 27712 27192 27776
rect 27256 27712 27264 27776
rect 26944 26688 27264 27712
rect 26944 26624 26952 26688
rect 27016 26624 27032 26688
rect 27096 26624 27112 26688
rect 27176 26624 27192 26688
rect 27256 26624 27264 26688
rect 26944 25600 27264 26624
rect 26944 25536 26952 25600
rect 27016 25536 27032 25600
rect 27096 25536 27112 25600
rect 27176 25536 27192 25600
rect 27256 25536 27264 25600
rect 26944 24512 27264 25536
rect 26944 24448 26952 24512
rect 27016 24448 27032 24512
rect 27096 24448 27112 24512
rect 27176 24448 27192 24512
rect 27256 24448 27264 24512
rect 26944 23424 27264 24448
rect 26944 23360 26952 23424
rect 27016 23360 27032 23424
rect 27096 23360 27112 23424
rect 27176 23360 27192 23424
rect 27256 23360 27264 23424
rect 26944 23294 27264 23360
rect 26944 23058 26986 23294
rect 27222 23058 27264 23294
rect 26944 22336 27264 23058
rect 26944 22272 26952 22336
rect 27016 22272 27032 22336
rect 27096 22272 27112 22336
rect 27176 22272 27192 22336
rect 27256 22272 27264 22336
rect 26944 21248 27264 22272
rect 26944 21184 26952 21248
rect 27016 21184 27032 21248
rect 27096 21184 27112 21248
rect 27176 21184 27192 21248
rect 27256 21184 27264 21248
rect 26944 20160 27264 21184
rect 26944 20096 26952 20160
rect 27016 20096 27032 20160
rect 27096 20096 27112 20160
rect 27176 20096 27192 20160
rect 27256 20096 27264 20160
rect 26944 19072 27264 20096
rect 26944 19008 26952 19072
rect 27016 19008 27032 19072
rect 27096 19008 27112 19072
rect 27176 19008 27192 19072
rect 27256 19008 27264 19072
rect 26944 18294 27264 19008
rect 26944 18058 26986 18294
rect 27222 18058 27264 18294
rect 26944 17984 27264 18058
rect 26944 17920 26952 17984
rect 27016 17920 27032 17984
rect 27096 17920 27112 17984
rect 27176 17920 27192 17984
rect 27256 17920 27264 17984
rect 26944 16896 27264 17920
rect 26944 16832 26952 16896
rect 27016 16832 27032 16896
rect 27096 16832 27112 16896
rect 27176 16832 27192 16896
rect 27256 16832 27264 16896
rect 26944 15808 27264 16832
rect 26944 15744 26952 15808
rect 27016 15744 27032 15808
rect 27096 15744 27112 15808
rect 27176 15744 27192 15808
rect 27256 15744 27264 15808
rect 24899 15060 24965 15061
rect 24899 14996 24900 15060
rect 24964 14996 24965 15060
rect 24899 14995 24965 14996
rect 22604 14112 22612 14176
rect 22676 14112 22692 14176
rect 22756 14112 22772 14176
rect 22836 14112 22852 14176
rect 22916 14112 22924 14176
rect 22604 13954 22924 14112
rect 22604 13718 22646 13954
rect 22882 13718 22924 13954
rect 22604 13088 22924 13718
rect 22604 13024 22612 13088
rect 22676 13024 22692 13088
rect 22756 13024 22772 13088
rect 22836 13024 22852 13088
rect 22916 13024 22924 13088
rect 22604 12000 22924 13024
rect 22604 11936 22612 12000
rect 22676 11936 22692 12000
rect 22756 11936 22772 12000
rect 22836 11936 22852 12000
rect 22916 11936 22924 12000
rect 22604 10912 22924 11936
rect 22604 10848 22612 10912
rect 22676 10848 22692 10912
rect 22756 10848 22772 10912
rect 22836 10848 22852 10912
rect 22916 10848 22924 10912
rect 22604 9824 22924 10848
rect 22604 9760 22612 9824
rect 22676 9760 22692 9824
rect 22756 9760 22772 9824
rect 22836 9760 22852 9824
rect 22916 9760 22924 9824
rect 22604 8954 22924 9760
rect 22604 8736 22646 8954
rect 22882 8736 22924 8954
rect 22604 8672 22612 8736
rect 22676 8672 22692 8718
rect 22756 8672 22772 8718
rect 22836 8672 22852 8718
rect 22916 8672 22924 8736
rect 22604 7648 22924 8672
rect 22604 7584 22612 7648
rect 22676 7584 22692 7648
rect 22756 7584 22772 7648
rect 22836 7584 22852 7648
rect 22916 7584 22924 7648
rect 22604 6560 22924 7584
rect 22604 6496 22612 6560
rect 22676 6496 22692 6560
rect 22756 6496 22772 6560
rect 22836 6496 22852 6560
rect 22916 6496 22924 6560
rect 22604 5472 22924 6496
rect 22604 5408 22612 5472
rect 22676 5408 22692 5472
rect 22756 5408 22772 5472
rect 22836 5408 22852 5472
rect 22916 5408 22924 5472
rect 22604 4384 22924 5408
rect 22604 4320 22612 4384
rect 22676 4320 22692 4384
rect 22756 4320 22772 4384
rect 22836 4320 22852 4384
rect 22916 4320 22924 4384
rect 22604 3954 22924 4320
rect 22604 3718 22646 3954
rect 22882 3718 22924 3954
rect 22604 3296 22924 3718
rect 22604 3232 22612 3296
rect 22676 3232 22692 3296
rect 22756 3232 22772 3296
rect 22836 3232 22852 3296
rect 22916 3232 22924 3296
rect 22604 2208 22924 3232
rect 22604 2144 22612 2208
rect 22676 2144 22692 2208
rect 22756 2144 22772 2208
rect 22836 2144 22852 2208
rect 22916 2144 22924 2208
rect 22604 2128 22924 2144
rect 26944 14720 27264 15744
rect 26944 14656 26952 14720
rect 27016 14656 27032 14720
rect 27096 14656 27112 14720
rect 27176 14656 27192 14720
rect 27256 14656 27264 14720
rect 26944 13632 27264 14656
rect 26944 13568 26952 13632
rect 27016 13568 27032 13632
rect 27096 13568 27112 13632
rect 27176 13568 27192 13632
rect 27256 13568 27264 13632
rect 26944 13294 27264 13568
rect 26944 13058 26986 13294
rect 27222 13058 27264 13294
rect 26944 12544 27264 13058
rect 26944 12480 26952 12544
rect 27016 12480 27032 12544
rect 27096 12480 27112 12544
rect 27176 12480 27192 12544
rect 27256 12480 27264 12544
rect 26944 11456 27264 12480
rect 26944 11392 26952 11456
rect 27016 11392 27032 11456
rect 27096 11392 27112 11456
rect 27176 11392 27192 11456
rect 27256 11392 27264 11456
rect 26944 10368 27264 11392
rect 26944 10304 26952 10368
rect 27016 10304 27032 10368
rect 27096 10304 27112 10368
rect 27176 10304 27192 10368
rect 27256 10304 27264 10368
rect 26944 9280 27264 10304
rect 26944 9216 26952 9280
rect 27016 9216 27032 9280
rect 27096 9216 27112 9280
rect 27176 9216 27192 9280
rect 27256 9216 27264 9280
rect 26944 8294 27264 9216
rect 26944 8192 26986 8294
rect 27222 8192 27264 8294
rect 26944 8128 26952 8192
rect 27256 8128 27264 8192
rect 26944 8058 26986 8128
rect 27222 8058 27264 8128
rect 26944 7104 27264 8058
rect 26944 7040 26952 7104
rect 27016 7040 27032 7104
rect 27096 7040 27112 7104
rect 27176 7040 27192 7104
rect 27256 7040 27264 7104
rect 26944 6016 27264 7040
rect 26944 5952 26952 6016
rect 27016 5952 27032 6016
rect 27096 5952 27112 6016
rect 27176 5952 27192 6016
rect 27256 5952 27264 6016
rect 26944 4928 27264 5952
rect 26944 4864 26952 4928
rect 27016 4864 27032 4928
rect 27096 4864 27112 4928
rect 27176 4864 27192 4928
rect 27256 4864 27264 4928
rect 26944 3840 27264 4864
rect 26944 3776 26952 3840
rect 27016 3776 27032 3840
rect 27096 3776 27112 3840
rect 27176 3776 27192 3840
rect 27256 3776 27264 3840
rect 26944 3294 27264 3776
rect 26944 3058 26986 3294
rect 27222 3058 27264 3294
rect 26944 2752 27264 3058
rect 26944 2688 26952 2752
rect 27016 2688 27032 2752
rect 27096 2688 27112 2752
rect 27176 2688 27192 2752
rect 27256 2688 27264 2752
rect 26944 2128 27264 2688
rect 27604 69664 27924 69680
rect 27604 69600 27612 69664
rect 27676 69600 27692 69664
rect 27756 69600 27772 69664
rect 27836 69600 27852 69664
rect 27916 69600 27924 69664
rect 27604 68954 27924 69600
rect 27604 68718 27646 68954
rect 27882 68718 27924 68954
rect 27604 68576 27924 68718
rect 27604 68512 27612 68576
rect 27676 68512 27692 68576
rect 27756 68512 27772 68576
rect 27836 68512 27852 68576
rect 27916 68512 27924 68576
rect 27604 67488 27924 68512
rect 27604 67424 27612 67488
rect 27676 67424 27692 67488
rect 27756 67424 27772 67488
rect 27836 67424 27852 67488
rect 27916 67424 27924 67488
rect 27604 66400 27924 67424
rect 27604 66336 27612 66400
rect 27676 66336 27692 66400
rect 27756 66336 27772 66400
rect 27836 66336 27852 66400
rect 27916 66336 27924 66400
rect 27604 65312 27924 66336
rect 27604 65248 27612 65312
rect 27676 65248 27692 65312
rect 27756 65248 27772 65312
rect 27836 65248 27852 65312
rect 27916 65248 27924 65312
rect 27604 64224 27924 65248
rect 27604 64160 27612 64224
rect 27676 64160 27692 64224
rect 27756 64160 27772 64224
rect 27836 64160 27852 64224
rect 27916 64160 27924 64224
rect 27604 63954 27924 64160
rect 27604 63718 27646 63954
rect 27882 63718 27924 63954
rect 27604 63136 27924 63718
rect 27604 63072 27612 63136
rect 27676 63072 27692 63136
rect 27756 63072 27772 63136
rect 27836 63072 27852 63136
rect 27916 63072 27924 63136
rect 27604 62048 27924 63072
rect 27604 61984 27612 62048
rect 27676 61984 27692 62048
rect 27756 61984 27772 62048
rect 27836 61984 27852 62048
rect 27916 61984 27924 62048
rect 27604 60960 27924 61984
rect 27604 60896 27612 60960
rect 27676 60896 27692 60960
rect 27756 60896 27772 60960
rect 27836 60896 27852 60960
rect 27916 60896 27924 60960
rect 27604 59872 27924 60896
rect 27604 59808 27612 59872
rect 27676 59808 27692 59872
rect 27756 59808 27772 59872
rect 27836 59808 27852 59872
rect 27916 59808 27924 59872
rect 27604 58954 27924 59808
rect 27604 58784 27646 58954
rect 27882 58784 27924 58954
rect 27604 58720 27612 58784
rect 27916 58720 27924 58784
rect 27604 58718 27646 58720
rect 27882 58718 27924 58720
rect 27604 57696 27924 58718
rect 27604 57632 27612 57696
rect 27676 57632 27692 57696
rect 27756 57632 27772 57696
rect 27836 57632 27852 57696
rect 27916 57632 27924 57696
rect 27604 56608 27924 57632
rect 27604 56544 27612 56608
rect 27676 56544 27692 56608
rect 27756 56544 27772 56608
rect 27836 56544 27852 56608
rect 27916 56544 27924 56608
rect 27604 55520 27924 56544
rect 27604 55456 27612 55520
rect 27676 55456 27692 55520
rect 27756 55456 27772 55520
rect 27836 55456 27852 55520
rect 27916 55456 27924 55520
rect 27604 54432 27924 55456
rect 27604 54368 27612 54432
rect 27676 54368 27692 54432
rect 27756 54368 27772 54432
rect 27836 54368 27852 54432
rect 27916 54368 27924 54432
rect 27604 53954 27924 54368
rect 27604 53718 27646 53954
rect 27882 53718 27924 53954
rect 27604 53344 27924 53718
rect 27604 53280 27612 53344
rect 27676 53280 27692 53344
rect 27756 53280 27772 53344
rect 27836 53280 27852 53344
rect 27916 53280 27924 53344
rect 27604 52256 27924 53280
rect 27604 52192 27612 52256
rect 27676 52192 27692 52256
rect 27756 52192 27772 52256
rect 27836 52192 27852 52256
rect 27916 52192 27924 52256
rect 27604 51168 27924 52192
rect 27604 51104 27612 51168
rect 27676 51104 27692 51168
rect 27756 51104 27772 51168
rect 27836 51104 27852 51168
rect 27916 51104 27924 51168
rect 27604 50080 27924 51104
rect 27604 50016 27612 50080
rect 27676 50016 27692 50080
rect 27756 50016 27772 50080
rect 27836 50016 27852 50080
rect 27916 50016 27924 50080
rect 27604 48992 27924 50016
rect 27604 48928 27612 48992
rect 27676 48954 27692 48992
rect 27756 48954 27772 48992
rect 27836 48954 27852 48992
rect 27916 48928 27924 48992
rect 27604 48718 27646 48928
rect 27882 48718 27924 48928
rect 27604 47904 27924 48718
rect 27604 47840 27612 47904
rect 27676 47840 27692 47904
rect 27756 47840 27772 47904
rect 27836 47840 27852 47904
rect 27916 47840 27924 47904
rect 27604 46816 27924 47840
rect 27604 46752 27612 46816
rect 27676 46752 27692 46816
rect 27756 46752 27772 46816
rect 27836 46752 27852 46816
rect 27916 46752 27924 46816
rect 27604 45728 27924 46752
rect 27604 45664 27612 45728
rect 27676 45664 27692 45728
rect 27756 45664 27772 45728
rect 27836 45664 27852 45728
rect 27916 45664 27924 45728
rect 27604 44640 27924 45664
rect 27604 44576 27612 44640
rect 27676 44576 27692 44640
rect 27756 44576 27772 44640
rect 27836 44576 27852 44640
rect 27916 44576 27924 44640
rect 27604 43954 27924 44576
rect 27604 43718 27646 43954
rect 27882 43718 27924 43954
rect 27604 43552 27924 43718
rect 27604 43488 27612 43552
rect 27676 43488 27692 43552
rect 27756 43488 27772 43552
rect 27836 43488 27852 43552
rect 27916 43488 27924 43552
rect 27604 42464 27924 43488
rect 27604 42400 27612 42464
rect 27676 42400 27692 42464
rect 27756 42400 27772 42464
rect 27836 42400 27852 42464
rect 27916 42400 27924 42464
rect 27604 41376 27924 42400
rect 27604 41312 27612 41376
rect 27676 41312 27692 41376
rect 27756 41312 27772 41376
rect 27836 41312 27852 41376
rect 27916 41312 27924 41376
rect 27604 40288 27924 41312
rect 27604 40224 27612 40288
rect 27676 40224 27692 40288
rect 27756 40224 27772 40288
rect 27836 40224 27852 40288
rect 27916 40224 27924 40288
rect 27604 39200 27924 40224
rect 31944 69120 32264 69680
rect 31944 69056 31952 69120
rect 32016 69056 32032 69120
rect 32096 69056 32112 69120
rect 32176 69056 32192 69120
rect 32256 69056 32264 69120
rect 31944 68294 32264 69056
rect 31944 68058 31986 68294
rect 32222 68058 32264 68294
rect 31944 68032 32264 68058
rect 31944 67968 31952 68032
rect 32016 67968 32032 68032
rect 32096 67968 32112 68032
rect 32176 67968 32192 68032
rect 32256 67968 32264 68032
rect 31944 66944 32264 67968
rect 31944 66880 31952 66944
rect 32016 66880 32032 66944
rect 32096 66880 32112 66944
rect 32176 66880 32192 66944
rect 32256 66880 32264 66944
rect 31944 65856 32264 66880
rect 31944 65792 31952 65856
rect 32016 65792 32032 65856
rect 32096 65792 32112 65856
rect 32176 65792 32192 65856
rect 32256 65792 32264 65856
rect 31944 64768 32264 65792
rect 31944 64704 31952 64768
rect 32016 64704 32032 64768
rect 32096 64704 32112 64768
rect 32176 64704 32192 64768
rect 32256 64704 32264 64768
rect 31944 63680 32264 64704
rect 31944 63616 31952 63680
rect 32016 63616 32032 63680
rect 32096 63616 32112 63680
rect 32176 63616 32192 63680
rect 32256 63616 32264 63680
rect 31944 63294 32264 63616
rect 31944 63058 31986 63294
rect 32222 63058 32264 63294
rect 31944 62592 32264 63058
rect 31944 62528 31952 62592
rect 32016 62528 32032 62592
rect 32096 62528 32112 62592
rect 32176 62528 32192 62592
rect 32256 62528 32264 62592
rect 31944 61504 32264 62528
rect 31944 61440 31952 61504
rect 32016 61440 32032 61504
rect 32096 61440 32112 61504
rect 32176 61440 32192 61504
rect 32256 61440 32264 61504
rect 31944 60416 32264 61440
rect 31944 60352 31952 60416
rect 32016 60352 32032 60416
rect 32096 60352 32112 60416
rect 32176 60352 32192 60416
rect 32256 60352 32264 60416
rect 31944 59328 32264 60352
rect 31944 59264 31952 59328
rect 32016 59264 32032 59328
rect 32096 59264 32112 59328
rect 32176 59264 32192 59328
rect 32256 59264 32264 59328
rect 31944 58294 32264 59264
rect 31944 58240 31986 58294
rect 32222 58240 32264 58294
rect 31944 58176 31952 58240
rect 32256 58176 32264 58240
rect 31944 58058 31986 58176
rect 32222 58058 32264 58176
rect 31944 57152 32264 58058
rect 31944 57088 31952 57152
rect 32016 57088 32032 57152
rect 32096 57088 32112 57152
rect 32176 57088 32192 57152
rect 32256 57088 32264 57152
rect 31944 56064 32264 57088
rect 31944 56000 31952 56064
rect 32016 56000 32032 56064
rect 32096 56000 32112 56064
rect 32176 56000 32192 56064
rect 32256 56000 32264 56064
rect 31944 54976 32264 56000
rect 31944 54912 31952 54976
rect 32016 54912 32032 54976
rect 32096 54912 32112 54976
rect 32176 54912 32192 54976
rect 32256 54912 32264 54976
rect 31944 53888 32264 54912
rect 31944 53824 31952 53888
rect 32016 53824 32032 53888
rect 32096 53824 32112 53888
rect 32176 53824 32192 53888
rect 32256 53824 32264 53888
rect 31944 53294 32264 53824
rect 31944 53058 31986 53294
rect 32222 53058 32264 53294
rect 31944 52800 32264 53058
rect 31944 52736 31952 52800
rect 32016 52736 32032 52800
rect 32096 52736 32112 52800
rect 32176 52736 32192 52800
rect 32256 52736 32264 52800
rect 31944 51712 32264 52736
rect 31944 51648 31952 51712
rect 32016 51648 32032 51712
rect 32096 51648 32112 51712
rect 32176 51648 32192 51712
rect 32256 51648 32264 51712
rect 31944 50624 32264 51648
rect 31944 50560 31952 50624
rect 32016 50560 32032 50624
rect 32096 50560 32112 50624
rect 32176 50560 32192 50624
rect 32256 50560 32264 50624
rect 31944 49536 32264 50560
rect 31944 49472 31952 49536
rect 32016 49472 32032 49536
rect 32096 49472 32112 49536
rect 32176 49472 32192 49536
rect 32256 49472 32264 49536
rect 31944 48448 32264 49472
rect 31944 48384 31952 48448
rect 32016 48384 32032 48448
rect 32096 48384 32112 48448
rect 32176 48384 32192 48448
rect 32256 48384 32264 48448
rect 31944 48294 32264 48384
rect 31944 48058 31986 48294
rect 32222 48058 32264 48294
rect 31944 47360 32264 48058
rect 31944 47296 31952 47360
rect 32016 47296 32032 47360
rect 32096 47296 32112 47360
rect 32176 47296 32192 47360
rect 32256 47296 32264 47360
rect 31944 46272 32264 47296
rect 31944 46208 31952 46272
rect 32016 46208 32032 46272
rect 32096 46208 32112 46272
rect 32176 46208 32192 46272
rect 32256 46208 32264 46272
rect 31944 45184 32264 46208
rect 31944 45120 31952 45184
rect 32016 45120 32032 45184
rect 32096 45120 32112 45184
rect 32176 45120 32192 45184
rect 32256 45120 32264 45184
rect 31944 44096 32264 45120
rect 31944 44032 31952 44096
rect 32016 44032 32032 44096
rect 32096 44032 32112 44096
rect 32176 44032 32192 44096
rect 32256 44032 32264 44096
rect 31944 43294 32264 44032
rect 31944 43058 31986 43294
rect 32222 43058 32264 43294
rect 31944 43008 32264 43058
rect 31944 42944 31952 43008
rect 32016 42944 32032 43008
rect 32096 42944 32112 43008
rect 32176 42944 32192 43008
rect 32256 42944 32264 43008
rect 31944 41920 32264 42944
rect 31944 41856 31952 41920
rect 32016 41856 32032 41920
rect 32096 41856 32112 41920
rect 32176 41856 32192 41920
rect 32256 41856 32264 41920
rect 31944 40832 32264 41856
rect 31944 40768 31952 40832
rect 32016 40768 32032 40832
rect 32096 40768 32112 40832
rect 32176 40768 32192 40832
rect 32256 40768 32264 40832
rect 30603 40084 30669 40085
rect 30603 40020 30604 40084
rect 30668 40020 30669 40084
rect 30603 40019 30669 40020
rect 27604 39136 27612 39200
rect 27676 39136 27692 39200
rect 27756 39136 27772 39200
rect 27836 39136 27852 39200
rect 27916 39136 27924 39200
rect 27604 38954 27924 39136
rect 27604 38718 27646 38954
rect 27882 38718 27924 38954
rect 27604 38112 27924 38718
rect 27604 38048 27612 38112
rect 27676 38048 27692 38112
rect 27756 38048 27772 38112
rect 27836 38048 27852 38112
rect 27916 38048 27924 38112
rect 27604 37024 27924 38048
rect 27604 36960 27612 37024
rect 27676 36960 27692 37024
rect 27756 36960 27772 37024
rect 27836 36960 27852 37024
rect 27916 36960 27924 37024
rect 27604 35936 27924 36960
rect 27604 35872 27612 35936
rect 27676 35872 27692 35936
rect 27756 35872 27772 35936
rect 27836 35872 27852 35936
rect 27916 35872 27924 35936
rect 27604 34848 27924 35872
rect 27604 34784 27612 34848
rect 27676 34784 27692 34848
rect 27756 34784 27772 34848
rect 27836 34784 27852 34848
rect 27916 34784 27924 34848
rect 27604 33954 27924 34784
rect 27604 33760 27646 33954
rect 27882 33760 27924 33954
rect 27604 33696 27612 33760
rect 27676 33696 27692 33718
rect 27756 33696 27772 33718
rect 27836 33696 27852 33718
rect 27916 33696 27924 33760
rect 27604 32672 27924 33696
rect 27604 32608 27612 32672
rect 27676 32608 27692 32672
rect 27756 32608 27772 32672
rect 27836 32608 27852 32672
rect 27916 32608 27924 32672
rect 27604 31584 27924 32608
rect 27604 31520 27612 31584
rect 27676 31520 27692 31584
rect 27756 31520 27772 31584
rect 27836 31520 27852 31584
rect 27916 31520 27924 31584
rect 27604 30496 27924 31520
rect 30606 31245 30666 40019
rect 31944 39744 32264 40768
rect 31944 39680 31952 39744
rect 32016 39680 32032 39744
rect 32096 39680 32112 39744
rect 32176 39680 32192 39744
rect 32256 39680 32264 39744
rect 31944 38656 32264 39680
rect 31944 38592 31952 38656
rect 32016 38592 32032 38656
rect 32096 38592 32112 38656
rect 32176 38592 32192 38656
rect 32256 38592 32264 38656
rect 31944 38294 32264 38592
rect 31944 38058 31986 38294
rect 32222 38058 32264 38294
rect 31944 37568 32264 38058
rect 31944 37504 31952 37568
rect 32016 37504 32032 37568
rect 32096 37504 32112 37568
rect 32176 37504 32192 37568
rect 32256 37504 32264 37568
rect 31944 36480 32264 37504
rect 31944 36416 31952 36480
rect 32016 36416 32032 36480
rect 32096 36416 32112 36480
rect 32176 36416 32192 36480
rect 32256 36416 32264 36480
rect 31944 35392 32264 36416
rect 31944 35328 31952 35392
rect 32016 35328 32032 35392
rect 32096 35328 32112 35392
rect 32176 35328 32192 35392
rect 32256 35328 32264 35392
rect 31944 34304 32264 35328
rect 31944 34240 31952 34304
rect 32016 34240 32032 34304
rect 32096 34240 32112 34304
rect 32176 34240 32192 34304
rect 32256 34240 32264 34304
rect 31944 33294 32264 34240
rect 31944 33216 31986 33294
rect 32222 33216 32264 33294
rect 31944 33152 31952 33216
rect 32256 33152 32264 33216
rect 31944 33058 31986 33152
rect 32222 33058 32264 33152
rect 31944 32128 32264 33058
rect 31944 32064 31952 32128
rect 32016 32064 32032 32128
rect 32096 32064 32112 32128
rect 32176 32064 32192 32128
rect 32256 32064 32264 32128
rect 30603 31244 30669 31245
rect 30603 31180 30604 31244
rect 30668 31180 30669 31244
rect 30603 31179 30669 31180
rect 27604 30432 27612 30496
rect 27676 30432 27692 30496
rect 27756 30432 27772 30496
rect 27836 30432 27852 30496
rect 27916 30432 27924 30496
rect 27604 29408 27924 30432
rect 27604 29344 27612 29408
rect 27676 29344 27692 29408
rect 27756 29344 27772 29408
rect 27836 29344 27852 29408
rect 27916 29344 27924 29408
rect 27604 28954 27924 29344
rect 27604 28718 27646 28954
rect 27882 28718 27924 28954
rect 27604 28320 27924 28718
rect 27604 28256 27612 28320
rect 27676 28256 27692 28320
rect 27756 28256 27772 28320
rect 27836 28256 27852 28320
rect 27916 28256 27924 28320
rect 27604 27232 27924 28256
rect 27604 27168 27612 27232
rect 27676 27168 27692 27232
rect 27756 27168 27772 27232
rect 27836 27168 27852 27232
rect 27916 27168 27924 27232
rect 27604 26144 27924 27168
rect 27604 26080 27612 26144
rect 27676 26080 27692 26144
rect 27756 26080 27772 26144
rect 27836 26080 27852 26144
rect 27916 26080 27924 26144
rect 27604 25056 27924 26080
rect 27604 24992 27612 25056
rect 27676 24992 27692 25056
rect 27756 24992 27772 25056
rect 27836 24992 27852 25056
rect 27916 24992 27924 25056
rect 27604 23968 27924 24992
rect 27604 23904 27612 23968
rect 27676 23954 27692 23968
rect 27756 23954 27772 23968
rect 27836 23954 27852 23968
rect 27916 23904 27924 23968
rect 27604 23718 27646 23904
rect 27882 23718 27924 23904
rect 27604 22880 27924 23718
rect 27604 22816 27612 22880
rect 27676 22816 27692 22880
rect 27756 22816 27772 22880
rect 27836 22816 27852 22880
rect 27916 22816 27924 22880
rect 27604 21792 27924 22816
rect 27604 21728 27612 21792
rect 27676 21728 27692 21792
rect 27756 21728 27772 21792
rect 27836 21728 27852 21792
rect 27916 21728 27924 21792
rect 27604 20704 27924 21728
rect 27604 20640 27612 20704
rect 27676 20640 27692 20704
rect 27756 20640 27772 20704
rect 27836 20640 27852 20704
rect 27916 20640 27924 20704
rect 27604 19616 27924 20640
rect 27604 19552 27612 19616
rect 27676 19552 27692 19616
rect 27756 19552 27772 19616
rect 27836 19552 27852 19616
rect 27916 19552 27924 19616
rect 27604 18954 27924 19552
rect 27604 18718 27646 18954
rect 27882 18718 27924 18954
rect 27604 18528 27924 18718
rect 27604 18464 27612 18528
rect 27676 18464 27692 18528
rect 27756 18464 27772 18528
rect 27836 18464 27852 18528
rect 27916 18464 27924 18528
rect 27604 17440 27924 18464
rect 27604 17376 27612 17440
rect 27676 17376 27692 17440
rect 27756 17376 27772 17440
rect 27836 17376 27852 17440
rect 27916 17376 27924 17440
rect 27604 16352 27924 17376
rect 27604 16288 27612 16352
rect 27676 16288 27692 16352
rect 27756 16288 27772 16352
rect 27836 16288 27852 16352
rect 27916 16288 27924 16352
rect 27604 15264 27924 16288
rect 27604 15200 27612 15264
rect 27676 15200 27692 15264
rect 27756 15200 27772 15264
rect 27836 15200 27852 15264
rect 27916 15200 27924 15264
rect 27604 14176 27924 15200
rect 27604 14112 27612 14176
rect 27676 14112 27692 14176
rect 27756 14112 27772 14176
rect 27836 14112 27852 14176
rect 27916 14112 27924 14176
rect 27604 13954 27924 14112
rect 27604 13718 27646 13954
rect 27882 13718 27924 13954
rect 27604 13088 27924 13718
rect 27604 13024 27612 13088
rect 27676 13024 27692 13088
rect 27756 13024 27772 13088
rect 27836 13024 27852 13088
rect 27916 13024 27924 13088
rect 27604 12000 27924 13024
rect 27604 11936 27612 12000
rect 27676 11936 27692 12000
rect 27756 11936 27772 12000
rect 27836 11936 27852 12000
rect 27916 11936 27924 12000
rect 27604 10912 27924 11936
rect 27604 10848 27612 10912
rect 27676 10848 27692 10912
rect 27756 10848 27772 10912
rect 27836 10848 27852 10912
rect 27916 10848 27924 10912
rect 27604 9824 27924 10848
rect 27604 9760 27612 9824
rect 27676 9760 27692 9824
rect 27756 9760 27772 9824
rect 27836 9760 27852 9824
rect 27916 9760 27924 9824
rect 27604 8954 27924 9760
rect 27604 8736 27646 8954
rect 27882 8736 27924 8954
rect 27604 8672 27612 8736
rect 27676 8672 27692 8718
rect 27756 8672 27772 8718
rect 27836 8672 27852 8718
rect 27916 8672 27924 8736
rect 27604 7648 27924 8672
rect 27604 7584 27612 7648
rect 27676 7584 27692 7648
rect 27756 7584 27772 7648
rect 27836 7584 27852 7648
rect 27916 7584 27924 7648
rect 27604 6560 27924 7584
rect 27604 6496 27612 6560
rect 27676 6496 27692 6560
rect 27756 6496 27772 6560
rect 27836 6496 27852 6560
rect 27916 6496 27924 6560
rect 27604 5472 27924 6496
rect 27604 5408 27612 5472
rect 27676 5408 27692 5472
rect 27756 5408 27772 5472
rect 27836 5408 27852 5472
rect 27916 5408 27924 5472
rect 27604 4384 27924 5408
rect 27604 4320 27612 4384
rect 27676 4320 27692 4384
rect 27756 4320 27772 4384
rect 27836 4320 27852 4384
rect 27916 4320 27924 4384
rect 27604 3954 27924 4320
rect 27604 3718 27646 3954
rect 27882 3718 27924 3954
rect 27604 3296 27924 3718
rect 27604 3232 27612 3296
rect 27676 3232 27692 3296
rect 27756 3232 27772 3296
rect 27836 3232 27852 3296
rect 27916 3232 27924 3296
rect 27604 2208 27924 3232
rect 27604 2144 27612 2208
rect 27676 2144 27692 2208
rect 27756 2144 27772 2208
rect 27836 2144 27852 2208
rect 27916 2144 27924 2208
rect 27604 2128 27924 2144
rect 31944 31040 32264 32064
rect 31944 30976 31952 31040
rect 32016 30976 32032 31040
rect 32096 30976 32112 31040
rect 32176 30976 32192 31040
rect 32256 30976 32264 31040
rect 31944 29952 32264 30976
rect 31944 29888 31952 29952
rect 32016 29888 32032 29952
rect 32096 29888 32112 29952
rect 32176 29888 32192 29952
rect 32256 29888 32264 29952
rect 31944 28864 32264 29888
rect 31944 28800 31952 28864
rect 32016 28800 32032 28864
rect 32096 28800 32112 28864
rect 32176 28800 32192 28864
rect 32256 28800 32264 28864
rect 31944 28294 32264 28800
rect 31944 28058 31986 28294
rect 32222 28058 32264 28294
rect 31944 27776 32264 28058
rect 31944 27712 31952 27776
rect 32016 27712 32032 27776
rect 32096 27712 32112 27776
rect 32176 27712 32192 27776
rect 32256 27712 32264 27776
rect 31944 26688 32264 27712
rect 31944 26624 31952 26688
rect 32016 26624 32032 26688
rect 32096 26624 32112 26688
rect 32176 26624 32192 26688
rect 32256 26624 32264 26688
rect 31944 25600 32264 26624
rect 31944 25536 31952 25600
rect 32016 25536 32032 25600
rect 32096 25536 32112 25600
rect 32176 25536 32192 25600
rect 32256 25536 32264 25600
rect 31944 24512 32264 25536
rect 31944 24448 31952 24512
rect 32016 24448 32032 24512
rect 32096 24448 32112 24512
rect 32176 24448 32192 24512
rect 32256 24448 32264 24512
rect 31944 23424 32264 24448
rect 31944 23360 31952 23424
rect 32016 23360 32032 23424
rect 32096 23360 32112 23424
rect 32176 23360 32192 23424
rect 32256 23360 32264 23424
rect 31944 23294 32264 23360
rect 31944 23058 31986 23294
rect 32222 23058 32264 23294
rect 31944 22336 32264 23058
rect 31944 22272 31952 22336
rect 32016 22272 32032 22336
rect 32096 22272 32112 22336
rect 32176 22272 32192 22336
rect 32256 22272 32264 22336
rect 31944 21248 32264 22272
rect 31944 21184 31952 21248
rect 32016 21184 32032 21248
rect 32096 21184 32112 21248
rect 32176 21184 32192 21248
rect 32256 21184 32264 21248
rect 31944 20160 32264 21184
rect 31944 20096 31952 20160
rect 32016 20096 32032 20160
rect 32096 20096 32112 20160
rect 32176 20096 32192 20160
rect 32256 20096 32264 20160
rect 31944 19072 32264 20096
rect 31944 19008 31952 19072
rect 32016 19008 32032 19072
rect 32096 19008 32112 19072
rect 32176 19008 32192 19072
rect 32256 19008 32264 19072
rect 31944 18294 32264 19008
rect 31944 18058 31986 18294
rect 32222 18058 32264 18294
rect 31944 17984 32264 18058
rect 31944 17920 31952 17984
rect 32016 17920 32032 17984
rect 32096 17920 32112 17984
rect 32176 17920 32192 17984
rect 32256 17920 32264 17984
rect 31944 16896 32264 17920
rect 31944 16832 31952 16896
rect 32016 16832 32032 16896
rect 32096 16832 32112 16896
rect 32176 16832 32192 16896
rect 32256 16832 32264 16896
rect 31944 15808 32264 16832
rect 31944 15744 31952 15808
rect 32016 15744 32032 15808
rect 32096 15744 32112 15808
rect 32176 15744 32192 15808
rect 32256 15744 32264 15808
rect 31944 14720 32264 15744
rect 31944 14656 31952 14720
rect 32016 14656 32032 14720
rect 32096 14656 32112 14720
rect 32176 14656 32192 14720
rect 32256 14656 32264 14720
rect 31944 13632 32264 14656
rect 31944 13568 31952 13632
rect 32016 13568 32032 13632
rect 32096 13568 32112 13632
rect 32176 13568 32192 13632
rect 32256 13568 32264 13632
rect 31944 13294 32264 13568
rect 31944 13058 31986 13294
rect 32222 13058 32264 13294
rect 31944 12544 32264 13058
rect 31944 12480 31952 12544
rect 32016 12480 32032 12544
rect 32096 12480 32112 12544
rect 32176 12480 32192 12544
rect 32256 12480 32264 12544
rect 31944 11456 32264 12480
rect 31944 11392 31952 11456
rect 32016 11392 32032 11456
rect 32096 11392 32112 11456
rect 32176 11392 32192 11456
rect 32256 11392 32264 11456
rect 31944 10368 32264 11392
rect 31944 10304 31952 10368
rect 32016 10304 32032 10368
rect 32096 10304 32112 10368
rect 32176 10304 32192 10368
rect 32256 10304 32264 10368
rect 31944 9280 32264 10304
rect 31944 9216 31952 9280
rect 32016 9216 32032 9280
rect 32096 9216 32112 9280
rect 32176 9216 32192 9280
rect 32256 9216 32264 9280
rect 31944 8294 32264 9216
rect 31944 8192 31986 8294
rect 32222 8192 32264 8294
rect 31944 8128 31952 8192
rect 32256 8128 32264 8192
rect 31944 8058 31986 8128
rect 32222 8058 32264 8128
rect 31944 7104 32264 8058
rect 31944 7040 31952 7104
rect 32016 7040 32032 7104
rect 32096 7040 32112 7104
rect 32176 7040 32192 7104
rect 32256 7040 32264 7104
rect 31944 6016 32264 7040
rect 31944 5952 31952 6016
rect 32016 5952 32032 6016
rect 32096 5952 32112 6016
rect 32176 5952 32192 6016
rect 32256 5952 32264 6016
rect 31944 4928 32264 5952
rect 31944 4864 31952 4928
rect 32016 4864 32032 4928
rect 32096 4864 32112 4928
rect 32176 4864 32192 4928
rect 32256 4864 32264 4928
rect 31944 3840 32264 4864
rect 31944 3776 31952 3840
rect 32016 3776 32032 3840
rect 32096 3776 32112 3840
rect 32176 3776 32192 3840
rect 32256 3776 32264 3840
rect 31944 3294 32264 3776
rect 31944 3058 31986 3294
rect 32222 3058 32264 3294
rect 31944 2752 32264 3058
rect 31944 2688 31952 2752
rect 32016 2688 32032 2752
rect 32096 2688 32112 2752
rect 32176 2688 32192 2752
rect 32256 2688 32264 2752
rect 31944 2128 32264 2688
rect 32604 69664 32924 69680
rect 32604 69600 32612 69664
rect 32676 69600 32692 69664
rect 32756 69600 32772 69664
rect 32836 69600 32852 69664
rect 32916 69600 32924 69664
rect 32604 68954 32924 69600
rect 32604 68718 32646 68954
rect 32882 68718 32924 68954
rect 32604 68576 32924 68718
rect 32604 68512 32612 68576
rect 32676 68512 32692 68576
rect 32756 68512 32772 68576
rect 32836 68512 32852 68576
rect 32916 68512 32924 68576
rect 32604 67488 32924 68512
rect 32604 67424 32612 67488
rect 32676 67424 32692 67488
rect 32756 67424 32772 67488
rect 32836 67424 32852 67488
rect 32916 67424 32924 67488
rect 32604 66400 32924 67424
rect 32604 66336 32612 66400
rect 32676 66336 32692 66400
rect 32756 66336 32772 66400
rect 32836 66336 32852 66400
rect 32916 66336 32924 66400
rect 32604 65312 32924 66336
rect 32604 65248 32612 65312
rect 32676 65248 32692 65312
rect 32756 65248 32772 65312
rect 32836 65248 32852 65312
rect 32916 65248 32924 65312
rect 32604 64224 32924 65248
rect 32604 64160 32612 64224
rect 32676 64160 32692 64224
rect 32756 64160 32772 64224
rect 32836 64160 32852 64224
rect 32916 64160 32924 64224
rect 32604 63954 32924 64160
rect 32604 63718 32646 63954
rect 32882 63718 32924 63954
rect 32604 63136 32924 63718
rect 32604 63072 32612 63136
rect 32676 63072 32692 63136
rect 32756 63072 32772 63136
rect 32836 63072 32852 63136
rect 32916 63072 32924 63136
rect 32604 62048 32924 63072
rect 32604 61984 32612 62048
rect 32676 61984 32692 62048
rect 32756 61984 32772 62048
rect 32836 61984 32852 62048
rect 32916 61984 32924 62048
rect 32604 60960 32924 61984
rect 32604 60896 32612 60960
rect 32676 60896 32692 60960
rect 32756 60896 32772 60960
rect 32836 60896 32852 60960
rect 32916 60896 32924 60960
rect 32604 59872 32924 60896
rect 32604 59808 32612 59872
rect 32676 59808 32692 59872
rect 32756 59808 32772 59872
rect 32836 59808 32852 59872
rect 32916 59808 32924 59872
rect 32604 58954 32924 59808
rect 32604 58784 32646 58954
rect 32882 58784 32924 58954
rect 32604 58720 32612 58784
rect 32916 58720 32924 58784
rect 32604 58718 32646 58720
rect 32882 58718 32924 58720
rect 32604 57696 32924 58718
rect 32604 57632 32612 57696
rect 32676 57632 32692 57696
rect 32756 57632 32772 57696
rect 32836 57632 32852 57696
rect 32916 57632 32924 57696
rect 32604 56608 32924 57632
rect 32604 56544 32612 56608
rect 32676 56544 32692 56608
rect 32756 56544 32772 56608
rect 32836 56544 32852 56608
rect 32916 56544 32924 56608
rect 32604 55520 32924 56544
rect 32604 55456 32612 55520
rect 32676 55456 32692 55520
rect 32756 55456 32772 55520
rect 32836 55456 32852 55520
rect 32916 55456 32924 55520
rect 32604 54432 32924 55456
rect 32604 54368 32612 54432
rect 32676 54368 32692 54432
rect 32756 54368 32772 54432
rect 32836 54368 32852 54432
rect 32916 54368 32924 54432
rect 32604 53954 32924 54368
rect 32604 53718 32646 53954
rect 32882 53718 32924 53954
rect 32604 53344 32924 53718
rect 32604 53280 32612 53344
rect 32676 53280 32692 53344
rect 32756 53280 32772 53344
rect 32836 53280 32852 53344
rect 32916 53280 32924 53344
rect 32604 52256 32924 53280
rect 32604 52192 32612 52256
rect 32676 52192 32692 52256
rect 32756 52192 32772 52256
rect 32836 52192 32852 52256
rect 32916 52192 32924 52256
rect 32604 51168 32924 52192
rect 32604 51104 32612 51168
rect 32676 51104 32692 51168
rect 32756 51104 32772 51168
rect 32836 51104 32852 51168
rect 32916 51104 32924 51168
rect 32604 50080 32924 51104
rect 36944 69120 37264 69680
rect 36944 69056 36952 69120
rect 37016 69056 37032 69120
rect 37096 69056 37112 69120
rect 37176 69056 37192 69120
rect 37256 69056 37264 69120
rect 36944 68294 37264 69056
rect 36944 68058 36986 68294
rect 37222 68058 37264 68294
rect 36944 68032 37264 68058
rect 36944 67968 36952 68032
rect 37016 67968 37032 68032
rect 37096 67968 37112 68032
rect 37176 67968 37192 68032
rect 37256 67968 37264 68032
rect 36944 66944 37264 67968
rect 36944 66880 36952 66944
rect 37016 66880 37032 66944
rect 37096 66880 37112 66944
rect 37176 66880 37192 66944
rect 37256 66880 37264 66944
rect 36944 65856 37264 66880
rect 36944 65792 36952 65856
rect 37016 65792 37032 65856
rect 37096 65792 37112 65856
rect 37176 65792 37192 65856
rect 37256 65792 37264 65856
rect 36944 64768 37264 65792
rect 36944 64704 36952 64768
rect 37016 64704 37032 64768
rect 37096 64704 37112 64768
rect 37176 64704 37192 64768
rect 37256 64704 37264 64768
rect 36944 63680 37264 64704
rect 36944 63616 36952 63680
rect 37016 63616 37032 63680
rect 37096 63616 37112 63680
rect 37176 63616 37192 63680
rect 37256 63616 37264 63680
rect 36944 63294 37264 63616
rect 36944 63058 36986 63294
rect 37222 63058 37264 63294
rect 36944 62592 37264 63058
rect 36944 62528 36952 62592
rect 37016 62528 37032 62592
rect 37096 62528 37112 62592
rect 37176 62528 37192 62592
rect 37256 62528 37264 62592
rect 36944 61504 37264 62528
rect 36944 61440 36952 61504
rect 37016 61440 37032 61504
rect 37096 61440 37112 61504
rect 37176 61440 37192 61504
rect 37256 61440 37264 61504
rect 36944 60416 37264 61440
rect 36944 60352 36952 60416
rect 37016 60352 37032 60416
rect 37096 60352 37112 60416
rect 37176 60352 37192 60416
rect 37256 60352 37264 60416
rect 36944 59328 37264 60352
rect 36944 59264 36952 59328
rect 37016 59264 37032 59328
rect 37096 59264 37112 59328
rect 37176 59264 37192 59328
rect 37256 59264 37264 59328
rect 36944 58294 37264 59264
rect 36944 58240 36986 58294
rect 37222 58240 37264 58294
rect 36944 58176 36952 58240
rect 37256 58176 37264 58240
rect 36944 58058 36986 58176
rect 37222 58058 37264 58176
rect 36944 57152 37264 58058
rect 36944 57088 36952 57152
rect 37016 57088 37032 57152
rect 37096 57088 37112 57152
rect 37176 57088 37192 57152
rect 37256 57088 37264 57152
rect 36944 56064 37264 57088
rect 36944 56000 36952 56064
rect 37016 56000 37032 56064
rect 37096 56000 37112 56064
rect 37176 56000 37192 56064
rect 37256 56000 37264 56064
rect 36944 54976 37264 56000
rect 36944 54912 36952 54976
rect 37016 54912 37032 54976
rect 37096 54912 37112 54976
rect 37176 54912 37192 54976
rect 37256 54912 37264 54976
rect 36944 53888 37264 54912
rect 36944 53824 36952 53888
rect 37016 53824 37032 53888
rect 37096 53824 37112 53888
rect 37176 53824 37192 53888
rect 37256 53824 37264 53888
rect 36944 53294 37264 53824
rect 36944 53058 36986 53294
rect 37222 53058 37264 53294
rect 36944 52800 37264 53058
rect 36944 52736 36952 52800
rect 37016 52736 37032 52800
rect 37096 52736 37112 52800
rect 37176 52736 37192 52800
rect 37256 52736 37264 52800
rect 36944 51712 37264 52736
rect 36944 51648 36952 51712
rect 37016 51648 37032 51712
rect 37096 51648 37112 51712
rect 37176 51648 37192 51712
rect 37256 51648 37264 51712
rect 34835 51100 34901 51101
rect 34835 51036 34836 51100
rect 34900 51036 34901 51100
rect 34835 51035 34901 51036
rect 32604 50016 32612 50080
rect 32676 50016 32692 50080
rect 32756 50016 32772 50080
rect 32836 50016 32852 50080
rect 32916 50016 32924 50080
rect 32604 48992 32924 50016
rect 32604 48928 32612 48992
rect 32676 48954 32692 48992
rect 32756 48954 32772 48992
rect 32836 48954 32852 48992
rect 32916 48928 32924 48992
rect 32604 48718 32646 48928
rect 32882 48718 32924 48928
rect 32604 47904 32924 48718
rect 32604 47840 32612 47904
rect 32676 47840 32692 47904
rect 32756 47840 32772 47904
rect 32836 47840 32852 47904
rect 32916 47840 32924 47904
rect 32604 46816 32924 47840
rect 32604 46752 32612 46816
rect 32676 46752 32692 46816
rect 32756 46752 32772 46816
rect 32836 46752 32852 46816
rect 32916 46752 32924 46816
rect 32604 45728 32924 46752
rect 32604 45664 32612 45728
rect 32676 45664 32692 45728
rect 32756 45664 32772 45728
rect 32836 45664 32852 45728
rect 32916 45664 32924 45728
rect 32604 44640 32924 45664
rect 32604 44576 32612 44640
rect 32676 44576 32692 44640
rect 32756 44576 32772 44640
rect 32836 44576 32852 44640
rect 32916 44576 32924 44640
rect 32604 43954 32924 44576
rect 32604 43718 32646 43954
rect 32882 43718 32924 43954
rect 32604 43552 32924 43718
rect 32604 43488 32612 43552
rect 32676 43488 32692 43552
rect 32756 43488 32772 43552
rect 32836 43488 32852 43552
rect 32916 43488 32924 43552
rect 32604 42464 32924 43488
rect 32604 42400 32612 42464
rect 32676 42400 32692 42464
rect 32756 42400 32772 42464
rect 32836 42400 32852 42464
rect 32916 42400 32924 42464
rect 32604 41376 32924 42400
rect 32604 41312 32612 41376
rect 32676 41312 32692 41376
rect 32756 41312 32772 41376
rect 32836 41312 32852 41376
rect 32916 41312 32924 41376
rect 32604 40288 32924 41312
rect 32604 40224 32612 40288
rect 32676 40224 32692 40288
rect 32756 40224 32772 40288
rect 32836 40224 32852 40288
rect 32916 40224 32924 40288
rect 32604 39200 32924 40224
rect 32604 39136 32612 39200
rect 32676 39136 32692 39200
rect 32756 39136 32772 39200
rect 32836 39136 32852 39200
rect 32916 39136 32924 39200
rect 32604 38954 32924 39136
rect 32604 38718 32646 38954
rect 32882 38718 32924 38954
rect 32604 38112 32924 38718
rect 32604 38048 32612 38112
rect 32676 38048 32692 38112
rect 32756 38048 32772 38112
rect 32836 38048 32852 38112
rect 32916 38048 32924 38112
rect 32604 37024 32924 38048
rect 32604 36960 32612 37024
rect 32676 36960 32692 37024
rect 32756 36960 32772 37024
rect 32836 36960 32852 37024
rect 32916 36960 32924 37024
rect 32604 35936 32924 36960
rect 32604 35872 32612 35936
rect 32676 35872 32692 35936
rect 32756 35872 32772 35936
rect 32836 35872 32852 35936
rect 32916 35872 32924 35936
rect 32604 34848 32924 35872
rect 32604 34784 32612 34848
rect 32676 34784 32692 34848
rect 32756 34784 32772 34848
rect 32836 34784 32852 34848
rect 32916 34784 32924 34848
rect 32604 33954 32924 34784
rect 32604 33760 32646 33954
rect 32882 33760 32924 33954
rect 32604 33696 32612 33760
rect 32676 33696 32692 33718
rect 32756 33696 32772 33718
rect 32836 33696 32852 33718
rect 32916 33696 32924 33760
rect 32604 32672 32924 33696
rect 32604 32608 32612 32672
rect 32676 32608 32692 32672
rect 32756 32608 32772 32672
rect 32836 32608 32852 32672
rect 32916 32608 32924 32672
rect 32604 31584 32924 32608
rect 32604 31520 32612 31584
rect 32676 31520 32692 31584
rect 32756 31520 32772 31584
rect 32836 31520 32852 31584
rect 32916 31520 32924 31584
rect 32604 30496 32924 31520
rect 32604 30432 32612 30496
rect 32676 30432 32692 30496
rect 32756 30432 32772 30496
rect 32836 30432 32852 30496
rect 32916 30432 32924 30496
rect 32604 29408 32924 30432
rect 32604 29344 32612 29408
rect 32676 29344 32692 29408
rect 32756 29344 32772 29408
rect 32836 29344 32852 29408
rect 32916 29344 32924 29408
rect 32604 28954 32924 29344
rect 32604 28718 32646 28954
rect 32882 28718 32924 28954
rect 32604 28320 32924 28718
rect 32604 28256 32612 28320
rect 32676 28256 32692 28320
rect 32756 28256 32772 28320
rect 32836 28256 32852 28320
rect 32916 28256 32924 28320
rect 32604 27232 32924 28256
rect 32604 27168 32612 27232
rect 32676 27168 32692 27232
rect 32756 27168 32772 27232
rect 32836 27168 32852 27232
rect 32916 27168 32924 27232
rect 32604 26144 32924 27168
rect 32604 26080 32612 26144
rect 32676 26080 32692 26144
rect 32756 26080 32772 26144
rect 32836 26080 32852 26144
rect 32916 26080 32924 26144
rect 32604 25056 32924 26080
rect 32604 24992 32612 25056
rect 32676 24992 32692 25056
rect 32756 24992 32772 25056
rect 32836 24992 32852 25056
rect 32916 24992 32924 25056
rect 32604 23968 32924 24992
rect 32604 23904 32612 23968
rect 32676 23954 32692 23968
rect 32756 23954 32772 23968
rect 32836 23954 32852 23968
rect 32916 23904 32924 23968
rect 32604 23718 32646 23904
rect 32882 23718 32924 23904
rect 32604 22880 32924 23718
rect 32604 22816 32612 22880
rect 32676 22816 32692 22880
rect 32756 22816 32772 22880
rect 32836 22816 32852 22880
rect 32916 22816 32924 22880
rect 32604 21792 32924 22816
rect 32604 21728 32612 21792
rect 32676 21728 32692 21792
rect 32756 21728 32772 21792
rect 32836 21728 32852 21792
rect 32916 21728 32924 21792
rect 32604 20704 32924 21728
rect 32604 20640 32612 20704
rect 32676 20640 32692 20704
rect 32756 20640 32772 20704
rect 32836 20640 32852 20704
rect 32916 20640 32924 20704
rect 32604 19616 32924 20640
rect 32604 19552 32612 19616
rect 32676 19552 32692 19616
rect 32756 19552 32772 19616
rect 32836 19552 32852 19616
rect 32916 19552 32924 19616
rect 32604 18954 32924 19552
rect 32604 18718 32646 18954
rect 32882 18718 32924 18954
rect 32604 18528 32924 18718
rect 32604 18464 32612 18528
rect 32676 18464 32692 18528
rect 32756 18464 32772 18528
rect 32836 18464 32852 18528
rect 32916 18464 32924 18528
rect 32604 17440 32924 18464
rect 32604 17376 32612 17440
rect 32676 17376 32692 17440
rect 32756 17376 32772 17440
rect 32836 17376 32852 17440
rect 32916 17376 32924 17440
rect 32604 16352 32924 17376
rect 32604 16288 32612 16352
rect 32676 16288 32692 16352
rect 32756 16288 32772 16352
rect 32836 16288 32852 16352
rect 32916 16288 32924 16352
rect 32604 15264 32924 16288
rect 32604 15200 32612 15264
rect 32676 15200 32692 15264
rect 32756 15200 32772 15264
rect 32836 15200 32852 15264
rect 32916 15200 32924 15264
rect 32604 14176 32924 15200
rect 32604 14112 32612 14176
rect 32676 14112 32692 14176
rect 32756 14112 32772 14176
rect 32836 14112 32852 14176
rect 32916 14112 32924 14176
rect 32604 13954 32924 14112
rect 32604 13718 32646 13954
rect 32882 13718 32924 13954
rect 32604 13088 32924 13718
rect 32604 13024 32612 13088
rect 32676 13024 32692 13088
rect 32756 13024 32772 13088
rect 32836 13024 32852 13088
rect 32916 13024 32924 13088
rect 32604 12000 32924 13024
rect 32604 11936 32612 12000
rect 32676 11936 32692 12000
rect 32756 11936 32772 12000
rect 32836 11936 32852 12000
rect 32916 11936 32924 12000
rect 32604 10912 32924 11936
rect 34838 11661 34898 51035
rect 36944 50624 37264 51648
rect 36944 50560 36952 50624
rect 37016 50560 37032 50624
rect 37096 50560 37112 50624
rect 37176 50560 37192 50624
rect 37256 50560 37264 50624
rect 36944 49536 37264 50560
rect 36944 49472 36952 49536
rect 37016 49472 37032 49536
rect 37096 49472 37112 49536
rect 37176 49472 37192 49536
rect 37256 49472 37264 49536
rect 36944 48448 37264 49472
rect 36944 48384 36952 48448
rect 37016 48384 37032 48448
rect 37096 48384 37112 48448
rect 37176 48384 37192 48448
rect 37256 48384 37264 48448
rect 36944 48294 37264 48384
rect 36944 48058 36986 48294
rect 37222 48058 37264 48294
rect 36944 47360 37264 48058
rect 36944 47296 36952 47360
rect 37016 47296 37032 47360
rect 37096 47296 37112 47360
rect 37176 47296 37192 47360
rect 37256 47296 37264 47360
rect 36944 46272 37264 47296
rect 36944 46208 36952 46272
rect 37016 46208 37032 46272
rect 37096 46208 37112 46272
rect 37176 46208 37192 46272
rect 37256 46208 37264 46272
rect 36944 45184 37264 46208
rect 36944 45120 36952 45184
rect 37016 45120 37032 45184
rect 37096 45120 37112 45184
rect 37176 45120 37192 45184
rect 37256 45120 37264 45184
rect 36944 44096 37264 45120
rect 36944 44032 36952 44096
rect 37016 44032 37032 44096
rect 37096 44032 37112 44096
rect 37176 44032 37192 44096
rect 37256 44032 37264 44096
rect 36944 43294 37264 44032
rect 36944 43058 36986 43294
rect 37222 43058 37264 43294
rect 36944 43008 37264 43058
rect 36944 42944 36952 43008
rect 37016 42944 37032 43008
rect 37096 42944 37112 43008
rect 37176 42944 37192 43008
rect 37256 42944 37264 43008
rect 36944 41920 37264 42944
rect 36944 41856 36952 41920
rect 37016 41856 37032 41920
rect 37096 41856 37112 41920
rect 37176 41856 37192 41920
rect 37256 41856 37264 41920
rect 36944 40832 37264 41856
rect 36944 40768 36952 40832
rect 37016 40768 37032 40832
rect 37096 40768 37112 40832
rect 37176 40768 37192 40832
rect 37256 40768 37264 40832
rect 36944 39744 37264 40768
rect 36944 39680 36952 39744
rect 37016 39680 37032 39744
rect 37096 39680 37112 39744
rect 37176 39680 37192 39744
rect 37256 39680 37264 39744
rect 36944 38656 37264 39680
rect 36944 38592 36952 38656
rect 37016 38592 37032 38656
rect 37096 38592 37112 38656
rect 37176 38592 37192 38656
rect 37256 38592 37264 38656
rect 36944 38294 37264 38592
rect 36944 38058 36986 38294
rect 37222 38058 37264 38294
rect 36944 37568 37264 38058
rect 36944 37504 36952 37568
rect 37016 37504 37032 37568
rect 37096 37504 37112 37568
rect 37176 37504 37192 37568
rect 37256 37504 37264 37568
rect 36944 36480 37264 37504
rect 36944 36416 36952 36480
rect 37016 36416 37032 36480
rect 37096 36416 37112 36480
rect 37176 36416 37192 36480
rect 37256 36416 37264 36480
rect 36944 35392 37264 36416
rect 36944 35328 36952 35392
rect 37016 35328 37032 35392
rect 37096 35328 37112 35392
rect 37176 35328 37192 35392
rect 37256 35328 37264 35392
rect 36944 34304 37264 35328
rect 36944 34240 36952 34304
rect 37016 34240 37032 34304
rect 37096 34240 37112 34304
rect 37176 34240 37192 34304
rect 37256 34240 37264 34304
rect 36944 33294 37264 34240
rect 36944 33216 36986 33294
rect 37222 33216 37264 33294
rect 36944 33152 36952 33216
rect 37256 33152 37264 33216
rect 36944 33058 36986 33152
rect 37222 33058 37264 33152
rect 36944 32128 37264 33058
rect 36944 32064 36952 32128
rect 37016 32064 37032 32128
rect 37096 32064 37112 32128
rect 37176 32064 37192 32128
rect 37256 32064 37264 32128
rect 36944 31040 37264 32064
rect 36944 30976 36952 31040
rect 37016 30976 37032 31040
rect 37096 30976 37112 31040
rect 37176 30976 37192 31040
rect 37256 30976 37264 31040
rect 36944 29952 37264 30976
rect 36944 29888 36952 29952
rect 37016 29888 37032 29952
rect 37096 29888 37112 29952
rect 37176 29888 37192 29952
rect 37256 29888 37264 29952
rect 36944 28864 37264 29888
rect 36944 28800 36952 28864
rect 37016 28800 37032 28864
rect 37096 28800 37112 28864
rect 37176 28800 37192 28864
rect 37256 28800 37264 28864
rect 36944 28294 37264 28800
rect 36944 28058 36986 28294
rect 37222 28058 37264 28294
rect 36944 27776 37264 28058
rect 36944 27712 36952 27776
rect 37016 27712 37032 27776
rect 37096 27712 37112 27776
rect 37176 27712 37192 27776
rect 37256 27712 37264 27776
rect 36944 26688 37264 27712
rect 36944 26624 36952 26688
rect 37016 26624 37032 26688
rect 37096 26624 37112 26688
rect 37176 26624 37192 26688
rect 37256 26624 37264 26688
rect 36944 25600 37264 26624
rect 36944 25536 36952 25600
rect 37016 25536 37032 25600
rect 37096 25536 37112 25600
rect 37176 25536 37192 25600
rect 37256 25536 37264 25600
rect 36944 24512 37264 25536
rect 36944 24448 36952 24512
rect 37016 24448 37032 24512
rect 37096 24448 37112 24512
rect 37176 24448 37192 24512
rect 37256 24448 37264 24512
rect 36944 23424 37264 24448
rect 36944 23360 36952 23424
rect 37016 23360 37032 23424
rect 37096 23360 37112 23424
rect 37176 23360 37192 23424
rect 37256 23360 37264 23424
rect 36944 23294 37264 23360
rect 36944 23058 36986 23294
rect 37222 23058 37264 23294
rect 36944 22336 37264 23058
rect 36944 22272 36952 22336
rect 37016 22272 37032 22336
rect 37096 22272 37112 22336
rect 37176 22272 37192 22336
rect 37256 22272 37264 22336
rect 36944 21248 37264 22272
rect 36944 21184 36952 21248
rect 37016 21184 37032 21248
rect 37096 21184 37112 21248
rect 37176 21184 37192 21248
rect 37256 21184 37264 21248
rect 36944 20160 37264 21184
rect 36944 20096 36952 20160
rect 37016 20096 37032 20160
rect 37096 20096 37112 20160
rect 37176 20096 37192 20160
rect 37256 20096 37264 20160
rect 36944 19072 37264 20096
rect 36944 19008 36952 19072
rect 37016 19008 37032 19072
rect 37096 19008 37112 19072
rect 37176 19008 37192 19072
rect 37256 19008 37264 19072
rect 36944 18294 37264 19008
rect 36944 18058 36986 18294
rect 37222 18058 37264 18294
rect 36944 17984 37264 18058
rect 36944 17920 36952 17984
rect 37016 17920 37032 17984
rect 37096 17920 37112 17984
rect 37176 17920 37192 17984
rect 37256 17920 37264 17984
rect 36944 16896 37264 17920
rect 36944 16832 36952 16896
rect 37016 16832 37032 16896
rect 37096 16832 37112 16896
rect 37176 16832 37192 16896
rect 37256 16832 37264 16896
rect 36944 15808 37264 16832
rect 36944 15744 36952 15808
rect 37016 15744 37032 15808
rect 37096 15744 37112 15808
rect 37176 15744 37192 15808
rect 37256 15744 37264 15808
rect 36944 14720 37264 15744
rect 36944 14656 36952 14720
rect 37016 14656 37032 14720
rect 37096 14656 37112 14720
rect 37176 14656 37192 14720
rect 37256 14656 37264 14720
rect 36944 13632 37264 14656
rect 36944 13568 36952 13632
rect 37016 13568 37032 13632
rect 37096 13568 37112 13632
rect 37176 13568 37192 13632
rect 37256 13568 37264 13632
rect 36944 13294 37264 13568
rect 36944 13058 36986 13294
rect 37222 13058 37264 13294
rect 36944 12544 37264 13058
rect 36944 12480 36952 12544
rect 37016 12480 37032 12544
rect 37096 12480 37112 12544
rect 37176 12480 37192 12544
rect 37256 12480 37264 12544
rect 34835 11660 34901 11661
rect 34835 11596 34836 11660
rect 34900 11596 34901 11660
rect 34835 11595 34901 11596
rect 32604 10848 32612 10912
rect 32676 10848 32692 10912
rect 32756 10848 32772 10912
rect 32836 10848 32852 10912
rect 32916 10848 32924 10912
rect 32604 9824 32924 10848
rect 32604 9760 32612 9824
rect 32676 9760 32692 9824
rect 32756 9760 32772 9824
rect 32836 9760 32852 9824
rect 32916 9760 32924 9824
rect 32604 8954 32924 9760
rect 32604 8736 32646 8954
rect 32882 8736 32924 8954
rect 32604 8672 32612 8736
rect 32676 8672 32692 8718
rect 32756 8672 32772 8718
rect 32836 8672 32852 8718
rect 32916 8672 32924 8736
rect 32604 7648 32924 8672
rect 32604 7584 32612 7648
rect 32676 7584 32692 7648
rect 32756 7584 32772 7648
rect 32836 7584 32852 7648
rect 32916 7584 32924 7648
rect 32604 6560 32924 7584
rect 32604 6496 32612 6560
rect 32676 6496 32692 6560
rect 32756 6496 32772 6560
rect 32836 6496 32852 6560
rect 32916 6496 32924 6560
rect 32604 5472 32924 6496
rect 32604 5408 32612 5472
rect 32676 5408 32692 5472
rect 32756 5408 32772 5472
rect 32836 5408 32852 5472
rect 32916 5408 32924 5472
rect 32604 4384 32924 5408
rect 32604 4320 32612 4384
rect 32676 4320 32692 4384
rect 32756 4320 32772 4384
rect 32836 4320 32852 4384
rect 32916 4320 32924 4384
rect 32604 3954 32924 4320
rect 32604 3718 32646 3954
rect 32882 3718 32924 3954
rect 32604 3296 32924 3718
rect 32604 3232 32612 3296
rect 32676 3232 32692 3296
rect 32756 3232 32772 3296
rect 32836 3232 32852 3296
rect 32916 3232 32924 3296
rect 32604 2208 32924 3232
rect 32604 2144 32612 2208
rect 32676 2144 32692 2208
rect 32756 2144 32772 2208
rect 32836 2144 32852 2208
rect 32916 2144 32924 2208
rect 32604 2128 32924 2144
rect 36944 11456 37264 12480
rect 36944 11392 36952 11456
rect 37016 11392 37032 11456
rect 37096 11392 37112 11456
rect 37176 11392 37192 11456
rect 37256 11392 37264 11456
rect 36944 10368 37264 11392
rect 36944 10304 36952 10368
rect 37016 10304 37032 10368
rect 37096 10304 37112 10368
rect 37176 10304 37192 10368
rect 37256 10304 37264 10368
rect 36944 9280 37264 10304
rect 36944 9216 36952 9280
rect 37016 9216 37032 9280
rect 37096 9216 37112 9280
rect 37176 9216 37192 9280
rect 37256 9216 37264 9280
rect 36944 8294 37264 9216
rect 36944 8192 36986 8294
rect 37222 8192 37264 8294
rect 36944 8128 36952 8192
rect 37256 8128 37264 8192
rect 36944 8058 36986 8128
rect 37222 8058 37264 8128
rect 36944 7104 37264 8058
rect 36944 7040 36952 7104
rect 37016 7040 37032 7104
rect 37096 7040 37112 7104
rect 37176 7040 37192 7104
rect 37256 7040 37264 7104
rect 36944 6016 37264 7040
rect 36944 5952 36952 6016
rect 37016 5952 37032 6016
rect 37096 5952 37112 6016
rect 37176 5952 37192 6016
rect 37256 5952 37264 6016
rect 36944 4928 37264 5952
rect 36944 4864 36952 4928
rect 37016 4864 37032 4928
rect 37096 4864 37112 4928
rect 37176 4864 37192 4928
rect 37256 4864 37264 4928
rect 36944 3840 37264 4864
rect 36944 3776 36952 3840
rect 37016 3776 37032 3840
rect 37096 3776 37112 3840
rect 37176 3776 37192 3840
rect 37256 3776 37264 3840
rect 36944 3294 37264 3776
rect 36944 3058 36986 3294
rect 37222 3058 37264 3294
rect 36944 2752 37264 3058
rect 36944 2688 36952 2752
rect 37016 2688 37032 2752
rect 37096 2688 37112 2752
rect 37176 2688 37192 2752
rect 37256 2688 37264 2752
rect 36944 2128 37264 2688
rect 37604 69664 37924 69680
rect 37604 69600 37612 69664
rect 37676 69600 37692 69664
rect 37756 69600 37772 69664
rect 37836 69600 37852 69664
rect 37916 69600 37924 69664
rect 37604 68954 37924 69600
rect 37604 68718 37646 68954
rect 37882 68718 37924 68954
rect 37604 68576 37924 68718
rect 37604 68512 37612 68576
rect 37676 68512 37692 68576
rect 37756 68512 37772 68576
rect 37836 68512 37852 68576
rect 37916 68512 37924 68576
rect 37604 67488 37924 68512
rect 37604 67424 37612 67488
rect 37676 67424 37692 67488
rect 37756 67424 37772 67488
rect 37836 67424 37852 67488
rect 37916 67424 37924 67488
rect 37604 66400 37924 67424
rect 37604 66336 37612 66400
rect 37676 66336 37692 66400
rect 37756 66336 37772 66400
rect 37836 66336 37852 66400
rect 37916 66336 37924 66400
rect 37604 65312 37924 66336
rect 37604 65248 37612 65312
rect 37676 65248 37692 65312
rect 37756 65248 37772 65312
rect 37836 65248 37852 65312
rect 37916 65248 37924 65312
rect 37604 64224 37924 65248
rect 37604 64160 37612 64224
rect 37676 64160 37692 64224
rect 37756 64160 37772 64224
rect 37836 64160 37852 64224
rect 37916 64160 37924 64224
rect 37604 63954 37924 64160
rect 37604 63718 37646 63954
rect 37882 63718 37924 63954
rect 37604 63136 37924 63718
rect 37604 63072 37612 63136
rect 37676 63072 37692 63136
rect 37756 63072 37772 63136
rect 37836 63072 37852 63136
rect 37916 63072 37924 63136
rect 37604 62048 37924 63072
rect 37604 61984 37612 62048
rect 37676 61984 37692 62048
rect 37756 61984 37772 62048
rect 37836 61984 37852 62048
rect 37916 61984 37924 62048
rect 37604 60960 37924 61984
rect 37604 60896 37612 60960
rect 37676 60896 37692 60960
rect 37756 60896 37772 60960
rect 37836 60896 37852 60960
rect 37916 60896 37924 60960
rect 37604 59872 37924 60896
rect 37604 59808 37612 59872
rect 37676 59808 37692 59872
rect 37756 59808 37772 59872
rect 37836 59808 37852 59872
rect 37916 59808 37924 59872
rect 37604 58954 37924 59808
rect 37604 58784 37646 58954
rect 37882 58784 37924 58954
rect 37604 58720 37612 58784
rect 37916 58720 37924 58784
rect 37604 58718 37646 58720
rect 37882 58718 37924 58720
rect 37604 57696 37924 58718
rect 37604 57632 37612 57696
rect 37676 57632 37692 57696
rect 37756 57632 37772 57696
rect 37836 57632 37852 57696
rect 37916 57632 37924 57696
rect 37604 56608 37924 57632
rect 37604 56544 37612 56608
rect 37676 56544 37692 56608
rect 37756 56544 37772 56608
rect 37836 56544 37852 56608
rect 37916 56544 37924 56608
rect 37604 55520 37924 56544
rect 37604 55456 37612 55520
rect 37676 55456 37692 55520
rect 37756 55456 37772 55520
rect 37836 55456 37852 55520
rect 37916 55456 37924 55520
rect 37604 54432 37924 55456
rect 37604 54368 37612 54432
rect 37676 54368 37692 54432
rect 37756 54368 37772 54432
rect 37836 54368 37852 54432
rect 37916 54368 37924 54432
rect 37604 53954 37924 54368
rect 37604 53718 37646 53954
rect 37882 53718 37924 53954
rect 37604 53344 37924 53718
rect 37604 53280 37612 53344
rect 37676 53280 37692 53344
rect 37756 53280 37772 53344
rect 37836 53280 37852 53344
rect 37916 53280 37924 53344
rect 37604 52256 37924 53280
rect 37604 52192 37612 52256
rect 37676 52192 37692 52256
rect 37756 52192 37772 52256
rect 37836 52192 37852 52256
rect 37916 52192 37924 52256
rect 37604 51168 37924 52192
rect 37604 51104 37612 51168
rect 37676 51104 37692 51168
rect 37756 51104 37772 51168
rect 37836 51104 37852 51168
rect 37916 51104 37924 51168
rect 37604 50080 37924 51104
rect 37604 50016 37612 50080
rect 37676 50016 37692 50080
rect 37756 50016 37772 50080
rect 37836 50016 37852 50080
rect 37916 50016 37924 50080
rect 37604 48992 37924 50016
rect 37604 48928 37612 48992
rect 37676 48954 37692 48992
rect 37756 48954 37772 48992
rect 37836 48954 37852 48992
rect 37916 48928 37924 48992
rect 37604 48718 37646 48928
rect 37882 48718 37924 48928
rect 37604 47904 37924 48718
rect 37604 47840 37612 47904
rect 37676 47840 37692 47904
rect 37756 47840 37772 47904
rect 37836 47840 37852 47904
rect 37916 47840 37924 47904
rect 37604 46816 37924 47840
rect 37604 46752 37612 46816
rect 37676 46752 37692 46816
rect 37756 46752 37772 46816
rect 37836 46752 37852 46816
rect 37916 46752 37924 46816
rect 37604 45728 37924 46752
rect 37604 45664 37612 45728
rect 37676 45664 37692 45728
rect 37756 45664 37772 45728
rect 37836 45664 37852 45728
rect 37916 45664 37924 45728
rect 37604 44640 37924 45664
rect 37604 44576 37612 44640
rect 37676 44576 37692 44640
rect 37756 44576 37772 44640
rect 37836 44576 37852 44640
rect 37916 44576 37924 44640
rect 37604 43954 37924 44576
rect 37604 43718 37646 43954
rect 37882 43718 37924 43954
rect 37604 43552 37924 43718
rect 37604 43488 37612 43552
rect 37676 43488 37692 43552
rect 37756 43488 37772 43552
rect 37836 43488 37852 43552
rect 37916 43488 37924 43552
rect 37604 42464 37924 43488
rect 37604 42400 37612 42464
rect 37676 42400 37692 42464
rect 37756 42400 37772 42464
rect 37836 42400 37852 42464
rect 37916 42400 37924 42464
rect 37604 41376 37924 42400
rect 37604 41312 37612 41376
rect 37676 41312 37692 41376
rect 37756 41312 37772 41376
rect 37836 41312 37852 41376
rect 37916 41312 37924 41376
rect 37604 40288 37924 41312
rect 37604 40224 37612 40288
rect 37676 40224 37692 40288
rect 37756 40224 37772 40288
rect 37836 40224 37852 40288
rect 37916 40224 37924 40288
rect 37604 39200 37924 40224
rect 37604 39136 37612 39200
rect 37676 39136 37692 39200
rect 37756 39136 37772 39200
rect 37836 39136 37852 39200
rect 37916 39136 37924 39200
rect 37604 38954 37924 39136
rect 37604 38718 37646 38954
rect 37882 38718 37924 38954
rect 37604 38112 37924 38718
rect 37604 38048 37612 38112
rect 37676 38048 37692 38112
rect 37756 38048 37772 38112
rect 37836 38048 37852 38112
rect 37916 38048 37924 38112
rect 37604 37024 37924 38048
rect 37604 36960 37612 37024
rect 37676 36960 37692 37024
rect 37756 36960 37772 37024
rect 37836 36960 37852 37024
rect 37916 36960 37924 37024
rect 37604 35936 37924 36960
rect 37604 35872 37612 35936
rect 37676 35872 37692 35936
rect 37756 35872 37772 35936
rect 37836 35872 37852 35936
rect 37916 35872 37924 35936
rect 37604 34848 37924 35872
rect 37604 34784 37612 34848
rect 37676 34784 37692 34848
rect 37756 34784 37772 34848
rect 37836 34784 37852 34848
rect 37916 34784 37924 34848
rect 37604 33954 37924 34784
rect 37604 33760 37646 33954
rect 37882 33760 37924 33954
rect 37604 33696 37612 33760
rect 37676 33696 37692 33718
rect 37756 33696 37772 33718
rect 37836 33696 37852 33718
rect 37916 33696 37924 33760
rect 37604 32672 37924 33696
rect 37604 32608 37612 32672
rect 37676 32608 37692 32672
rect 37756 32608 37772 32672
rect 37836 32608 37852 32672
rect 37916 32608 37924 32672
rect 37604 31584 37924 32608
rect 37604 31520 37612 31584
rect 37676 31520 37692 31584
rect 37756 31520 37772 31584
rect 37836 31520 37852 31584
rect 37916 31520 37924 31584
rect 37604 30496 37924 31520
rect 37604 30432 37612 30496
rect 37676 30432 37692 30496
rect 37756 30432 37772 30496
rect 37836 30432 37852 30496
rect 37916 30432 37924 30496
rect 37604 29408 37924 30432
rect 37604 29344 37612 29408
rect 37676 29344 37692 29408
rect 37756 29344 37772 29408
rect 37836 29344 37852 29408
rect 37916 29344 37924 29408
rect 37604 28954 37924 29344
rect 37604 28718 37646 28954
rect 37882 28718 37924 28954
rect 37604 28320 37924 28718
rect 37604 28256 37612 28320
rect 37676 28256 37692 28320
rect 37756 28256 37772 28320
rect 37836 28256 37852 28320
rect 37916 28256 37924 28320
rect 37604 27232 37924 28256
rect 37604 27168 37612 27232
rect 37676 27168 37692 27232
rect 37756 27168 37772 27232
rect 37836 27168 37852 27232
rect 37916 27168 37924 27232
rect 37604 26144 37924 27168
rect 37604 26080 37612 26144
rect 37676 26080 37692 26144
rect 37756 26080 37772 26144
rect 37836 26080 37852 26144
rect 37916 26080 37924 26144
rect 37604 25056 37924 26080
rect 37604 24992 37612 25056
rect 37676 24992 37692 25056
rect 37756 24992 37772 25056
rect 37836 24992 37852 25056
rect 37916 24992 37924 25056
rect 37604 23968 37924 24992
rect 37604 23904 37612 23968
rect 37676 23954 37692 23968
rect 37756 23954 37772 23968
rect 37836 23954 37852 23968
rect 37916 23904 37924 23968
rect 37604 23718 37646 23904
rect 37882 23718 37924 23904
rect 37604 22880 37924 23718
rect 37604 22816 37612 22880
rect 37676 22816 37692 22880
rect 37756 22816 37772 22880
rect 37836 22816 37852 22880
rect 37916 22816 37924 22880
rect 37604 21792 37924 22816
rect 37604 21728 37612 21792
rect 37676 21728 37692 21792
rect 37756 21728 37772 21792
rect 37836 21728 37852 21792
rect 37916 21728 37924 21792
rect 37604 20704 37924 21728
rect 37604 20640 37612 20704
rect 37676 20640 37692 20704
rect 37756 20640 37772 20704
rect 37836 20640 37852 20704
rect 37916 20640 37924 20704
rect 37604 19616 37924 20640
rect 37604 19552 37612 19616
rect 37676 19552 37692 19616
rect 37756 19552 37772 19616
rect 37836 19552 37852 19616
rect 37916 19552 37924 19616
rect 37604 18954 37924 19552
rect 37604 18718 37646 18954
rect 37882 18718 37924 18954
rect 37604 18528 37924 18718
rect 37604 18464 37612 18528
rect 37676 18464 37692 18528
rect 37756 18464 37772 18528
rect 37836 18464 37852 18528
rect 37916 18464 37924 18528
rect 37604 17440 37924 18464
rect 37604 17376 37612 17440
rect 37676 17376 37692 17440
rect 37756 17376 37772 17440
rect 37836 17376 37852 17440
rect 37916 17376 37924 17440
rect 37604 16352 37924 17376
rect 37604 16288 37612 16352
rect 37676 16288 37692 16352
rect 37756 16288 37772 16352
rect 37836 16288 37852 16352
rect 37916 16288 37924 16352
rect 37604 15264 37924 16288
rect 37604 15200 37612 15264
rect 37676 15200 37692 15264
rect 37756 15200 37772 15264
rect 37836 15200 37852 15264
rect 37916 15200 37924 15264
rect 37604 14176 37924 15200
rect 37604 14112 37612 14176
rect 37676 14112 37692 14176
rect 37756 14112 37772 14176
rect 37836 14112 37852 14176
rect 37916 14112 37924 14176
rect 37604 13954 37924 14112
rect 37604 13718 37646 13954
rect 37882 13718 37924 13954
rect 37604 13088 37924 13718
rect 37604 13024 37612 13088
rect 37676 13024 37692 13088
rect 37756 13024 37772 13088
rect 37836 13024 37852 13088
rect 37916 13024 37924 13088
rect 37604 12000 37924 13024
rect 37604 11936 37612 12000
rect 37676 11936 37692 12000
rect 37756 11936 37772 12000
rect 37836 11936 37852 12000
rect 37916 11936 37924 12000
rect 37604 10912 37924 11936
rect 37604 10848 37612 10912
rect 37676 10848 37692 10912
rect 37756 10848 37772 10912
rect 37836 10848 37852 10912
rect 37916 10848 37924 10912
rect 37604 9824 37924 10848
rect 37604 9760 37612 9824
rect 37676 9760 37692 9824
rect 37756 9760 37772 9824
rect 37836 9760 37852 9824
rect 37916 9760 37924 9824
rect 37604 8954 37924 9760
rect 37604 8736 37646 8954
rect 37882 8736 37924 8954
rect 37604 8672 37612 8736
rect 37676 8672 37692 8718
rect 37756 8672 37772 8718
rect 37836 8672 37852 8718
rect 37916 8672 37924 8736
rect 37604 7648 37924 8672
rect 37604 7584 37612 7648
rect 37676 7584 37692 7648
rect 37756 7584 37772 7648
rect 37836 7584 37852 7648
rect 37916 7584 37924 7648
rect 37604 6560 37924 7584
rect 37604 6496 37612 6560
rect 37676 6496 37692 6560
rect 37756 6496 37772 6560
rect 37836 6496 37852 6560
rect 37916 6496 37924 6560
rect 37604 5472 37924 6496
rect 37604 5408 37612 5472
rect 37676 5408 37692 5472
rect 37756 5408 37772 5472
rect 37836 5408 37852 5472
rect 37916 5408 37924 5472
rect 37604 4384 37924 5408
rect 37604 4320 37612 4384
rect 37676 4320 37692 4384
rect 37756 4320 37772 4384
rect 37836 4320 37852 4384
rect 37916 4320 37924 4384
rect 37604 3954 37924 4320
rect 37604 3718 37646 3954
rect 37882 3718 37924 3954
rect 37604 3296 37924 3718
rect 37604 3232 37612 3296
rect 37676 3232 37692 3296
rect 37756 3232 37772 3296
rect 37836 3232 37852 3296
rect 37916 3232 37924 3296
rect 37604 2208 37924 3232
rect 37604 2144 37612 2208
rect 37676 2144 37692 2208
rect 37756 2144 37772 2208
rect 37836 2144 37852 2208
rect 37916 2144 37924 2208
rect 37604 2128 37924 2144
<< via4 >>
rect 1986 68058 2222 68294
rect 1986 63058 2222 63294
rect 1986 58240 2222 58294
rect 1986 58176 2016 58240
rect 2016 58176 2032 58240
rect 2032 58176 2096 58240
rect 2096 58176 2112 58240
rect 2112 58176 2176 58240
rect 2176 58176 2192 58240
rect 2192 58176 2222 58240
rect 1986 58058 2222 58176
rect 1986 53058 2222 53294
rect 1986 48058 2222 48294
rect 1986 43058 2222 43294
rect 1986 38058 2222 38294
rect 1986 33216 2222 33294
rect 1986 33152 2016 33216
rect 2016 33152 2032 33216
rect 2032 33152 2096 33216
rect 2096 33152 2112 33216
rect 2112 33152 2176 33216
rect 2176 33152 2192 33216
rect 2192 33152 2222 33216
rect 1986 33058 2222 33152
rect 1986 28058 2222 28294
rect 1986 23058 2222 23294
rect 1986 18058 2222 18294
rect 1986 13058 2222 13294
rect 1986 8192 2222 8294
rect 1986 8128 2016 8192
rect 2016 8128 2032 8192
rect 2032 8128 2096 8192
rect 2096 8128 2112 8192
rect 2112 8128 2176 8192
rect 2176 8128 2192 8192
rect 2192 8128 2222 8192
rect 1986 8058 2222 8128
rect 1986 3058 2222 3294
rect 2646 68718 2882 68954
rect 6986 68058 7222 68294
rect 2646 63718 2882 63954
rect 2646 58784 2882 58954
rect 2646 58720 2676 58784
rect 2676 58720 2692 58784
rect 2692 58720 2756 58784
rect 2756 58720 2772 58784
rect 2772 58720 2836 58784
rect 2836 58720 2852 58784
rect 2852 58720 2882 58784
rect 2646 58718 2882 58720
rect 2646 53718 2882 53954
rect 2646 48928 2676 48954
rect 2676 48928 2692 48954
rect 2692 48928 2756 48954
rect 2756 48928 2772 48954
rect 2772 48928 2836 48954
rect 2836 48928 2852 48954
rect 2852 48928 2882 48954
rect 2646 48718 2882 48928
rect 2646 43718 2882 43954
rect 2646 38718 2882 38954
rect 2646 33760 2882 33954
rect 2646 33718 2676 33760
rect 2676 33718 2692 33760
rect 2692 33718 2756 33760
rect 2756 33718 2772 33760
rect 2772 33718 2836 33760
rect 2836 33718 2852 33760
rect 2852 33718 2882 33760
rect 2646 28718 2882 28954
rect 2646 23904 2676 23954
rect 2676 23904 2692 23954
rect 2692 23904 2756 23954
rect 2756 23904 2772 23954
rect 2772 23904 2836 23954
rect 2836 23904 2852 23954
rect 2852 23904 2882 23954
rect 2646 23718 2882 23904
rect 2646 18718 2882 18954
rect 2646 13718 2882 13954
rect 6986 63058 7222 63294
rect 6986 58240 7222 58294
rect 6986 58176 7016 58240
rect 7016 58176 7032 58240
rect 7032 58176 7096 58240
rect 7096 58176 7112 58240
rect 7112 58176 7176 58240
rect 7176 58176 7192 58240
rect 7192 58176 7222 58240
rect 6986 58058 7222 58176
rect 6986 53058 7222 53294
rect 6986 48058 7222 48294
rect 6986 43058 7222 43294
rect 6986 38058 7222 38294
rect 6986 33216 7222 33294
rect 6986 33152 7016 33216
rect 7016 33152 7032 33216
rect 7032 33152 7096 33216
rect 7096 33152 7112 33216
rect 7112 33152 7176 33216
rect 7176 33152 7192 33216
rect 7192 33152 7222 33216
rect 6986 33058 7222 33152
rect 6986 28058 7222 28294
rect 6986 23058 7222 23294
rect 6986 18058 7222 18294
rect 6986 13058 7222 13294
rect 2646 8736 2882 8954
rect 2646 8718 2676 8736
rect 2676 8718 2692 8736
rect 2692 8718 2756 8736
rect 2756 8718 2772 8736
rect 2772 8718 2836 8736
rect 2836 8718 2852 8736
rect 2852 8718 2882 8736
rect 2646 3718 2882 3954
rect 6986 8192 7222 8294
rect 6986 8128 7016 8192
rect 7016 8128 7032 8192
rect 7032 8128 7096 8192
rect 7096 8128 7112 8192
rect 7112 8128 7176 8192
rect 7176 8128 7192 8192
rect 7192 8128 7222 8192
rect 6986 8058 7222 8128
rect 6986 3058 7222 3294
rect 7646 68718 7882 68954
rect 7646 63718 7882 63954
rect 7646 58784 7882 58954
rect 7646 58720 7676 58784
rect 7676 58720 7692 58784
rect 7692 58720 7756 58784
rect 7756 58720 7772 58784
rect 7772 58720 7836 58784
rect 7836 58720 7852 58784
rect 7852 58720 7882 58784
rect 7646 58718 7882 58720
rect 7646 53718 7882 53954
rect 7646 48928 7676 48954
rect 7676 48928 7692 48954
rect 7692 48928 7756 48954
rect 7756 48928 7772 48954
rect 7772 48928 7836 48954
rect 7836 48928 7852 48954
rect 7852 48928 7882 48954
rect 7646 48718 7882 48928
rect 7646 43718 7882 43954
rect 7646 38718 7882 38954
rect 7646 33760 7882 33954
rect 7646 33718 7676 33760
rect 7676 33718 7692 33760
rect 7692 33718 7756 33760
rect 7756 33718 7772 33760
rect 7772 33718 7836 33760
rect 7836 33718 7852 33760
rect 7852 33718 7882 33760
rect 7646 28718 7882 28954
rect 7646 23904 7676 23954
rect 7676 23904 7692 23954
rect 7692 23904 7756 23954
rect 7756 23904 7772 23954
rect 7772 23904 7836 23954
rect 7836 23904 7852 23954
rect 7852 23904 7882 23954
rect 7646 23718 7882 23904
rect 7646 18718 7882 18954
rect 7646 13718 7882 13954
rect 7646 8736 7882 8954
rect 7646 8718 7676 8736
rect 7676 8718 7692 8736
rect 7692 8718 7756 8736
rect 7756 8718 7772 8736
rect 7772 8718 7836 8736
rect 7836 8718 7852 8736
rect 7852 8718 7882 8736
rect 7646 3718 7882 3954
rect 11986 68058 12222 68294
rect 11986 63058 12222 63294
rect 11986 58240 12222 58294
rect 11986 58176 12016 58240
rect 12016 58176 12032 58240
rect 12032 58176 12096 58240
rect 12096 58176 12112 58240
rect 12112 58176 12176 58240
rect 12176 58176 12192 58240
rect 12192 58176 12222 58240
rect 11986 58058 12222 58176
rect 11986 53058 12222 53294
rect 11986 48058 12222 48294
rect 11986 43058 12222 43294
rect 11986 38058 12222 38294
rect 11986 33216 12222 33294
rect 11986 33152 12016 33216
rect 12016 33152 12032 33216
rect 12032 33152 12096 33216
rect 12096 33152 12112 33216
rect 12112 33152 12176 33216
rect 12176 33152 12192 33216
rect 12192 33152 12222 33216
rect 11986 33058 12222 33152
rect 11986 28058 12222 28294
rect 11986 23058 12222 23294
rect 11986 18058 12222 18294
rect 11986 13058 12222 13294
rect 11986 8192 12222 8294
rect 11986 8128 12016 8192
rect 12016 8128 12032 8192
rect 12032 8128 12096 8192
rect 12096 8128 12112 8192
rect 12112 8128 12176 8192
rect 12176 8128 12192 8192
rect 12192 8128 12222 8192
rect 11986 8058 12222 8128
rect 11986 3058 12222 3294
rect 12646 68718 12882 68954
rect 16986 68058 17222 68294
rect 12646 63718 12882 63954
rect 12646 58784 12882 58954
rect 12646 58720 12676 58784
rect 12676 58720 12692 58784
rect 12692 58720 12756 58784
rect 12756 58720 12772 58784
rect 12772 58720 12836 58784
rect 12836 58720 12852 58784
rect 12852 58720 12882 58784
rect 12646 58718 12882 58720
rect 12646 53718 12882 53954
rect 12646 48928 12676 48954
rect 12676 48928 12692 48954
rect 12692 48928 12756 48954
rect 12756 48928 12772 48954
rect 12772 48928 12836 48954
rect 12836 48928 12852 48954
rect 12852 48928 12882 48954
rect 12646 48718 12882 48928
rect 12646 43718 12882 43954
rect 12646 38718 12882 38954
rect 12646 33760 12882 33954
rect 12646 33718 12676 33760
rect 12676 33718 12692 33760
rect 12692 33718 12756 33760
rect 12756 33718 12772 33760
rect 12772 33718 12836 33760
rect 12836 33718 12852 33760
rect 12852 33718 12882 33760
rect 12646 28718 12882 28954
rect 12646 23904 12676 23954
rect 12676 23904 12692 23954
rect 12692 23904 12756 23954
rect 12756 23904 12772 23954
rect 12772 23904 12836 23954
rect 12836 23904 12852 23954
rect 12852 23904 12882 23954
rect 12646 23718 12882 23904
rect 16986 63058 17222 63294
rect 16986 58240 17222 58294
rect 16986 58176 17016 58240
rect 17016 58176 17032 58240
rect 17032 58176 17096 58240
rect 17096 58176 17112 58240
rect 17112 58176 17176 58240
rect 17176 58176 17192 58240
rect 17192 58176 17222 58240
rect 16986 58058 17222 58176
rect 12646 18718 12882 18954
rect 12646 13718 12882 13954
rect 12646 8736 12882 8954
rect 12646 8718 12676 8736
rect 12676 8718 12692 8736
rect 12692 8718 12756 8736
rect 12756 8718 12772 8736
rect 12772 8718 12836 8736
rect 12836 8718 12852 8736
rect 12852 8718 12882 8736
rect 12646 3718 12882 3954
rect 16986 53058 17222 53294
rect 16986 48058 17222 48294
rect 16986 43058 17222 43294
rect 16986 38058 17222 38294
rect 16986 33216 17222 33294
rect 16986 33152 17016 33216
rect 17016 33152 17032 33216
rect 17032 33152 17096 33216
rect 17096 33152 17112 33216
rect 17112 33152 17176 33216
rect 17176 33152 17192 33216
rect 17192 33152 17222 33216
rect 16986 33058 17222 33152
rect 16986 28058 17222 28294
rect 16986 23058 17222 23294
rect 16986 18058 17222 18294
rect 16986 13058 17222 13294
rect 16986 8192 17222 8294
rect 16986 8128 17016 8192
rect 17016 8128 17032 8192
rect 17032 8128 17096 8192
rect 17096 8128 17112 8192
rect 17112 8128 17176 8192
rect 17176 8128 17192 8192
rect 17192 8128 17222 8192
rect 16986 8058 17222 8128
rect 16986 3058 17222 3294
rect 17646 68718 17882 68954
rect 17646 63718 17882 63954
rect 21986 68058 22222 68294
rect 17646 58784 17882 58954
rect 17646 58720 17676 58784
rect 17676 58720 17692 58784
rect 17692 58720 17756 58784
rect 17756 58720 17772 58784
rect 17772 58720 17836 58784
rect 17836 58720 17852 58784
rect 17852 58720 17882 58784
rect 17646 58718 17882 58720
rect 17646 53718 17882 53954
rect 17646 48928 17676 48954
rect 17676 48928 17692 48954
rect 17692 48928 17756 48954
rect 17756 48928 17772 48954
rect 17772 48928 17836 48954
rect 17836 48928 17852 48954
rect 17852 48928 17882 48954
rect 17646 48718 17882 48928
rect 17646 43718 17882 43954
rect 17646 38718 17882 38954
rect 17646 33760 17882 33954
rect 17646 33718 17676 33760
rect 17676 33718 17692 33760
rect 17692 33718 17756 33760
rect 17756 33718 17772 33760
rect 17772 33718 17836 33760
rect 17836 33718 17852 33760
rect 17852 33718 17882 33760
rect 17646 28718 17882 28954
rect 17646 23904 17676 23954
rect 17676 23904 17692 23954
rect 17692 23904 17756 23954
rect 17756 23904 17772 23954
rect 17772 23904 17836 23954
rect 17836 23904 17852 23954
rect 17852 23904 17882 23954
rect 17646 23718 17882 23904
rect 17646 18718 17882 18954
rect 17646 13718 17882 13954
rect 21986 63058 22222 63294
rect 21986 58240 22222 58294
rect 21986 58176 22016 58240
rect 22016 58176 22032 58240
rect 22032 58176 22096 58240
rect 22096 58176 22112 58240
rect 22112 58176 22176 58240
rect 22176 58176 22192 58240
rect 22192 58176 22222 58240
rect 21986 58058 22222 58176
rect 21986 53058 22222 53294
rect 21986 48058 22222 48294
rect 21986 43058 22222 43294
rect 21986 38058 22222 38294
rect 21986 33216 22222 33294
rect 21986 33152 22016 33216
rect 22016 33152 22032 33216
rect 22032 33152 22096 33216
rect 22096 33152 22112 33216
rect 22112 33152 22176 33216
rect 22176 33152 22192 33216
rect 22192 33152 22222 33216
rect 21986 33058 22222 33152
rect 21986 28058 22222 28294
rect 21986 23058 22222 23294
rect 21986 18058 22222 18294
rect 21986 13058 22222 13294
rect 17646 8736 17882 8954
rect 17646 8718 17676 8736
rect 17676 8718 17692 8736
rect 17692 8718 17756 8736
rect 17756 8718 17772 8736
rect 17772 8718 17836 8736
rect 17836 8718 17852 8736
rect 17852 8718 17882 8736
rect 17646 3718 17882 3954
rect 21986 8192 22222 8294
rect 21986 8128 22016 8192
rect 22016 8128 22032 8192
rect 22032 8128 22096 8192
rect 22096 8128 22112 8192
rect 22112 8128 22176 8192
rect 22176 8128 22192 8192
rect 22192 8128 22222 8192
rect 21986 8058 22222 8128
rect 21986 3058 22222 3294
rect 22646 68718 22882 68954
rect 26986 68058 27222 68294
rect 22646 63718 22882 63954
rect 22646 58784 22882 58954
rect 22646 58720 22676 58784
rect 22676 58720 22692 58784
rect 22692 58720 22756 58784
rect 22756 58720 22772 58784
rect 22772 58720 22836 58784
rect 22836 58720 22852 58784
rect 22852 58720 22882 58784
rect 22646 58718 22882 58720
rect 22646 53718 22882 53954
rect 22646 48928 22676 48954
rect 22676 48928 22692 48954
rect 22692 48928 22756 48954
rect 22756 48928 22772 48954
rect 22772 48928 22836 48954
rect 22836 48928 22852 48954
rect 22852 48928 22882 48954
rect 22646 48718 22882 48928
rect 22646 43718 22882 43954
rect 26986 63058 27222 63294
rect 22646 38718 22882 38954
rect 22646 33760 22882 33954
rect 22646 33718 22676 33760
rect 22676 33718 22692 33760
rect 22692 33718 22756 33760
rect 22756 33718 22772 33760
rect 22772 33718 22836 33760
rect 22836 33718 22852 33760
rect 22852 33718 22882 33760
rect 22646 28718 22882 28954
rect 22646 23904 22676 23954
rect 22676 23904 22692 23954
rect 22692 23904 22756 23954
rect 22756 23904 22772 23954
rect 22772 23904 22836 23954
rect 22836 23904 22852 23954
rect 22852 23904 22882 23954
rect 22646 23718 22882 23904
rect 22646 18718 22882 18954
rect 26986 58240 27222 58294
rect 26986 58176 27016 58240
rect 27016 58176 27032 58240
rect 27032 58176 27096 58240
rect 27096 58176 27112 58240
rect 27112 58176 27176 58240
rect 27176 58176 27192 58240
rect 27192 58176 27222 58240
rect 26986 58058 27222 58176
rect 26986 53058 27222 53294
rect 26986 48058 27222 48294
rect 26986 43058 27222 43294
rect 26986 38058 27222 38294
rect 26986 33216 27222 33294
rect 26986 33152 27016 33216
rect 27016 33152 27032 33216
rect 27032 33152 27096 33216
rect 27096 33152 27112 33216
rect 27112 33152 27176 33216
rect 27176 33152 27192 33216
rect 27192 33152 27222 33216
rect 26986 33058 27222 33152
rect 26986 28058 27222 28294
rect 26986 23058 27222 23294
rect 26986 18058 27222 18294
rect 22646 13718 22882 13954
rect 22646 8736 22882 8954
rect 22646 8718 22676 8736
rect 22676 8718 22692 8736
rect 22692 8718 22756 8736
rect 22756 8718 22772 8736
rect 22772 8718 22836 8736
rect 22836 8718 22852 8736
rect 22852 8718 22882 8736
rect 22646 3718 22882 3954
rect 26986 13058 27222 13294
rect 26986 8192 27222 8294
rect 26986 8128 27016 8192
rect 27016 8128 27032 8192
rect 27032 8128 27096 8192
rect 27096 8128 27112 8192
rect 27112 8128 27176 8192
rect 27176 8128 27192 8192
rect 27192 8128 27222 8192
rect 26986 8058 27222 8128
rect 26986 3058 27222 3294
rect 27646 68718 27882 68954
rect 27646 63718 27882 63954
rect 27646 58784 27882 58954
rect 27646 58720 27676 58784
rect 27676 58720 27692 58784
rect 27692 58720 27756 58784
rect 27756 58720 27772 58784
rect 27772 58720 27836 58784
rect 27836 58720 27852 58784
rect 27852 58720 27882 58784
rect 27646 58718 27882 58720
rect 27646 53718 27882 53954
rect 27646 48928 27676 48954
rect 27676 48928 27692 48954
rect 27692 48928 27756 48954
rect 27756 48928 27772 48954
rect 27772 48928 27836 48954
rect 27836 48928 27852 48954
rect 27852 48928 27882 48954
rect 27646 48718 27882 48928
rect 27646 43718 27882 43954
rect 31986 68058 32222 68294
rect 31986 63058 32222 63294
rect 31986 58240 32222 58294
rect 31986 58176 32016 58240
rect 32016 58176 32032 58240
rect 32032 58176 32096 58240
rect 32096 58176 32112 58240
rect 32112 58176 32176 58240
rect 32176 58176 32192 58240
rect 32192 58176 32222 58240
rect 31986 58058 32222 58176
rect 31986 53058 32222 53294
rect 31986 48058 32222 48294
rect 31986 43058 32222 43294
rect 27646 38718 27882 38954
rect 27646 33760 27882 33954
rect 27646 33718 27676 33760
rect 27676 33718 27692 33760
rect 27692 33718 27756 33760
rect 27756 33718 27772 33760
rect 27772 33718 27836 33760
rect 27836 33718 27852 33760
rect 27852 33718 27882 33760
rect 31986 38058 32222 38294
rect 31986 33216 32222 33294
rect 31986 33152 32016 33216
rect 32016 33152 32032 33216
rect 32032 33152 32096 33216
rect 32096 33152 32112 33216
rect 32112 33152 32176 33216
rect 32176 33152 32192 33216
rect 32192 33152 32222 33216
rect 31986 33058 32222 33152
rect 27646 28718 27882 28954
rect 27646 23904 27676 23954
rect 27676 23904 27692 23954
rect 27692 23904 27756 23954
rect 27756 23904 27772 23954
rect 27772 23904 27836 23954
rect 27836 23904 27852 23954
rect 27852 23904 27882 23954
rect 27646 23718 27882 23904
rect 27646 18718 27882 18954
rect 27646 13718 27882 13954
rect 27646 8736 27882 8954
rect 27646 8718 27676 8736
rect 27676 8718 27692 8736
rect 27692 8718 27756 8736
rect 27756 8718 27772 8736
rect 27772 8718 27836 8736
rect 27836 8718 27852 8736
rect 27852 8718 27882 8736
rect 27646 3718 27882 3954
rect 31986 28058 32222 28294
rect 31986 23058 32222 23294
rect 31986 18058 32222 18294
rect 31986 13058 32222 13294
rect 31986 8192 32222 8294
rect 31986 8128 32016 8192
rect 32016 8128 32032 8192
rect 32032 8128 32096 8192
rect 32096 8128 32112 8192
rect 32112 8128 32176 8192
rect 32176 8128 32192 8192
rect 32192 8128 32222 8192
rect 31986 8058 32222 8128
rect 31986 3058 32222 3294
rect 32646 68718 32882 68954
rect 32646 63718 32882 63954
rect 32646 58784 32882 58954
rect 32646 58720 32676 58784
rect 32676 58720 32692 58784
rect 32692 58720 32756 58784
rect 32756 58720 32772 58784
rect 32772 58720 32836 58784
rect 32836 58720 32852 58784
rect 32852 58720 32882 58784
rect 32646 58718 32882 58720
rect 32646 53718 32882 53954
rect 36986 68058 37222 68294
rect 36986 63058 37222 63294
rect 36986 58240 37222 58294
rect 36986 58176 37016 58240
rect 37016 58176 37032 58240
rect 37032 58176 37096 58240
rect 37096 58176 37112 58240
rect 37112 58176 37176 58240
rect 37176 58176 37192 58240
rect 37192 58176 37222 58240
rect 36986 58058 37222 58176
rect 36986 53058 37222 53294
rect 32646 48928 32676 48954
rect 32676 48928 32692 48954
rect 32692 48928 32756 48954
rect 32756 48928 32772 48954
rect 32772 48928 32836 48954
rect 32836 48928 32852 48954
rect 32852 48928 32882 48954
rect 32646 48718 32882 48928
rect 32646 43718 32882 43954
rect 32646 38718 32882 38954
rect 32646 33760 32882 33954
rect 32646 33718 32676 33760
rect 32676 33718 32692 33760
rect 32692 33718 32756 33760
rect 32756 33718 32772 33760
rect 32772 33718 32836 33760
rect 32836 33718 32852 33760
rect 32852 33718 32882 33760
rect 32646 28718 32882 28954
rect 32646 23904 32676 23954
rect 32676 23904 32692 23954
rect 32692 23904 32756 23954
rect 32756 23904 32772 23954
rect 32772 23904 32836 23954
rect 32836 23904 32852 23954
rect 32852 23904 32882 23954
rect 32646 23718 32882 23904
rect 32646 18718 32882 18954
rect 32646 13718 32882 13954
rect 36986 48058 37222 48294
rect 36986 43058 37222 43294
rect 36986 38058 37222 38294
rect 36986 33216 37222 33294
rect 36986 33152 37016 33216
rect 37016 33152 37032 33216
rect 37032 33152 37096 33216
rect 37096 33152 37112 33216
rect 37112 33152 37176 33216
rect 37176 33152 37192 33216
rect 37192 33152 37222 33216
rect 36986 33058 37222 33152
rect 36986 28058 37222 28294
rect 36986 23058 37222 23294
rect 36986 18058 37222 18294
rect 36986 13058 37222 13294
rect 32646 8736 32882 8954
rect 32646 8718 32676 8736
rect 32676 8718 32692 8736
rect 32692 8718 32756 8736
rect 32756 8718 32772 8736
rect 32772 8718 32836 8736
rect 32836 8718 32852 8736
rect 32852 8718 32882 8736
rect 32646 3718 32882 3954
rect 36986 8192 37222 8294
rect 36986 8128 37016 8192
rect 37016 8128 37032 8192
rect 37032 8128 37096 8192
rect 37096 8128 37112 8192
rect 37112 8128 37176 8192
rect 37176 8128 37192 8192
rect 37192 8128 37222 8192
rect 36986 8058 37222 8128
rect 36986 3058 37222 3294
rect 37646 68718 37882 68954
rect 37646 63718 37882 63954
rect 37646 58784 37882 58954
rect 37646 58720 37676 58784
rect 37676 58720 37692 58784
rect 37692 58720 37756 58784
rect 37756 58720 37772 58784
rect 37772 58720 37836 58784
rect 37836 58720 37852 58784
rect 37852 58720 37882 58784
rect 37646 58718 37882 58720
rect 37646 53718 37882 53954
rect 37646 48928 37676 48954
rect 37676 48928 37692 48954
rect 37692 48928 37756 48954
rect 37756 48928 37772 48954
rect 37772 48928 37836 48954
rect 37836 48928 37852 48954
rect 37852 48928 37882 48954
rect 37646 48718 37882 48928
rect 37646 43718 37882 43954
rect 37646 38718 37882 38954
rect 37646 33760 37882 33954
rect 37646 33718 37676 33760
rect 37676 33718 37692 33760
rect 37692 33718 37756 33760
rect 37756 33718 37772 33760
rect 37772 33718 37836 33760
rect 37836 33718 37852 33760
rect 37852 33718 37882 33760
rect 37646 28718 37882 28954
rect 37646 23904 37676 23954
rect 37676 23904 37692 23954
rect 37692 23904 37756 23954
rect 37756 23904 37772 23954
rect 37772 23904 37836 23954
rect 37836 23904 37852 23954
rect 37852 23904 37882 23954
rect 37646 23718 37882 23904
rect 37646 18718 37882 18954
rect 37646 13718 37882 13954
rect 37646 8736 37882 8954
rect 37646 8718 37676 8736
rect 37676 8718 37692 8736
rect 37692 8718 37756 8736
rect 37756 8718 37772 8736
rect 37772 8718 37836 8736
rect 37836 8718 37852 8736
rect 37852 8718 37882 8736
rect 37646 3718 37882 3954
<< metal5 >>
rect 1056 68954 40896 68996
rect 1056 68718 2646 68954
rect 2882 68718 7646 68954
rect 7882 68718 12646 68954
rect 12882 68718 17646 68954
rect 17882 68718 22646 68954
rect 22882 68718 27646 68954
rect 27882 68718 32646 68954
rect 32882 68718 37646 68954
rect 37882 68718 40896 68954
rect 1056 68676 40896 68718
rect 1056 68294 40896 68336
rect 1056 68058 1986 68294
rect 2222 68058 6986 68294
rect 7222 68058 11986 68294
rect 12222 68058 16986 68294
rect 17222 68058 21986 68294
rect 22222 68058 26986 68294
rect 27222 68058 31986 68294
rect 32222 68058 36986 68294
rect 37222 68058 40896 68294
rect 1056 68016 40896 68058
rect 1056 63954 40896 63996
rect 1056 63718 2646 63954
rect 2882 63718 7646 63954
rect 7882 63718 12646 63954
rect 12882 63718 17646 63954
rect 17882 63718 22646 63954
rect 22882 63718 27646 63954
rect 27882 63718 32646 63954
rect 32882 63718 37646 63954
rect 37882 63718 40896 63954
rect 1056 63676 40896 63718
rect 1056 63294 40896 63336
rect 1056 63058 1986 63294
rect 2222 63058 6986 63294
rect 7222 63058 11986 63294
rect 12222 63058 16986 63294
rect 17222 63058 21986 63294
rect 22222 63058 26986 63294
rect 27222 63058 31986 63294
rect 32222 63058 36986 63294
rect 37222 63058 40896 63294
rect 1056 63016 40896 63058
rect 1056 58954 40896 58996
rect 1056 58718 2646 58954
rect 2882 58718 7646 58954
rect 7882 58718 12646 58954
rect 12882 58718 17646 58954
rect 17882 58718 22646 58954
rect 22882 58718 27646 58954
rect 27882 58718 32646 58954
rect 32882 58718 37646 58954
rect 37882 58718 40896 58954
rect 1056 58676 40896 58718
rect 1056 58294 40896 58336
rect 1056 58058 1986 58294
rect 2222 58058 6986 58294
rect 7222 58058 11986 58294
rect 12222 58058 16986 58294
rect 17222 58058 21986 58294
rect 22222 58058 26986 58294
rect 27222 58058 31986 58294
rect 32222 58058 36986 58294
rect 37222 58058 40896 58294
rect 1056 58016 40896 58058
rect 1056 53954 40896 53996
rect 1056 53718 2646 53954
rect 2882 53718 7646 53954
rect 7882 53718 12646 53954
rect 12882 53718 17646 53954
rect 17882 53718 22646 53954
rect 22882 53718 27646 53954
rect 27882 53718 32646 53954
rect 32882 53718 37646 53954
rect 37882 53718 40896 53954
rect 1056 53676 40896 53718
rect 1056 53294 40896 53336
rect 1056 53058 1986 53294
rect 2222 53058 6986 53294
rect 7222 53058 11986 53294
rect 12222 53058 16986 53294
rect 17222 53058 21986 53294
rect 22222 53058 26986 53294
rect 27222 53058 31986 53294
rect 32222 53058 36986 53294
rect 37222 53058 40896 53294
rect 1056 53016 40896 53058
rect 1056 48954 40896 48996
rect 1056 48718 2646 48954
rect 2882 48718 7646 48954
rect 7882 48718 12646 48954
rect 12882 48718 17646 48954
rect 17882 48718 22646 48954
rect 22882 48718 27646 48954
rect 27882 48718 32646 48954
rect 32882 48718 37646 48954
rect 37882 48718 40896 48954
rect 1056 48676 40896 48718
rect 1056 48294 40896 48336
rect 1056 48058 1986 48294
rect 2222 48058 6986 48294
rect 7222 48058 11986 48294
rect 12222 48058 16986 48294
rect 17222 48058 21986 48294
rect 22222 48058 26986 48294
rect 27222 48058 31986 48294
rect 32222 48058 36986 48294
rect 37222 48058 40896 48294
rect 1056 48016 40896 48058
rect 1056 43954 40896 43996
rect 1056 43718 2646 43954
rect 2882 43718 7646 43954
rect 7882 43718 12646 43954
rect 12882 43718 17646 43954
rect 17882 43718 22646 43954
rect 22882 43718 27646 43954
rect 27882 43718 32646 43954
rect 32882 43718 37646 43954
rect 37882 43718 40896 43954
rect 1056 43676 40896 43718
rect 1056 43294 40896 43336
rect 1056 43058 1986 43294
rect 2222 43058 6986 43294
rect 7222 43058 11986 43294
rect 12222 43058 16986 43294
rect 17222 43058 21986 43294
rect 22222 43058 26986 43294
rect 27222 43058 31986 43294
rect 32222 43058 36986 43294
rect 37222 43058 40896 43294
rect 1056 43016 40896 43058
rect 1056 38954 40896 38996
rect 1056 38718 2646 38954
rect 2882 38718 7646 38954
rect 7882 38718 12646 38954
rect 12882 38718 17646 38954
rect 17882 38718 22646 38954
rect 22882 38718 27646 38954
rect 27882 38718 32646 38954
rect 32882 38718 37646 38954
rect 37882 38718 40896 38954
rect 1056 38676 40896 38718
rect 1056 38294 40896 38336
rect 1056 38058 1986 38294
rect 2222 38058 6986 38294
rect 7222 38058 11986 38294
rect 12222 38058 16986 38294
rect 17222 38058 21986 38294
rect 22222 38058 26986 38294
rect 27222 38058 31986 38294
rect 32222 38058 36986 38294
rect 37222 38058 40896 38294
rect 1056 38016 40896 38058
rect 1056 33954 40896 33996
rect 1056 33718 2646 33954
rect 2882 33718 7646 33954
rect 7882 33718 12646 33954
rect 12882 33718 17646 33954
rect 17882 33718 22646 33954
rect 22882 33718 27646 33954
rect 27882 33718 32646 33954
rect 32882 33718 37646 33954
rect 37882 33718 40896 33954
rect 1056 33676 40896 33718
rect 1056 33294 40896 33336
rect 1056 33058 1986 33294
rect 2222 33058 6986 33294
rect 7222 33058 11986 33294
rect 12222 33058 16986 33294
rect 17222 33058 21986 33294
rect 22222 33058 26986 33294
rect 27222 33058 31986 33294
rect 32222 33058 36986 33294
rect 37222 33058 40896 33294
rect 1056 33016 40896 33058
rect 1056 28954 40896 28996
rect 1056 28718 2646 28954
rect 2882 28718 7646 28954
rect 7882 28718 12646 28954
rect 12882 28718 17646 28954
rect 17882 28718 22646 28954
rect 22882 28718 27646 28954
rect 27882 28718 32646 28954
rect 32882 28718 37646 28954
rect 37882 28718 40896 28954
rect 1056 28676 40896 28718
rect 1056 28294 40896 28336
rect 1056 28058 1986 28294
rect 2222 28058 6986 28294
rect 7222 28058 11986 28294
rect 12222 28058 16986 28294
rect 17222 28058 21986 28294
rect 22222 28058 26986 28294
rect 27222 28058 31986 28294
rect 32222 28058 36986 28294
rect 37222 28058 40896 28294
rect 1056 28016 40896 28058
rect 1056 23954 40896 23996
rect 1056 23718 2646 23954
rect 2882 23718 7646 23954
rect 7882 23718 12646 23954
rect 12882 23718 17646 23954
rect 17882 23718 22646 23954
rect 22882 23718 27646 23954
rect 27882 23718 32646 23954
rect 32882 23718 37646 23954
rect 37882 23718 40896 23954
rect 1056 23676 40896 23718
rect 1056 23294 40896 23336
rect 1056 23058 1986 23294
rect 2222 23058 6986 23294
rect 7222 23058 11986 23294
rect 12222 23058 16986 23294
rect 17222 23058 21986 23294
rect 22222 23058 26986 23294
rect 27222 23058 31986 23294
rect 32222 23058 36986 23294
rect 37222 23058 40896 23294
rect 1056 23016 40896 23058
rect 1056 18954 40896 18996
rect 1056 18718 2646 18954
rect 2882 18718 7646 18954
rect 7882 18718 12646 18954
rect 12882 18718 17646 18954
rect 17882 18718 22646 18954
rect 22882 18718 27646 18954
rect 27882 18718 32646 18954
rect 32882 18718 37646 18954
rect 37882 18718 40896 18954
rect 1056 18676 40896 18718
rect 1056 18294 40896 18336
rect 1056 18058 1986 18294
rect 2222 18058 6986 18294
rect 7222 18058 11986 18294
rect 12222 18058 16986 18294
rect 17222 18058 21986 18294
rect 22222 18058 26986 18294
rect 27222 18058 31986 18294
rect 32222 18058 36986 18294
rect 37222 18058 40896 18294
rect 1056 18016 40896 18058
rect 1056 13954 40896 13996
rect 1056 13718 2646 13954
rect 2882 13718 7646 13954
rect 7882 13718 12646 13954
rect 12882 13718 17646 13954
rect 17882 13718 22646 13954
rect 22882 13718 27646 13954
rect 27882 13718 32646 13954
rect 32882 13718 37646 13954
rect 37882 13718 40896 13954
rect 1056 13676 40896 13718
rect 1056 13294 40896 13336
rect 1056 13058 1986 13294
rect 2222 13058 6986 13294
rect 7222 13058 11986 13294
rect 12222 13058 16986 13294
rect 17222 13058 21986 13294
rect 22222 13058 26986 13294
rect 27222 13058 31986 13294
rect 32222 13058 36986 13294
rect 37222 13058 40896 13294
rect 1056 13016 40896 13058
rect 1056 8954 40896 8996
rect 1056 8718 2646 8954
rect 2882 8718 7646 8954
rect 7882 8718 12646 8954
rect 12882 8718 17646 8954
rect 17882 8718 22646 8954
rect 22882 8718 27646 8954
rect 27882 8718 32646 8954
rect 32882 8718 37646 8954
rect 37882 8718 40896 8954
rect 1056 8676 40896 8718
rect 1056 8294 40896 8336
rect 1056 8058 1986 8294
rect 2222 8058 6986 8294
rect 7222 8058 11986 8294
rect 12222 8058 16986 8294
rect 17222 8058 21986 8294
rect 22222 8058 26986 8294
rect 27222 8058 31986 8294
rect 32222 8058 36986 8294
rect 37222 8058 40896 8294
rect 1056 8016 40896 8058
rect 1056 3954 40896 3996
rect 1056 3718 2646 3954
rect 2882 3718 7646 3954
rect 7882 3718 12646 3954
rect 12882 3718 17646 3954
rect 17882 3718 22646 3954
rect 22882 3718 27646 3954
rect 27882 3718 32646 3954
rect 32882 3718 37646 3954
rect 37882 3718 40896 3954
rect 1056 3676 40896 3718
rect 1056 3294 40896 3336
rect 1056 3058 1986 3294
rect 2222 3058 6986 3294
rect 7222 3058 11986 3294
rect 12222 3058 16986 3294
rect 17222 3058 21986 3294
rect 22222 3058 26986 3294
rect 27222 3058 31986 3294
rect 32222 3058 36986 3294
rect 37222 3058 40896 3294
rect 1056 3016 40896 3058
use sky130_fd_sc_hd__buf_8  _248_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 2576 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_4  _249_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4140 0 1 58752
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _250_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6348 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_16  _251_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 5612 0 1 54400
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_12  _252_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 15732 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__or2_1  _253_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 31372 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_4  _254_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3772 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__inv_4  _255_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 11868 0 1 65280
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_8  _256_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 38732 0 -1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__nand3_4  _257_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 33672 0 -1 15232
box -38 -48 1326 592
use sky130_fd_sc_hd__nor2_8  _258_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 33856 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__nor2_4  _259_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 37260 0 -1 48960
box -38 -48 866 592
use sky130_fd_sc_hd__o211a_4  _260_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 1564 0 1 8704
box -38 -48 1326 592
use sky130_fd_sc_hd__a31o_2  _261_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 38088 0 1 67456
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_2  _262_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 14260 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__buf_8  _263_
timestamp 1704896540
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_2  _264_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 15548 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_8  _265_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 32568 0 1 33728
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_12  _266_
timestamp 1704896540
transform 1 0 9016 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_8  _267_
timestamp 1704896540
transform 1 0 7452 0 -1 45696
box -38 -48 1050 592
use sky130_fd_sc_hd__nor2_8  _268_
timestamp 1704896540
transform 1 0 7084 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__or3b_2  _269_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 27968 0 1 63104
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_8  _270_
timestamp 1704896540
transform 1 0 31004 0 -1 47872
box -38 -48 1050 592
use sky130_fd_sc_hd__a21oi_2  _271_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 27232 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _272_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 17388 0 -1 48960
box -38 -48 682 592
use sky130_fd_sc_hd__and3_4  _273_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 13524 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__or2b_2  _274_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 18584 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__nand3b_4  _275_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 33948 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__a21oi_2  _276_
timestamp 1704896540
transform 1 0 10212 0 -1 48960
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _277_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 17112 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_2  _278_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 10212 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__or3_4  _279_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 16284 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__or2b_1  _280_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 19872 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _281_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 8556 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and4_2  _282_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 37996 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _283_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 39008 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__and3b_1  _284_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 19228 0 1 59840
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_2  _285_
timestamp 1704896540
transform -1 0 23092 0 1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_2  _286_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 2852 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_2  _287_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 18584 0 -1 63104
box -38 -48 866 592
use sky130_fd_sc_hd__buf_8  _288_
timestamp 1704896540
transform 1 0 12696 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_12  _289_
timestamp 1704896540
transform -1 0 37720 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__nand2_2  _290_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 6808 0 -1 45696
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _291_
timestamp 1704896540
transform -1 0 18860 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _292_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6992 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_2  _293_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 12696 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_4  _294_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5888 0 1 44608
box -38 -48 2062 592
use sky130_fd_sc_hd__and2_4  _295_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 32200 0 1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_2  _296_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 32292 0 1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _297_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 9936 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_4  _298_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 37536 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__xnor2_4  _299_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 23000 0 -1 36992
box -38 -48 2062 592
use sky130_fd_sc_hd__xor2_4  _300_
timestamp 1704896540
transform -1 0 28060 0 1 8704
box -38 -48 2062 592
use sky130_fd_sc_hd__a21o_4  _301_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 38456 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_2  _302_
timestamp 1704896540
transform -1 0 37812 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_2  _303_
timestamp 1704896540
transform 1 0 12972 0 1 67456
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_8  _304_
timestamp 1704896540
transform 1 0 17480 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__and2b_2  _305_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 37444 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _306_
timestamp 1704896540
transform -1 0 20700 0 1 64192
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_2  _307_
timestamp 1704896540
transform -1 0 25024 0 1 48960
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _308_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 1840 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_2  _309_
timestamp 1704896540
transform -1 0 16652 0 1 55488
box -38 -48 866 592
use sky130_fd_sc_hd__buf_12  _310_
timestamp 1704896540
transform 1 0 38272 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__and2_1  _311_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 31556 0 1 68544
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_4  _312_
timestamp 1704896540
transform 1 0 7360 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  _313_
timestamp 1704896540
transform 1 0 35696 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__a211oi_4  _314_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 38732 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__o311a_4  _315_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 13524 0 1 68544
box -38 -48 1602 592
use sky130_fd_sc_hd__o21ai_4  _316_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 16192 0 -1 53312
box -38 -48 1234 592
use sky130_fd_sc_hd__or3_4  _317_
timestamp 1704896540
transform 1 0 16652 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__and3_2  _318_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 4324 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _319_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 39192 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_2  _320_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 27140 0 1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  _321_
timestamp 1704896540
transform 1 0 16284 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  _322_
timestamp 1704896540
transform -1 0 8280 0 1 66368
box -38 -48 866 592
use sky130_fd_sc_hd__and4_4  _323_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 19228 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__a22oi_4  _324_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 39008 0 -1 57664
box -38 -48 1602 592
use sky130_fd_sc_hd__or3_4  _325_
timestamp 1704896540
transform 1 0 24380 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_4  _326_
timestamp 1704896540
transform -1 0 11408 0 -1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__and4_4  _327_
timestamp 1704896540
transform -1 0 28980 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_4  _328_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 20332 0 1 42432
box -38 -48 1326 592
use sky130_fd_sc_hd__and3_1  _329_
timestamp 1704896540
transform 1 0 32108 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_4  _330_
timestamp 1704896540
transform 1 0 7544 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__and2b_2  _331_
timestamp 1704896540
transform 1 0 38824 0 1 52224
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_4  _332_
timestamp 1704896540
transform -1 0 32844 0 1 51136
box -38 -48 2062 592
use sky130_fd_sc_hd__nand2_4  _333_
timestamp 1704896540
transform 1 0 3864 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _334_
timestamp 1704896540
transform 1 0 8096 0 -1 63104
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _335_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 3588 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _336_
timestamp 1704896540
transform -1 0 6992 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a311o_1  _337_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 10488 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _338_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 9384 0 -1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _339_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 2668 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  _340_
timestamp 1704896540
transform 1 0 2208 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__a31o_4  _341_
timestamp 1704896540
transform -1 0 30636 0 -1 35904
box -38 -48 1326 592
use sky130_fd_sc_hd__buf_8  _342_
timestamp 1704896540
transform 1 0 26956 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_2  _343_
timestamp 1704896540
transform 1 0 8188 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__and4_2  _344_
timestamp 1704896540
transform 1 0 6532 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__clkinv_4  _345_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 33764 0 1 54400
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _346_
timestamp 1704896540
transform 1 0 13156 0 -1 62016
box -38 -48 682 592
use sky130_fd_sc_hd__and4_4  _347_
timestamp 1704896540
transform 1 0 11500 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__a22oi_4  _348_
timestamp 1704896540
transform 1 0 6624 0 -1 26112
box -38 -48 1602 592
use sky130_fd_sc_hd__or3_4  _349_
timestamp 1704896540
transform -1 0 2576 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_4  _350_
timestamp 1704896540
transform -1 0 32016 0 -1 28288
box -38 -48 1234 592
use sky130_fd_sc_hd__o21bai_4  _351_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 22264 0 1 40256
box -38 -48 1418 592
use sky130_fd_sc_hd__and3_4  _352_
timestamp 1704896540
transform 1 0 22908 0 1 58752
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_4  _353_
timestamp 1704896540
transform -1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__or2b_4  _354_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 31832 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_4  _355_
timestamp 1704896540
transform 1 0 3864 0 -1 55488
box -38 -48 2062 592
use sky130_fd_sc_hd__nand2_8  _356_
timestamp 1704896540
transform 1 0 6348 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__or2_4  _357_
timestamp 1704896540
transform 1 0 24656 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _358_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 17848 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__nand3b_4  _359_
timestamp 1704896540
transform 1 0 35696 0 -1 50048
box -38 -48 1510 592
use sky130_fd_sc_hd__and3_2  _360_
timestamp 1704896540
transform 1 0 16652 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_4  _361_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 14536 0 -1 15232
box -38 -48 1326 592
use sky130_fd_sc_hd__xnor2_4  _362_
timestamp 1704896540
transform -1 0 29164 0 1 7616
box -38 -48 2062 592
use sky130_fd_sc_hd__and2_2  _363_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 12420 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _364_
timestamp 1704896540
transform -1 0 27416 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _365_
timestamp 1704896540
transform 1 0 13616 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_2  _366_
timestamp 1704896540
transform 1 0 31556 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_2  _367_
timestamp 1704896540
transform 1 0 19780 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _368_
timestamp 1704896540
transform 1 0 16836 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_4  _369_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 29900 0 1 58752
box -38 -48 1234 592
use sky130_fd_sc_hd__o22a_2  _370_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 7360 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__a311o_1  _371_
timestamp 1704896540
transform -1 0 22356 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _372_
timestamp 1704896540
transform 1 0 38640 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_2  _373_
timestamp 1704896540
transform 1 0 36156 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__buf_12  _374_
timestamp 1704896540
transform 1 0 32108 0 -1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__a21o_4  _375_
timestamp 1704896540
transform -1 0 16560 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__a21o_4  _376_
timestamp 1704896540
transform -1 0 5060 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__xnor2_4  _377_
timestamp 1704896540
transform -1 0 26864 0 -1 33728
box -38 -48 2062 592
use sky130_fd_sc_hd__and2_4  _378_
timestamp 1704896540
transform -1 0 7176 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _379_
timestamp 1704896540
transform 1 0 7360 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _380_
timestamp 1704896540
transform 1 0 3772 0 1 53312
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _381_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 35604 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_4  _382_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 21344 0 -1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__a22o_4  _383_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 9200 0 -1 60928
box -38 -48 1326 592
use sky130_fd_sc_hd__and2_4  _384_
timestamp 1704896540
transform -1 0 17296 0 -1 57664
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_4  _385_
timestamp 1704896540
transform 1 0 6440 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__nand3_4  _386_
timestamp 1704896540
transform 1 0 34684 0 1 27200
box -38 -48 1326 592
use sky130_fd_sc_hd__o21bai_4  _387_
timestamp 1704896540
transform -1 0 3588 0 1 40256
box -38 -48 1418 592
use sky130_fd_sc_hd__nand3_4  _388_
timestamp 1704896540
transform -1 0 35972 0 1 6528
box -38 -48 1326 592
use sky130_fd_sc_hd__a21o_4  _389_
timestamp 1704896540
transform -1 0 38916 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_4  _390_
timestamp 1704896540
transform -1 0 38824 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__and4_4  _391_
timestamp 1704896540
transform 1 0 15088 0 1 53312
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_2  _392_
timestamp 1704896540
transform 1 0 6624 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_2  _393_
timestamp 1704896540
transform 1 0 29624 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_4  _394_
timestamp 1704896540
transform -1 0 18676 0 -1 22848
box -38 -48 2062 592
use sky130_fd_sc_hd__a21o_4  _395_
timestamp 1704896540
transform 1 0 37260 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__nand3_4  _396_
timestamp 1704896540
transform -1 0 15364 0 1 4352
box -38 -48 1326 592
use sky130_fd_sc_hd__a21o_4  _397_
timestamp 1704896540
transform -1 0 39744 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__and3_4  _398_
timestamp 1704896540
transform 1 0 20148 0 1 62016
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_4  _399_
timestamp 1704896540
transform -1 0 10856 0 -1 67456
box -38 -48 1234 592
use sky130_fd_sc_hd__o21ai_4  _400_
timestamp 1704896540
transform 1 0 6900 0 1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__or3_4  _401_
timestamp 1704896540
transform 1 0 38456 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  _402_
timestamp 1704896540
transform -1 0 32016 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_4  _403_
timestamp 1704896540
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__nand3_2  _404_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 9016 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_2  _405_
timestamp 1704896540
transform -1 0 26220 0 1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _406_
timestamp 1704896540
transform 1 0 3864 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a311o_2  _407_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 22632 0 -1 51136
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _408_
timestamp 1704896540
transform 1 0 39008 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _409_
timestamp 1704896540
transform 1 0 33120 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_2  _410_
timestamp 1704896540
transform 1 0 24104 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_4  _411_
timestamp 1704896540
transform 1 0 28244 0 -1 54400
box -38 -48 1326 592
use sky130_fd_sc_hd__a31o_2  _412_
timestamp 1704896540
transform -1 0 26680 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__and3_4  _413_
timestamp 1704896540
transform -1 0 18768 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_4  _414_
timestamp 1704896540
transform 1 0 31648 0 1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_4  _415_
timestamp 1704896540
transform 1 0 13708 0 -1 50048
box -38 -48 866 592
use sky130_fd_sc_hd__nand4_4  _416_
timestamp 1704896540
transform 1 0 13616 0 -1 33728
box -38 -48 1602 592
use sky130_fd_sc_hd__a22o_4  _417_
timestamp 1704896540
transform -1 0 34960 0 -1 23936
box -38 -48 1326 592
use sky130_fd_sc_hd__and2_4  _418_
timestamp 1704896540
transform -1 0 25116 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_2  _419_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 36616 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_2  _420_
timestamp 1704896540
transform -1 0 5244 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_4  _421_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 30268 0 -1 30464
box -38 -48 1234 592
use sky130_fd_sc_hd__nand3_4  _422_
timestamp 1704896540
transform -1 0 5520 0 -1 52224
box -38 -48 1326 592
use sky130_fd_sc_hd__a21o_4  _423_
timestamp 1704896540
transform -1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_4  _424_
timestamp 1704896540
transform 1 0 26036 0 1 56576
box -38 -48 866 592
use sky130_fd_sc_hd__and3_4  _425_
timestamp 1704896540
transform -1 0 38640 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_2  _426_
timestamp 1704896540
transform -1 0 21620 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_4  _427_
timestamp 1704896540
transform -1 0 2576 0 1 60928
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_4  _428_
timestamp 1704896540
transform 1 0 32568 0 1 19584
box -38 -48 2062 592
use sky130_fd_sc_hd__a21o_4  _429_
timestamp 1704896540
transform 1 0 2208 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__nand3_4  _430_
timestamp 1704896540
transform 1 0 17756 0 1 23936
box -38 -48 1326 592
use sky130_fd_sc_hd__a21bo_4  _431_
timestamp 1704896540
transform 1 0 35144 0 1 67456
box -38 -48 1234 592
use sky130_fd_sc_hd__nand3_4  _432_
timestamp 1704896540
transform -1 0 7912 0 -1 19584
box -38 -48 1326 592
use sky130_fd_sc_hd__a21o_4  _433_
timestamp 1704896540
transform 1 0 30084 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__and3_4  _434_
timestamp 1704896540
transform 1 0 8924 0 1 60928
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_4  _435_
timestamp 1704896540
transform -1 0 11224 0 1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__a211oi_4  _436_
timestamp 1704896540
transform -1 0 21712 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__o211a_2  _437_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 28612 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__a2111oi_4  _438_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 32568 0 1 59840
box -38 -48 2062 592
use sky130_fd_sc_hd__or2_4  _439_
timestamp 1704896540
transform -1 0 31004 0 -1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_2  _440_
timestamp 1704896540
transform 1 0 2208 0 1 65280
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _441_
timestamp 1704896540
transform -1 0 2024 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_4  _442_
timestamp 1704896540
transform 1 0 21252 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_4  _443_
timestamp 1704896540
transform 1 0 14812 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_4  _444_
timestamp 1704896540
transform 1 0 28980 0 -1 60928
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_4  _445_
timestamp 1704896540
transform -1 0 24012 0 -1 33728
box -38 -48 2062 592
use sky130_fd_sc_hd__xor2_4  _446_
timestamp 1704896540
transform 1 0 22908 0 -1 68544
box -38 -48 2062 592
use sky130_fd_sc_hd__nand2_1  _447_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 23460 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _448_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 35236 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _449_
timestamp 1704896540
transform -1 0 33764 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _450_
timestamp 1704896540
transform 1 0 38088 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a311o_2  _451_
timestamp 1704896540
transform 1 0 22908 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_4  _452_
timestamp 1704896540
transform 1 0 24748 0 -1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__a22oi_4  _453_
timestamp 1704896540
transform 1 0 10028 0 1 56576
box -38 -48 1602 592
use sky130_fd_sc_hd__and2_2  _454_
timestamp 1704896540
transform -1 0 19872 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _455_
timestamp 1704896540
transform 1 0 34684 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_4  _456_
timestamp 1704896540
transform -1 0 19044 0 -1 67456
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_2  _457_
timestamp 1704896540
transform -1 0 34040 0 1 64192
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _458_
timestamp 1704896540
transform -1 0 37076 0 -1 53312
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _459_
timestamp 1704896540
transform 1 0 10764 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_2  _460_
timestamp 1704896540
transform -1 0 18124 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_2  _461_
timestamp 1704896540
transform -1 0 19044 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _462_
timestamp 1704896540
transform 1 0 17664 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_2  _463_
timestamp 1704896540
transform 1 0 12696 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__o311a_2  _464_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 26956 0 1 66368
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_4  _465_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 30360 0 -1 39168
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_4  _466_
timestamp 1704896540
transform -1 0 23092 0 1 20672
box -38 -48 1326 592
use sky130_fd_sc_hd__nand4_4  _467_
timestamp 1704896540
transform 1 0 35420 0 -1 66368
box -38 -48 1602 592
use sky130_fd_sc_hd__a22oi_4  _468_
timestamp 1704896540
transform 1 0 28520 0 -1 41344
box -38 -48 1602 592
use sky130_fd_sc_hd__and4_2  _469_
timestamp 1704896540
transform -1 0 4508 0 1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_4  _470_
timestamp 1704896540
transform 1 0 22908 0 -1 42432
box -38 -48 1326 592
use sky130_fd_sc_hd__o211ai_4  _471_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 23552 0 -1 50048
box -38 -48 1602 592
use sky130_fd_sc_hd__a22o_4  _472_
timestamp 1704896540
transform 1 0 25760 0 1 18496
box -38 -48 1326 592
use sky130_fd_sc_hd__nand4_4  _473_
timestamp 1704896540
transform 1 0 11868 0 1 62016
box -38 -48 1602 592
use sky130_fd_sc_hd__a21bo_2  _474_
timestamp 1704896540
transform -1 0 10212 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_2  _475_
timestamp 1704896540
transform -1 0 38548 0 1 58752
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_4  _476_
timestamp 1704896540
transform -1 0 39284 0 -1 67456
box -38 -48 2062 592
use sky130_fd_sc_hd__a21o_4  _477_
timestamp 1704896540
transform -1 0 15824 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__nand3_4  _478_
timestamp 1704896540
transform 1 0 20700 0 1 64192
box -38 -48 1326 592
use sky130_fd_sc_hd__and4_4  _479_
timestamp 1704896540
transform -1 0 4600 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_2  _480_
timestamp 1704896540
transform -1 0 35328 0 1 52224
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_4  _481_
timestamp 1704896540
transform 1 0 18584 0 -1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_2  _482_
timestamp 1704896540
transform 1 0 37812 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_4  _483_
timestamp 1704896540
transform 1 0 37996 0 -1 58752
box -38 -48 2062 592
use sky130_fd_sc_hd__xnor2_2  _484_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 11316 0 -1 51136
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_4  _485_
timestamp 1704896540
transform 1 0 5428 0 1 52224
box -38 -48 2062 592
use sky130_fd_sc_hd__a21o_4  _486_
timestamp 1704896540
transform -1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__nand3_4  _487_
timestamp 1704896540
transform -1 0 21160 0 1 57664
box -38 -48 1326 592
use sky130_fd_sc_hd__nand2_4  _488_
timestamp 1704896540
transform -1 0 32936 0 1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_2  _489_
timestamp 1704896540
transform -1 0 31648 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_4  _490_
timestamp 1704896540
transform -1 0 14812 0 -1 58752
box -38 -48 1326 592
use sky130_fd_sc_hd__a21boi_4  _491_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 3312 0 1 50048
box -38 -48 1418 592
use sky130_fd_sc_hd__a21oi_4  _492_
timestamp 1704896540
transform 1 0 29440 0 -1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__and3_4  _493_
timestamp 1704896540
transform -1 0 26036 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__or3_4  _494_
timestamp 1704896540
transform -1 0 6256 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_4  _495_
timestamp 1704896540
transform -1 0 35880 0 1 62016
box -38 -48 1234 592
use sky130_fd_sc_hd__and3_1  _496_
timestamp 1704896540
transform 1 0 12236 0 -1 51136
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_4  _497_
timestamp 1704896540
transform 1 0 29532 0 1 66368
box -38 -48 1234 592
use sky130_fd_sc_hd__o21a_1  _498_
timestamp 1704896540
transform 1 0 16744 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_4  _499_
timestamp 1704896540
transform 1 0 12788 0 1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__o221a_1  _500_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 24380 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _501_
timestamp 1704896540
transform -1 0 22632 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _502_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 14352 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o32a_4  _503_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 13984 0 1 34816
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 32936 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1704896540
transform 1 0 20516 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1704896540
transform 1 0 38640 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1704896540
transform 1 0 35604 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1704896540
transform -1 0 36984 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1704896540
transform -1 0 35696 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1704896540
transform -1 0 2024 0 1 65280
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1704896540
transform 1 0 17572 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1704896540
transform -1 0 3312 0 1 65280
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1704896540
transform -1 0 37260 0 1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1704896540
transform -1 0 39192 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp 1704896540
transform 1 0 39008 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp 1704896540
transform -1 0 19412 0 -1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp 1704896540
transform -1 0 19412 0 -1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp 1704896540
transform 1 0 38272 0 -1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp 1704896540
transform 1 0 30820 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp 1704896540
transform 1 0 32476 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp 1704896540
transform -1 0 26956 0 1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_19
timestamp 1704896540
transform 1 0 4692 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_20
timestamp 1704896540
transform 1 0 7544 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_21
timestamp 1704896540
transform 1 0 14444 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_22
timestamp 1704896540
transform 1 0 26588 0 1 63104
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_23
timestamp 1704896540
transform 1 0 39008 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_24
timestamp 1704896540
transform -1 0 17940 0 1 62016
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_25
timestamp 1704896540
transform -1 0 34316 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_26
timestamp 1704896540
transform 1 0 28612 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_27
timestamp 1704896540
transform 1 0 23276 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_28
timestamp 1704896540
transform -1 0 18216 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_29
timestamp 1704896540
transform -1 0 12236 0 1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_30
timestamp 1704896540
transform -1 0 5244 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_31
timestamp 1704896540
transform 1 0 31188 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_32
timestamp 1704896540
transform 1 0 26956 0 1 63104
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_33
timestamp 1704896540
transform -1 0 17940 0 1 63104
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_34
timestamp 1704896540
transform -1 0 34316 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_35
timestamp 1704896540
transform -1 0 17940 0 -1 62016
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_36
timestamp 1704896540
transform -1 0 34316 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clone15
timestamp 1704896540
transform 1 0 18308 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clone16
timestamp 1704896540
transform 1 0 23184 0 -1 45696
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clone17
timestamp 1704896540
transform 1 0 12788 0 -1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_12  clone31
timestamp 1704896540
transform 1 0 21804 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 1380 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_21
timestamp 1704896540
transform 1 0 3036 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 1704896540
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1704896540
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_78
timestamp 1704896540
transform 1 0 8280 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 1704896540
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_97
timestamp 1704896540
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109
timestamp 1704896540
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp 1704896540
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_125
timestamp 1704896540
transform 1 0 12604 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_135 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 13524 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_139
timestamp 1704896540
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 1704896540
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_153
timestamp 1704896540
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_165
timestamp 1704896540
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_169
timestamp 1704896540
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_181
timestamp 1704896540
transform 1 0 17756 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_186 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 18216 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_192
timestamp 1704896540
transform 1 0 18768 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_197
timestamp 1704896540
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_209
timestamp 1704896540
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_221
timestamp 1704896540
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_225
timestamp 1704896540
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_237
timestamp 1704896540
transform 1 0 22908 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_243
timestamp 1704896540
transform 1 0 23460 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_249
timestamp 1704896540
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_253
timestamp 1704896540
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_265
timestamp 1704896540
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_277
timestamp 1704896540
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_281
timestamp 1704896540
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_293
timestamp 1704896540
transform 1 0 28060 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_301
timestamp 1704896540
transform 1 0 28796 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_307
timestamp 1704896540
transform 1 0 29348 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_309
timestamp 1704896540
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_321
timestamp 1704896540
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_333
timestamp 1704896540
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_337
timestamp 1704896540
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_349 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 33212 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_357
timestamp 1704896540
transform 1 0 33948 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_363
timestamp 1704896540
transform 1 0 34500 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_365
timestamp 1704896540
transform 1 0 34684 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_377
timestamp 1704896540
transform 1 0 35788 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_389
timestamp 1704896540
transform 1 0 36892 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_393
timestamp 1704896540
transform 1 0 37260 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_405
timestamp 1704896540
transform 1 0 38364 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_411
timestamp 1704896540
transform 1 0 38916 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_414
timestamp 1704896540
transform 1 0 39192 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_421
timestamp 1704896540
transform 1 0 39836 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1704896540
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1704896540
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1704896540
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1704896540
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 1704896540
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1704896540
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1704896540
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1704896540
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 1704896540
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 1704896540
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105
timestamp 1704896540
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1704896540
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1704896540
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 1704896540
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_137
timestamp 1704896540
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_149
timestamp 1704896540
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_161
timestamp 1704896540
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 1704896540
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_169
timestamp 1704896540
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_181
timestamp 1704896540
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_193
timestamp 1704896540
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_205
timestamp 1704896540
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_217
timestamp 1704896540
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_223
timestamp 1704896540
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_225
timestamp 1704896540
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_237
timestamp 1704896540
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_249
timestamp 1704896540
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_261
timestamp 1704896540
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_273
timestamp 1704896540
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_279
timestamp 1704896540
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_281
timestamp 1704896540
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_293
timestamp 1704896540
transform 1 0 28060 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_303
timestamp 1704896540
transform 1 0 28980 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_309
timestamp 1704896540
transform 1 0 29532 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_317
timestamp 1704896540
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_329
timestamp 1704896540
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_335
timestamp 1704896540
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_337
timestamp 1704896540
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_349
timestamp 1704896540
transform 1 0 33212 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_357
timestamp 1704896540
transform 1 0 33948 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_361
timestamp 1704896540
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_373
timestamp 1704896540
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_385
timestamp 1704896540
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_391
timestamp 1704896540
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_393
timestamp 1704896540
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_405
timestamp 1704896540
transform 1 0 38364 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_417
timestamp 1704896540
transform 1 0 39468 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1704896540
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1704896540
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1704896540
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1704896540
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1704896540
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1704896540
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_81
timestamp 1704896540
transform 1 0 8556 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1704896540
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_110
timestamp 1704896540
transform 1 0 11224 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_122
timestamp 1704896540
transform 1 0 12328 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_126
timestamp 1704896540
transform 1 0 12696 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 1704896540
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_153
timestamp 1704896540
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_165
timestamp 1704896540
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_177
timestamp 1704896540
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_189
timestamp 1704896540
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 1704896540
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_197
timestamp 1704896540
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_209
timestamp 1704896540
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_221
timestamp 1704896540
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_233
timestamp 1704896540
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_245
timestamp 1704896540
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_251
timestamp 1704896540
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_253
timestamp 1704896540
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_265
timestamp 1704896540
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_277
timestamp 1704896540
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_289
timestamp 1704896540
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_301
timestamp 1704896540
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_307
timestamp 1704896540
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_309
timestamp 1704896540
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_321
timestamp 1704896540
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_333
timestamp 1704896540
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_345
timestamp 1704896540
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_357
timestamp 1704896540
transform 1 0 33948 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_361
timestamp 1704896540
transform 1 0 34316 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_365
timestamp 1704896540
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_377
timestamp 1704896540
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_389
timestamp 1704896540
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_401
timestamp 1704896540
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_413
timestamp 1704896540
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_419
timestamp 1704896540
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_421
timestamp 1704896540
transform 1 0 39836 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1704896540
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1704896540
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1704896540
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1704896540
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1704896540
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1704896540
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_73
timestamp 1704896540
transform 1 0 7820 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_85
timestamp 1704896540
transform 1 0 8924 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_97
timestamp 1704896540
transform 1 0 10028 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_109
timestamp 1704896540
transform 1 0 11132 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1704896540
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1704896540
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 1704896540
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp 1704896540
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_161
timestamp 1704896540
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1704896540
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 1704896540
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_181
timestamp 1704896540
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_193
timestamp 1704896540
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_205
timestamp 1704896540
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_217
timestamp 1704896540
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_223
timestamp 1704896540
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_225
timestamp 1704896540
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_237
timestamp 1704896540
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_249
timestamp 1704896540
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_261
timestamp 1704896540
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_273
timestamp 1704896540
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_279
timestamp 1704896540
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_281
timestamp 1704896540
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_293
timestamp 1704896540
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_305
timestamp 1704896540
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_317
timestamp 1704896540
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_329
timestamp 1704896540
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_335
timestamp 1704896540
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_337
timestamp 1704896540
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_349
timestamp 1704896540
transform 1 0 33212 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_357
timestamp 1704896540
transform 1 0 33948 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_361
timestamp 1704896540
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_373
timestamp 1704896540
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_385
timestamp 1704896540
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_391
timestamp 1704896540
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_393
timestamp 1704896540
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_405
timestamp 1704896540
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_417
timestamp 1704896540
transform 1 0 39468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1704896540
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1704896540
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_38
timestamp 1704896540
transform 1 0 4600 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_50
timestamp 1704896540
transform 1 0 5704 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_58
timestamp 1704896540
transform 1 0 6440 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_68
timestamp 1704896540
transform 1 0 7360 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_80
timestamp 1704896540
transform 1 0 8464 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1704896540
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1704896540
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 1704896540
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 1704896540
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 1704896540
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 1704896540
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_155
timestamp 1704896540
transform 1 0 15364 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_167
timestamp 1704896540
transform 1 0 16468 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_179
timestamp 1704896540
transform 1 0 17572 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_191
timestamp 1704896540
transform 1 0 18676 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 1704896540
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_206
timestamp 1704896540
transform 1 0 20056 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_218
timestamp 1704896540
transform 1 0 21160 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_230
timestamp 1704896540
transform 1 0 22264 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_242
timestamp 1704896540
transform 1 0 23368 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_250
timestamp 1704896540
transform 1 0 24104 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_253
timestamp 1704896540
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_265
timestamp 1704896540
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_277
timestamp 1704896540
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_289
timestamp 1704896540
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_301
timestamp 1704896540
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_307
timestamp 1704896540
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_309
timestamp 1704896540
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_321
timestamp 1704896540
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_333
timestamp 1704896540
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_345
timestamp 1704896540
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_357
timestamp 1704896540
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_363
timestamp 1704896540
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_365
timestamp 1704896540
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_377
timestamp 1704896540
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_389
timestamp 1704896540
transform 1 0 36892 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_393
timestamp 1704896540
transform 1 0 37260 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_411
timestamp 1704896540
transform 1 0 38916 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_419
timestamp 1704896540
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_421
timestamp 1704896540
transform 1 0 39836 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1704896540
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1704896540
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1704896540
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1704896540
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1704896540
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1704896540
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1704896540
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_69
timestamp 1704896540
transform 1 0 7452 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_85
timestamp 1704896540
transform 1 0 8924 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_97
timestamp 1704896540
transform 1 0 10028 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_109
timestamp 1704896540
transform 1 0 11132 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1704896540
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 1704896540
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_137
timestamp 1704896540
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_149
timestamp 1704896540
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_161
timestamp 1704896540
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 1704896540
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 1704896540
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_181
timestamp 1704896540
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_193
timestamp 1704896540
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_205
timestamp 1704896540
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_217
timestamp 1704896540
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 1704896540
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_225
timestamp 1704896540
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_237
timestamp 1704896540
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_249
timestamp 1704896540
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_261
timestamp 1704896540
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_273
timestamp 1704896540
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_279
timestamp 1704896540
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_281
timestamp 1704896540
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_293
timestamp 1704896540
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_305
timestamp 1704896540
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_317
timestamp 1704896540
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_329
timestamp 1704896540
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_335
timestamp 1704896540
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_337
timestamp 1704896540
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_349
timestamp 1704896540
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_361
timestamp 1704896540
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_373
timestamp 1704896540
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_385
timestamp 1704896540
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_391
timestamp 1704896540
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_393
timestamp 1704896540
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_405
timestamp 1704896540
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_417
timestamp 1704896540
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1704896540
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1704896540
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1704896540
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1704896540
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1704896540
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1704896540
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1704896540
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 1704896540
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1704896540
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1704896540
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 1704896540
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_109
timestamp 1704896540
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_121
timestamp 1704896540
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_133
timestamp 1704896540
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1704896540
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 1704896540
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_153
timestamp 1704896540
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_165
timestamp 1704896540
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_177
timestamp 1704896540
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_189
timestamp 1704896540
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp 1704896540
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_197
timestamp 1704896540
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_209
timestamp 1704896540
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_221
timestamp 1704896540
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_233
timestamp 1704896540
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_245
timestamp 1704896540
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_251
timestamp 1704896540
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_253
timestamp 1704896540
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_265
timestamp 1704896540
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_277
timestamp 1704896540
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_289
timestamp 1704896540
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_301
timestamp 1704896540
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_307
timestamp 1704896540
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_309
timestamp 1704896540
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_321
timestamp 1704896540
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_333
timestamp 1704896540
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_345
timestamp 1704896540
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_357
timestamp 1704896540
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_363
timestamp 1704896540
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_365
timestamp 1704896540
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_377
timestamp 1704896540
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_389
timestamp 1704896540
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_401
timestamp 1704896540
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_413
timestamp 1704896540
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_419
timestamp 1704896540
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_421
timestamp 1704896540
transform 1 0 39836 0 1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1704896540
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1704896540
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1704896540
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_39
timestamp 1704896540
transform 1 0 4692 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_45
timestamp 1704896540
transform 1 0 5244 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1704896540
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 1704896540
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_81
timestamp 1704896540
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_93
timestamp 1704896540
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_105
timestamp 1704896540
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1704896540
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 1704896540
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_125
timestamp 1704896540
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_137
timestamp 1704896540
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_149
timestamp 1704896540
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_161
timestamp 1704896540
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 1704896540
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_178
timestamp 1704896540
transform 1 0 17480 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_190
timestamp 1704896540
transform 1 0 18584 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_202
timestamp 1704896540
transform 1 0 19688 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_214
timestamp 1704896540
transform 1 0 20792 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_222
timestamp 1704896540
transform 1 0 21528 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_225
timestamp 1704896540
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_237
timestamp 1704896540
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_249
timestamp 1704896540
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_261
timestamp 1704896540
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_273
timestamp 1704896540
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_279
timestamp 1704896540
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_281
timestamp 1704896540
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_293
timestamp 1704896540
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_305
timestamp 1704896540
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_317
timestamp 1704896540
transform 1 0 30268 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_325
timestamp 1704896540
transform 1 0 31004 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_337
timestamp 1704896540
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_349
timestamp 1704896540
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_361
timestamp 1704896540
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_373
timestamp 1704896540
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_385
timestamp 1704896540
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_391
timestamp 1704896540
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_393
timestamp 1704896540
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_405
timestamp 1704896540
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_417
timestamp 1704896540
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1704896540
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1704896540
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1704896540
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1704896540
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1704896540
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 1704896540
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp 1704896540
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_77
timestamp 1704896540
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1704896540
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 1704896540
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 1704896540
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_109
timestamp 1704896540
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_121
timestamp 1704896540
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_133
timestamp 1704896540
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 1704896540
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 1704896540
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_153
timestamp 1704896540
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_165
timestamp 1704896540
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_177
timestamp 1704896540
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_189
timestamp 1704896540
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_195
timestamp 1704896540
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_197
timestamp 1704896540
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_209
timestamp 1704896540
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_221
timestamp 1704896540
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_233
timestamp 1704896540
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_245
timestamp 1704896540
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_251
timestamp 1704896540
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_253
timestamp 1704896540
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_265
timestamp 1704896540
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_277
timestamp 1704896540
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_289
timestamp 1704896540
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_301
timestamp 1704896540
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_307
timestamp 1704896540
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_309
timestamp 1704896540
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_321
timestamp 1704896540
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_333
timestamp 1704896540
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_345
timestamp 1704896540
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_357
timestamp 1704896540
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_363
timestamp 1704896540
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_379
timestamp 1704896540
transform 1 0 35972 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_391
timestamp 1704896540
transform 1 0 37076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_403
timestamp 1704896540
transform 1 0 38180 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_415
timestamp 1704896540
transform 1 0 39284 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_419
timestamp 1704896540
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_421
timestamp 1704896540
transform 1 0 39836 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1704896540
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1704896540
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1704896540
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_39
timestamp 1704896540
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_51
timestamp 1704896540
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1704896540
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1704896540
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_69
timestamp 1704896540
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_81
timestamp 1704896540
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_93
timestamp 1704896540
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_105
timestamp 1704896540
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1704896540
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_113
timestamp 1704896540
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_125
timestamp 1704896540
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_137
timestamp 1704896540
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_149
timestamp 1704896540
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_161
timestamp 1704896540
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_167
timestamp 1704896540
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_169
timestamp 1704896540
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_181
timestamp 1704896540
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_193
timestamp 1704896540
transform 1 0 18860 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_201
timestamp 1704896540
transform 1 0 19596 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_220
timestamp 1704896540
transform 1 0 21344 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_225
timestamp 1704896540
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_237
timestamp 1704896540
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_249
timestamp 1704896540
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_261
timestamp 1704896540
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_273
timestamp 1704896540
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_279
timestamp 1704896540
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_281
timestamp 1704896540
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_293
timestamp 1704896540
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_305
timestamp 1704896540
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_317
timestamp 1704896540
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_329
timestamp 1704896540
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_335
timestamp 1704896540
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_337
timestamp 1704896540
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_349
timestamp 1704896540
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_361
timestamp 1704896540
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_373
timestamp 1704896540
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_385
timestamp 1704896540
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_391
timestamp 1704896540
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_393
timestamp 1704896540
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_405
timestamp 1704896540
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_417
timestamp 1704896540
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1704896540
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1704896540
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1704896540
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1704896540
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1704896540
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_53
timestamp 1704896540
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_65
timestamp 1704896540
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_77
timestamp 1704896540
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1704896540
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 1704896540
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_97
timestamp 1704896540
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_109
timestamp 1704896540
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_121
timestamp 1704896540
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_133
timestamp 1704896540
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_139
timestamp 1704896540
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_141
timestamp 1704896540
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_153
timestamp 1704896540
transform 1 0 15180 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_168
timestamp 1704896540
transform 1 0 16560 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_180
timestamp 1704896540
transform 1 0 17664 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_192
timestamp 1704896540
transform 1 0 18768 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_197
timestamp 1704896540
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_209
timestamp 1704896540
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_221
timestamp 1704896540
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_233
timestamp 1704896540
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_245
timestamp 1704896540
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_251
timestamp 1704896540
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_253
timestamp 1704896540
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_265
timestamp 1704896540
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_277
timestamp 1704896540
transform 1 0 26588 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_305
timestamp 1704896540
transform 1 0 29164 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_309
timestamp 1704896540
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_321
timestamp 1704896540
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_333
timestamp 1704896540
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_345
timestamp 1704896540
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_357
timestamp 1704896540
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_363
timestamp 1704896540
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_365
timestamp 1704896540
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_377
timestamp 1704896540
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_389
timestamp 1704896540
transform 1 0 36892 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_402
timestamp 1704896540
transform 1 0 38088 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_414
timestamp 1704896540
transform 1 0 39192 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_421
timestamp 1704896540
transform 1 0 39836 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1704896540
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 1704896540
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 1704896540
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_39
timestamp 1704896540
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_51
timestamp 1704896540
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1704896540
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 1704896540
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_69
timestamp 1704896540
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_81
timestamp 1704896540
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_93
timestamp 1704896540
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_105
timestamp 1704896540
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 1704896540
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_113
timestamp 1704896540
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_125
timestamp 1704896540
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_137
timestamp 1704896540
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_149
timestamp 1704896540
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_161
timestamp 1704896540
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_167
timestamp 1704896540
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_169
timestamp 1704896540
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_181
timestamp 1704896540
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_193
timestamp 1704896540
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_205
timestamp 1704896540
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_217
timestamp 1704896540
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_223
timestamp 1704896540
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_225
timestamp 1704896540
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_237
timestamp 1704896540
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_249
timestamp 1704896540
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_261
timestamp 1704896540
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_273
timestamp 1704896540
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_279
timestamp 1704896540
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_281
timestamp 1704896540
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_293
timestamp 1704896540
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_305
timestamp 1704896540
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_317
timestamp 1704896540
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_329
timestamp 1704896540
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_335
timestamp 1704896540
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_337
timestamp 1704896540
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_349
timestamp 1704896540
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_361
timestamp 1704896540
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_373
timestamp 1704896540
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_385
timestamp 1704896540
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_391
timestamp 1704896540
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_393
timestamp 1704896540
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_405
timestamp 1704896540
transform 1 0 38364 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_417
timestamp 1704896540
transform 1 0 39468 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_3
timestamp 1704896540
transform 1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_19
timestamp 1704896540
transform 1 0 2852 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1704896540
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 1704896540
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 1704896540
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_53
timestamp 1704896540
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_65
timestamp 1704896540
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_77
timestamp 1704896540
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 1704896540
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_85
timestamp 1704896540
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_97
timestamp 1704896540
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_109
timestamp 1704896540
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_121
timestamp 1704896540
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_133
timestamp 1704896540
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_139
timestamp 1704896540
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_141
timestamp 1704896540
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_153
timestamp 1704896540
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_165
timestamp 1704896540
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_177
timestamp 1704896540
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_189
timestamp 1704896540
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_195
timestamp 1704896540
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_197
timestamp 1704896540
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_209
timestamp 1704896540
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_221
timestamp 1704896540
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_233
timestamp 1704896540
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_245
timestamp 1704896540
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_251
timestamp 1704896540
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_253
timestamp 1704896540
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_265
timestamp 1704896540
transform 1 0 25484 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_293
timestamp 1704896540
transform 1 0 28060 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_305
timestamp 1704896540
transform 1 0 29164 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_309
timestamp 1704896540
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_321
timestamp 1704896540
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_333
timestamp 1704896540
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_345
timestamp 1704896540
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_357
timestamp 1704896540
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_363
timestamp 1704896540
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_371
timestamp 1704896540
transform 1 0 35236 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_383
timestamp 1704896540
transform 1 0 36340 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_395
timestamp 1704896540
transform 1 0 37444 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_407
timestamp 1704896540
transform 1 0 38548 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_419
timestamp 1704896540
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_421
timestamp 1704896540
transform 1 0 39836 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1704896540
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_15
timestamp 1704896540
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_27
timestamp 1704896540
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_39
timestamp 1704896540
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_51
timestamp 1704896540
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 1704896540
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_57
timestamp 1704896540
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_69
timestamp 1704896540
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_81
timestamp 1704896540
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_93
timestamp 1704896540
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_105
timestamp 1704896540
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_111
timestamp 1704896540
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_113
timestamp 1704896540
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_125
timestamp 1704896540
transform 1 0 12604 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_133
timestamp 1704896540
transform 1 0 13340 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_144
timestamp 1704896540
transform 1 0 14352 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_156
timestamp 1704896540
transform 1 0 15456 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_175
timestamp 1704896540
transform 1 0 17204 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_187
timestamp 1704896540
transform 1 0 18308 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_199
timestamp 1704896540
transform 1 0 19412 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_211
timestamp 1704896540
transform 1 0 20516 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_223
timestamp 1704896540
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_225
timestamp 1704896540
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_237
timestamp 1704896540
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_249
timestamp 1704896540
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_261
timestamp 1704896540
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_273
timestamp 1704896540
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_279
timestamp 1704896540
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_281
timestamp 1704896540
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_293
timestamp 1704896540
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_305
timestamp 1704896540
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_317
timestamp 1704896540
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_329
timestamp 1704896540
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_335
timestamp 1704896540
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_337
timestamp 1704896540
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_349
timestamp 1704896540
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_361
timestamp 1704896540
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_373
timestamp 1704896540
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_385
timestamp 1704896540
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_391
timestamp 1704896540
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_393
timestamp 1704896540
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_405
timestamp 1704896540
transform 1 0 38364 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_417
timestamp 1704896540
transform 1 0 39468 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1704896540
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_15
timestamp 1704896540
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1704896540
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 1704896540
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_41
timestamp 1704896540
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_53
timestamp 1704896540
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_65
timestamp 1704896540
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_77
timestamp 1704896540
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_83
timestamp 1704896540
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_85
timestamp 1704896540
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_97
timestamp 1704896540
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_109
timestamp 1704896540
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_121
timestamp 1704896540
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_133
timestamp 1704896540
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_139
timestamp 1704896540
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_141
timestamp 1704896540
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_153
timestamp 1704896540
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_165
timestamp 1704896540
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_177
timestamp 1704896540
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_189
timestamp 1704896540
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_195
timestamp 1704896540
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_197
timestamp 1704896540
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_209
timestamp 1704896540
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_221
timestamp 1704896540
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_233
timestamp 1704896540
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_245
timestamp 1704896540
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_251
timestamp 1704896540
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_253
timestamp 1704896540
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_265
timestamp 1704896540
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_277
timestamp 1704896540
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_289
timestamp 1704896540
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_301
timestamp 1704896540
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_307
timestamp 1704896540
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_309
timestamp 1704896540
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_321
timestamp 1704896540
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_333
timestamp 1704896540
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_345
timestamp 1704896540
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_357
timestamp 1704896540
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_363
timestamp 1704896540
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_365
timestamp 1704896540
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_377
timestamp 1704896540
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_389
timestamp 1704896540
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_401
timestamp 1704896540
transform 1 0 37996 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_413
timestamp 1704896540
transform 1 0 39100 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_419
timestamp 1704896540
transform 1 0 39652 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_421
timestamp 1704896540
transform 1 0 39836 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_3
timestamp 1704896540
transform 1 0 1380 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_11
timestamp 1704896540
transform 1 0 2116 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_24
timestamp 1704896540
transform 1 0 3312 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_36
timestamp 1704896540
transform 1 0 4416 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_48
timestamp 1704896540
transform 1 0 5520 0 -1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_57
timestamp 1704896540
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_69
timestamp 1704896540
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_81
timestamp 1704896540
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_93
timestamp 1704896540
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_105
timestamp 1704896540
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_111
timestamp 1704896540
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_113
timestamp 1704896540
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_125
timestamp 1704896540
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_137
timestamp 1704896540
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_149
timestamp 1704896540
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_161
timestamp 1704896540
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_167
timestamp 1704896540
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_169
timestamp 1704896540
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_181
timestamp 1704896540
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_193
timestamp 1704896540
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_205
timestamp 1704896540
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_217
timestamp 1704896540
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_223
timestamp 1704896540
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_225
timestamp 1704896540
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_237
timestamp 1704896540
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_249
timestamp 1704896540
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_261
timestamp 1704896540
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_273
timestamp 1704896540
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_279
timestamp 1704896540
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_281
timestamp 1704896540
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_293
timestamp 1704896540
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_305
timestamp 1704896540
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_317
timestamp 1704896540
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_329
timestamp 1704896540
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_335
timestamp 1704896540
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_337
timestamp 1704896540
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_349
timestamp 1704896540
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_361
timestamp 1704896540
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_373
timestamp 1704896540
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_385
timestamp 1704896540
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_391
timestamp 1704896540
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_393
timestamp 1704896540
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_405
timestamp 1704896540
transform 1 0 38364 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_417
timestamp 1704896540
transform 1 0 39468 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_3
timestamp 1704896540
transform 1 0 1380 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_11
timestamp 1704896540
transform 1 0 2116 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_29
timestamp 1704896540
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_41
timestamp 1704896540
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_53
timestamp 1704896540
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_65
timestamp 1704896540
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_77
timestamp 1704896540
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_83
timestamp 1704896540
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_85
timestamp 1704896540
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_97
timestamp 1704896540
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_109
timestamp 1704896540
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_121
timestamp 1704896540
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_133
timestamp 1704896540
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_139
timestamp 1704896540
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_141
timestamp 1704896540
transform 1 0 14076 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_147
timestamp 1704896540
transform 1 0 14628 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_160
timestamp 1704896540
transform 1 0 15824 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_172
timestamp 1704896540
transform 1 0 16928 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_184
timestamp 1704896540
transform 1 0 18032 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_197
timestamp 1704896540
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_209
timestamp 1704896540
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_221
timestamp 1704896540
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_233
timestamp 1704896540
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_245
timestamp 1704896540
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_251
timestamp 1704896540
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_253
timestamp 1704896540
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_265
timestamp 1704896540
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_277
timestamp 1704896540
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_289
timestamp 1704896540
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_301
timestamp 1704896540
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_307
timestamp 1704896540
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_309
timestamp 1704896540
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_321
timestamp 1704896540
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_333
timestamp 1704896540
transform 1 0 31740 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_339
timestamp 1704896540
transform 1 0 32292 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_356
timestamp 1704896540
transform 1 0 33856 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_365
timestamp 1704896540
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_377
timestamp 1704896540
transform 1 0 35788 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_381
timestamp 1704896540
transform 1 0 36156 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_398
timestamp 1704896540
transform 1 0 37720 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_410
timestamp 1704896540
transform 1 0 38824 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_418
timestamp 1704896540
transform 1 0 39560 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_421
timestamp 1704896540
transform 1 0 39836 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 1704896540
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_15
timestamp 1704896540
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_27
timestamp 1704896540
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_39
timestamp 1704896540
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_51
timestamp 1704896540
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_55
timestamp 1704896540
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_57
timestamp 1704896540
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_69
timestamp 1704896540
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_81
timestamp 1704896540
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_93
timestamp 1704896540
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_105
timestamp 1704896540
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_111
timestamp 1704896540
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_113
timestamp 1704896540
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_125
timestamp 1704896540
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_137
timestamp 1704896540
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_149
timestamp 1704896540
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_161
timestamp 1704896540
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_167
timestamp 1704896540
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_169
timestamp 1704896540
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_181
timestamp 1704896540
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_193
timestamp 1704896540
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_205
timestamp 1704896540
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_217
timestamp 1704896540
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_223
timestamp 1704896540
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_225
timestamp 1704896540
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_237
timestamp 1704896540
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_249
timestamp 1704896540
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_261
timestamp 1704896540
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_273
timestamp 1704896540
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_279
timestamp 1704896540
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_281
timestamp 1704896540
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_293
timestamp 1704896540
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_305
timestamp 1704896540
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_317
timestamp 1704896540
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_329
timestamp 1704896540
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_335
timestamp 1704896540
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_337
timestamp 1704896540
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_349
timestamp 1704896540
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_361
timestamp 1704896540
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_373
timestamp 1704896540
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_385
timestamp 1704896540
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_391
timestamp 1704896540
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_393
timestamp 1704896540
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_405
timestamp 1704896540
transform 1 0 38364 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_417
timestamp 1704896540
transform 1 0 39468 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 1704896540
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_15
timestamp 1704896540
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 1704896540
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_29
timestamp 1704896540
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_41
timestamp 1704896540
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_53
timestamp 1704896540
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_65
timestamp 1704896540
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_77
timestamp 1704896540
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_83
timestamp 1704896540
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_85
timestamp 1704896540
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_97
timestamp 1704896540
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_109
timestamp 1704896540
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_121
timestamp 1704896540
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_133
timestamp 1704896540
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_139
timestamp 1704896540
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_141
timestamp 1704896540
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_153
timestamp 1704896540
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_177
timestamp 1704896540
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_189
timestamp 1704896540
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_195
timestamp 1704896540
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_197
timestamp 1704896540
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_209
timestamp 1704896540
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_221
timestamp 1704896540
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_233
timestamp 1704896540
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_245
timestamp 1704896540
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_251
timestamp 1704896540
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_253
timestamp 1704896540
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_265
timestamp 1704896540
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_277
timestamp 1704896540
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_289
timestamp 1704896540
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_301
timestamp 1704896540
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_307
timestamp 1704896540
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_309
timestamp 1704896540
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_321
timestamp 1704896540
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_333
timestamp 1704896540
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_345
timestamp 1704896540
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_357
timestamp 1704896540
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_363
timestamp 1704896540
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_365
timestamp 1704896540
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_377
timestamp 1704896540
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_389
timestamp 1704896540
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_401
timestamp 1704896540
transform 1 0 37996 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_413
timestamp 1704896540
transform 1 0 39100 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_419
timestamp 1704896540
transform 1 0 39652 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_421
timestamp 1704896540
transform 1 0 39836 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 1704896540
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_15
timestamp 1704896540
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_27
timestamp 1704896540
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_39
timestamp 1704896540
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_51
timestamp 1704896540
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_55
timestamp 1704896540
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_57
timestamp 1704896540
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_69
timestamp 1704896540
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_81
timestamp 1704896540
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_93
timestamp 1704896540
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_105
timestamp 1704896540
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_111
timestamp 1704896540
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_113
timestamp 1704896540
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_125
timestamp 1704896540
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_137
timestamp 1704896540
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_149
timestamp 1704896540
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_161
timestamp 1704896540
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_167
timestamp 1704896540
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_169
timestamp 1704896540
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_181
timestamp 1704896540
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_193
timestamp 1704896540
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_205
timestamp 1704896540
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_217
timestamp 1704896540
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_223
timestamp 1704896540
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_225
timestamp 1704896540
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_237
timestamp 1704896540
transform 1 0 22908 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_243
timestamp 1704896540
transform 1 0 23460 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_255
timestamp 1704896540
transform 1 0 24564 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_267
timestamp 1704896540
transform 1 0 25668 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_279
timestamp 1704896540
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_281
timestamp 1704896540
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_293
timestamp 1704896540
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_305
timestamp 1704896540
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_317
timestamp 1704896540
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_329
timestamp 1704896540
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_335
timestamp 1704896540
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_337
timestamp 1704896540
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_349
timestamp 1704896540
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_361
timestamp 1704896540
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_373
timestamp 1704896540
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_385
timestamp 1704896540
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_391
timestamp 1704896540
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_393
timestamp 1704896540
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_405
timestamp 1704896540
transform 1 0 38364 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_411
timestamp 1704896540
transform 1 0 38916 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_414
timestamp 1704896540
transform 1 0 39192 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_426
timestamp 1704896540
transform 1 0 40296 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_3
timestamp 1704896540
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_15
timestamp 1704896540
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1704896540
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_29
timestamp 1704896540
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_41
timestamp 1704896540
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_53
timestamp 1704896540
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_65
timestamp 1704896540
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_77
timestamp 1704896540
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_83
timestamp 1704896540
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_85
timestamp 1704896540
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_97
timestamp 1704896540
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_109
timestamp 1704896540
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_121
timestamp 1704896540
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_133
timestamp 1704896540
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_139
timestamp 1704896540
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_141
timestamp 1704896540
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_153
timestamp 1704896540
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_165
timestamp 1704896540
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_177
timestamp 1704896540
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_189
timestamp 1704896540
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_195
timestamp 1704896540
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_197
timestamp 1704896540
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_209
timestamp 1704896540
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_221
timestamp 1704896540
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_233
timestamp 1704896540
transform 1 0 22540 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_245
timestamp 1704896540
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_251
timestamp 1704896540
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_253
timestamp 1704896540
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_265
timestamp 1704896540
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_277
timestamp 1704896540
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_289
timestamp 1704896540
transform 1 0 27692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_301
timestamp 1704896540
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_307
timestamp 1704896540
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_309
timestamp 1704896540
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_321
timestamp 1704896540
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_333
timestamp 1704896540
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_345
timestamp 1704896540
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_357
timestamp 1704896540
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_363
timestamp 1704896540
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_365
timestamp 1704896540
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_377
timestamp 1704896540
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_389
timestamp 1704896540
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_401
timestamp 1704896540
transform 1 0 37996 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_409
timestamp 1704896540
transform 1 0 38732 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_421
timestamp 1704896540
transform 1 0 39836 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_23
timestamp 1704896540
transform 1 0 3220 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_35
timestamp 1704896540
transform 1 0 4324 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_47
timestamp 1704896540
transform 1 0 5428 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_55
timestamp 1704896540
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_57
timestamp 1704896540
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_69
timestamp 1704896540
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_81
timestamp 1704896540
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_93
timestamp 1704896540
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_105
timestamp 1704896540
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_111
timestamp 1704896540
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_113
timestamp 1704896540
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_125
timestamp 1704896540
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_137
timestamp 1704896540
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_149
timestamp 1704896540
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_161
timestamp 1704896540
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_167
timestamp 1704896540
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_169
timestamp 1704896540
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_181
timestamp 1704896540
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_193
timestamp 1704896540
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_205
timestamp 1704896540
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_217
timestamp 1704896540
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_223
timestamp 1704896540
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_225
timestamp 1704896540
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_237
timestamp 1704896540
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_249
timestamp 1704896540
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_261
timestamp 1704896540
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_273
timestamp 1704896540
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_279
timestamp 1704896540
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_281
timestamp 1704896540
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_293
timestamp 1704896540
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_305
timestamp 1704896540
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_317
timestamp 1704896540
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_329
timestamp 1704896540
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_335
timestamp 1704896540
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_337
timestamp 1704896540
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_349
timestamp 1704896540
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_361
timestamp 1704896540
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_373
timestamp 1704896540
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_385
timestamp 1704896540
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_391
timestamp 1704896540
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_393
timestamp 1704896540
transform 1 0 37260 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_410
timestamp 1704896540
transform 1 0 38824 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_414
timestamp 1704896540
transform 1 0 39192 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_3
timestamp 1704896540
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_15
timestamp 1704896540
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 1704896540
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_29
timestamp 1704896540
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_41
timestamp 1704896540
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_53
timestamp 1704896540
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_65
timestamp 1704896540
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_77
timestamp 1704896540
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_83
timestamp 1704896540
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_85
timestamp 1704896540
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_97
timestamp 1704896540
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_109
timestamp 1704896540
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_121
timestamp 1704896540
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_133
timestamp 1704896540
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_139
timestamp 1704896540
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_141
timestamp 1704896540
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_153
timestamp 1704896540
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_165
timestamp 1704896540
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_177
timestamp 1704896540
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_189
timestamp 1704896540
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_195
timestamp 1704896540
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_197
timestamp 1704896540
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_209
timestamp 1704896540
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_221
timestamp 1704896540
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_233
timestamp 1704896540
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_245
timestamp 1704896540
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_251
timestamp 1704896540
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_253
timestamp 1704896540
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_265
timestamp 1704896540
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_277
timestamp 1704896540
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_289
timestamp 1704896540
transform 1 0 27692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_301
timestamp 1704896540
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_307
timestamp 1704896540
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_309
timestamp 1704896540
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_321
timestamp 1704896540
transform 1 0 30636 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_345
timestamp 1704896540
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_357
timestamp 1704896540
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_363
timestamp 1704896540
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_365
timestamp 1704896540
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_377
timestamp 1704896540
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_389
timestamp 1704896540
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_401
timestamp 1704896540
transform 1 0 37996 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_407
timestamp 1704896540
transform 1 0 38548 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_410
timestamp 1704896540
transform 1 0 38824 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_419
timestamp 1704896540
transform 1 0 39652 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_421
timestamp 1704896540
transform 1 0 39836 0 1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_3
timestamp 1704896540
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_15
timestamp 1704896540
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_27
timestamp 1704896540
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_39
timestamp 1704896540
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_51
timestamp 1704896540
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_55
timestamp 1704896540
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_57
timestamp 1704896540
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_69
timestamp 1704896540
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_81
timestamp 1704896540
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_93
timestamp 1704896540
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_105
timestamp 1704896540
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_111
timestamp 1704896540
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_113
timestamp 1704896540
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_125
timestamp 1704896540
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_137
timestamp 1704896540
transform 1 0 13708 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_145
timestamp 1704896540
transform 1 0 14444 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_160
timestamp 1704896540
transform 1 0 15824 0 -1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_169
timestamp 1704896540
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_181
timestamp 1704896540
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_193
timestamp 1704896540
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_205
timestamp 1704896540
transform 1 0 19964 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_217
timestamp 1704896540
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_223
timestamp 1704896540
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_225
timestamp 1704896540
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_237
timestamp 1704896540
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_249
timestamp 1704896540
transform 1 0 24012 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_261
timestamp 1704896540
transform 1 0 25116 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_273
timestamp 1704896540
transform 1 0 26220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_279
timestamp 1704896540
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_281
timestamp 1704896540
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_293
timestamp 1704896540
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_305
timestamp 1704896540
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_317
timestamp 1704896540
transform 1 0 30268 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_334
timestamp 1704896540
transform 1 0 31832 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_337
timestamp 1704896540
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_349
timestamp 1704896540
transform 1 0 33212 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_353
timestamp 1704896540
transform 1 0 33580 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_375
timestamp 1704896540
transform 1 0 35604 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_387
timestamp 1704896540
transform 1 0 36708 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_391
timestamp 1704896540
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_393
timestamp 1704896540
transform 1 0 37260 0 -1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_408
timestamp 1704896540
transform 1 0 38640 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_420
timestamp 1704896540
transform 1 0 39744 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_428
timestamp 1704896540
transform 1 0 40480 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_3
timestamp 1704896540
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_15
timestamp 1704896540
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_27
timestamp 1704896540
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_29
timestamp 1704896540
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_41
timestamp 1704896540
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_53
timestamp 1704896540
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_65
timestamp 1704896540
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_77
timestamp 1704896540
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_83
timestamp 1704896540
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_85
timestamp 1704896540
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_97
timestamp 1704896540
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_109
timestamp 1704896540
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_121
timestamp 1704896540
transform 1 0 12236 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_125
timestamp 1704896540
transform 1 0 12604 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_135
timestamp 1704896540
transform 1 0 13524 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_139
timestamp 1704896540
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_141
timestamp 1704896540
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_153
timestamp 1704896540
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_165
timestamp 1704896540
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_177
timestamp 1704896540
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_189
timestamp 1704896540
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_195
timestamp 1704896540
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_197
timestamp 1704896540
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_209
timestamp 1704896540
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_221
timestamp 1704896540
transform 1 0 21436 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_233
timestamp 1704896540
transform 1 0 22540 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_245
timestamp 1704896540
transform 1 0 23644 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_251
timestamp 1704896540
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_253
timestamp 1704896540
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_265
timestamp 1704896540
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_277
timestamp 1704896540
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_289
timestamp 1704896540
transform 1 0 27692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_301
timestamp 1704896540
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_307
timestamp 1704896540
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_309
timestamp 1704896540
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_321
timestamp 1704896540
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_333
timestamp 1704896540
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_345
timestamp 1704896540
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_357
timestamp 1704896540
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_363
timestamp 1704896540
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_377
timestamp 1704896540
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_389
timestamp 1704896540
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_401
timestamp 1704896540
transform 1 0 37996 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_413
timestamp 1704896540
transform 1 0 39100 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_419
timestamp 1704896540
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_421
timestamp 1704896540
transform 1 0 39836 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_3
timestamp 1704896540
transform 1 0 1380 0 -1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_17
timestamp 1704896540
transform 1 0 2668 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_29
timestamp 1704896540
transform 1 0 3772 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_41
timestamp 1704896540
transform 1 0 4876 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_53
timestamp 1704896540
transform 1 0 5980 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_57
timestamp 1704896540
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_69
timestamp 1704896540
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_81
timestamp 1704896540
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_93
timestamp 1704896540
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_105
timestamp 1704896540
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_111
timestamp 1704896540
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_113
timestamp 1704896540
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_125
timestamp 1704896540
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_137
timestamp 1704896540
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_149
timestamp 1704896540
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_161
timestamp 1704896540
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_167
timestamp 1704896540
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_169
timestamp 1704896540
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_181
timestamp 1704896540
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_193
timestamp 1704896540
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_205
timestamp 1704896540
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_217
timestamp 1704896540
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_223
timestamp 1704896540
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_225
timestamp 1704896540
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_237
timestamp 1704896540
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_249
timestamp 1704896540
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_261
timestamp 1704896540
transform 1 0 25116 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_273
timestamp 1704896540
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_279
timestamp 1704896540
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_281
timestamp 1704896540
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_293
timestamp 1704896540
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_305
timestamp 1704896540
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_317
timestamp 1704896540
transform 1 0 30268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_329
timestamp 1704896540
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_335
timestamp 1704896540
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_337
timestamp 1704896540
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_349
timestamp 1704896540
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_361
timestamp 1704896540
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_373
timestamp 1704896540
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_385
timestamp 1704896540
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_391
timestamp 1704896540
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_393
timestamp 1704896540
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_405
timestamp 1704896540
transform 1 0 38364 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_417
timestamp 1704896540
transform 1 0 39468 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_3
timestamp 1704896540
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_15
timestamp 1704896540
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_27
timestamp 1704896540
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_29
timestamp 1704896540
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_41
timestamp 1704896540
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_53
timestamp 1704896540
transform 1 0 5980 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_66
timestamp 1704896540
transform 1 0 7176 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_78
timestamp 1704896540
transform 1 0 8280 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_85
timestamp 1704896540
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_97
timestamp 1704896540
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_109
timestamp 1704896540
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_121
timestamp 1704896540
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_133
timestamp 1704896540
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_139
timestamp 1704896540
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_141
timestamp 1704896540
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_153
timestamp 1704896540
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_165
timestamp 1704896540
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_177
timestamp 1704896540
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_189
timestamp 1704896540
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_195
timestamp 1704896540
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_197
timestamp 1704896540
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_209
timestamp 1704896540
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_221
timestamp 1704896540
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_233
timestamp 1704896540
transform 1 0 22540 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_245
timestamp 1704896540
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_251
timestamp 1704896540
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_253
timestamp 1704896540
transform 1 0 24380 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_261
timestamp 1704896540
transform 1 0 25116 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_273
timestamp 1704896540
transform 1 0 26220 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_285
timestamp 1704896540
transform 1 0 27324 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_297
timestamp 1704896540
transform 1 0 28428 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_305
timestamp 1704896540
transform 1 0 29164 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_309
timestamp 1704896540
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_321
timestamp 1704896540
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_333
timestamp 1704896540
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_345
timestamp 1704896540
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_357
timestamp 1704896540
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_363
timestamp 1704896540
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_365
timestamp 1704896540
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_377
timestamp 1704896540
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_389
timestamp 1704896540
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_401
timestamp 1704896540
transform 1 0 37996 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_413
timestamp 1704896540
transform 1 0 39100 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_419
timestamp 1704896540
transform 1 0 39652 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_421
timestamp 1704896540
transform 1 0 39836 0 1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_3
timestamp 1704896540
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_15
timestamp 1704896540
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_27
timestamp 1704896540
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_39
timestamp 1704896540
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_51
timestamp 1704896540
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_55
timestamp 1704896540
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_57
timestamp 1704896540
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_69
timestamp 1704896540
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_81
timestamp 1704896540
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_93
timestamp 1704896540
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_105
timestamp 1704896540
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_111
timestamp 1704896540
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_113
timestamp 1704896540
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_125
timestamp 1704896540
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_137
timestamp 1704896540
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_149
timestamp 1704896540
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_161
timestamp 1704896540
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_167
timestamp 1704896540
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_169
timestamp 1704896540
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_181
timestamp 1704896540
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_193
timestamp 1704896540
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_205
timestamp 1704896540
transform 1 0 19964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_217
timestamp 1704896540
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_223
timestamp 1704896540
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_225
timestamp 1704896540
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_237
timestamp 1704896540
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_249
timestamp 1704896540
transform 1 0 24012 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_261
timestamp 1704896540
transform 1 0 25116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_273
timestamp 1704896540
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_279
timestamp 1704896540
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_281
timestamp 1704896540
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_293
timestamp 1704896540
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_305
timestamp 1704896540
transform 1 0 29164 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_317
timestamp 1704896540
transform 1 0 30268 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_329
timestamp 1704896540
transform 1 0 31372 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_335
timestamp 1704896540
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_337
timestamp 1704896540
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_349
timestamp 1704896540
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_361
timestamp 1704896540
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_373
timestamp 1704896540
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_385
timestamp 1704896540
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_391
timestamp 1704896540
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_393
timestamp 1704896540
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_405
timestamp 1704896540
transform 1 0 38364 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_417
timestamp 1704896540
transform 1 0 39468 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_3
timestamp 1704896540
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_15
timestamp 1704896540
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_27
timestamp 1704896540
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_29
timestamp 1704896540
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_41
timestamp 1704896540
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_53
timestamp 1704896540
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_65
timestamp 1704896540
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_77
timestamp 1704896540
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_83
timestamp 1704896540
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_85
timestamp 1704896540
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_97
timestamp 1704896540
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_109
timestamp 1704896540
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_121
timestamp 1704896540
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_133
timestamp 1704896540
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_139
timestamp 1704896540
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_141
timestamp 1704896540
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_153
timestamp 1704896540
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_165
timestamp 1704896540
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_177
timestamp 1704896540
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_189
timestamp 1704896540
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_195
timestamp 1704896540
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_197
timestamp 1704896540
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_209
timestamp 1704896540
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_221
timestamp 1704896540
transform 1 0 21436 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_233
timestamp 1704896540
transform 1 0 22540 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_245
timestamp 1704896540
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_251
timestamp 1704896540
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_253
timestamp 1704896540
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_265
timestamp 1704896540
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_277
timestamp 1704896540
transform 1 0 26588 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_289
timestamp 1704896540
transform 1 0 27692 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_301
timestamp 1704896540
transform 1 0 28796 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_307
timestamp 1704896540
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_309
timestamp 1704896540
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_321
timestamp 1704896540
transform 1 0 30636 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_333
timestamp 1704896540
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_345
timestamp 1704896540
transform 1 0 32844 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_357
timestamp 1704896540
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_363
timestamp 1704896540
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_365
timestamp 1704896540
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_377
timestamp 1704896540
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_389
timestamp 1704896540
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_401
timestamp 1704896540
transform 1 0 37996 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_407
timestamp 1704896540
transform 1 0 38548 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_415
timestamp 1704896540
transform 1 0 39284 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_419
timestamp 1704896540
transform 1 0 39652 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_421
timestamp 1704896540
transform 1 0 39836 0 1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_3
timestamp 1704896540
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_15
timestamp 1704896540
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_27
timestamp 1704896540
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_39
timestamp 1704896540
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_51
timestamp 1704896540
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_55
timestamp 1704896540
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_57
timestamp 1704896540
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_69
timestamp 1704896540
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_81
timestamp 1704896540
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_93
timestamp 1704896540
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_105
timestamp 1704896540
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_111
timestamp 1704896540
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_113
timestamp 1704896540
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_125
timestamp 1704896540
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_137
timestamp 1704896540
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_149
timestamp 1704896540
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_161
timestamp 1704896540
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_167
timestamp 1704896540
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_169
timestamp 1704896540
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_181
timestamp 1704896540
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_193
timestamp 1704896540
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_205
timestamp 1704896540
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_217
timestamp 1704896540
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_223
timestamp 1704896540
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_225
timestamp 1704896540
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_237
timestamp 1704896540
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_249
timestamp 1704896540
transform 1 0 24012 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_261
timestamp 1704896540
transform 1 0 25116 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_273
timestamp 1704896540
transform 1 0 26220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_279
timestamp 1704896540
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_281
timestamp 1704896540
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_293
timestamp 1704896540
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_305
timestamp 1704896540
transform 1 0 29164 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_321
timestamp 1704896540
transform 1 0 30636 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_333
timestamp 1704896540
transform 1 0 31740 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_337
timestamp 1704896540
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_349
timestamp 1704896540
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_361
timestamp 1704896540
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_373
timestamp 1704896540
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_385
timestamp 1704896540
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_391
timestamp 1704896540
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_393
timestamp 1704896540
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_405
timestamp 1704896540
transform 1 0 38364 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_417
timestamp 1704896540
transform 1 0 39468 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_3
timestamp 1704896540
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_15
timestamp 1704896540
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_27
timestamp 1704896540
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_29
timestamp 1704896540
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_41
timestamp 1704896540
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_53
timestamp 1704896540
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_65
timestamp 1704896540
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_77
timestamp 1704896540
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_83
timestamp 1704896540
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_85
timestamp 1704896540
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_97
timestamp 1704896540
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_109
timestamp 1704896540
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_121
timestamp 1704896540
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_133
timestamp 1704896540
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_139
timestamp 1704896540
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_141
timestamp 1704896540
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_153
timestamp 1704896540
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_165
timestamp 1704896540
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_177
timestamp 1704896540
transform 1 0 17388 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_194
timestamp 1704896540
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_201
timestamp 1704896540
transform 1 0 19596 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_213
timestamp 1704896540
transform 1 0 20700 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_225
timestamp 1704896540
transform 1 0 21804 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_237
timestamp 1704896540
transform 1 0 22908 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_249
timestamp 1704896540
transform 1 0 24012 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_253
timestamp 1704896540
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_265
timestamp 1704896540
transform 1 0 25484 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_282
timestamp 1704896540
transform 1 0 27048 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_294
timestamp 1704896540
transform 1 0 28152 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_306
timestamp 1704896540
transform 1 0 29256 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_309
timestamp 1704896540
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_321
timestamp 1704896540
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_333
timestamp 1704896540
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_345
timestamp 1704896540
transform 1 0 32844 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_357
timestamp 1704896540
transform 1 0 33948 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_363
timestamp 1704896540
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_365
timestamp 1704896540
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_377
timestamp 1704896540
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_389
timestamp 1704896540
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_401
timestamp 1704896540
transform 1 0 37996 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_413
timestamp 1704896540
transform 1 0 39100 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_419
timestamp 1704896540
transform 1 0 39652 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_421
timestamp 1704896540
transform 1 0 39836 0 1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_3
timestamp 1704896540
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_15
timestamp 1704896540
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_27
timestamp 1704896540
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_39
timestamp 1704896540
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_51
timestamp 1704896540
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_55
timestamp 1704896540
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_57
timestamp 1704896540
transform 1 0 6348 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_74
timestamp 1704896540
transform 1 0 7912 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_86
timestamp 1704896540
transform 1 0 9016 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_98
timestamp 1704896540
transform 1 0 10120 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_110
timestamp 1704896540
transform 1 0 11224 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_113
timestamp 1704896540
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_125
timestamp 1704896540
transform 1 0 12604 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_138
timestamp 1704896540
transform 1 0 13800 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_150
timestamp 1704896540
transform 1 0 14904 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_162
timestamp 1704896540
transform 1 0 16008 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_169
timestamp 1704896540
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_181
timestamp 1704896540
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_193
timestamp 1704896540
transform 1 0 18860 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_205
timestamp 1704896540
transform 1 0 19964 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_217
timestamp 1704896540
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_223
timestamp 1704896540
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_225
timestamp 1704896540
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_237
timestamp 1704896540
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_249
timestamp 1704896540
transform 1 0 24012 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_261
timestamp 1704896540
transform 1 0 25116 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_273
timestamp 1704896540
transform 1 0 26220 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_279
timestamp 1704896540
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_281
timestamp 1704896540
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_293
timestamp 1704896540
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_305
timestamp 1704896540
transform 1 0 29164 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_317
timestamp 1704896540
transform 1 0 30268 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_329
timestamp 1704896540
transform 1 0 31372 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_335
timestamp 1704896540
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_337
timestamp 1704896540
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_349
timestamp 1704896540
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_361
timestamp 1704896540
transform 1 0 34316 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_373
timestamp 1704896540
transform 1 0 35420 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_385
timestamp 1704896540
transform 1 0 36524 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_391
timestamp 1704896540
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_393
timestamp 1704896540
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_405
timestamp 1704896540
transform 1 0 38364 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_417
timestamp 1704896540
transform 1 0 39468 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_3
timestamp 1704896540
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_15
timestamp 1704896540
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_27
timestamp 1704896540
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_38
timestamp 1704896540
transform 1 0 4600 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_50
timestamp 1704896540
transform 1 0 5704 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_62
timestamp 1704896540
transform 1 0 6808 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_71
timestamp 1704896540
transform 1 0 7636 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_83
timestamp 1704896540
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_85
timestamp 1704896540
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_97
timestamp 1704896540
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_109
timestamp 1704896540
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_121
timestamp 1704896540
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_133
timestamp 1704896540
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_139
timestamp 1704896540
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_141
timestamp 1704896540
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_153
timestamp 1704896540
transform 1 0 15180 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_175
timestamp 1704896540
transform 1 0 17204 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_187
timestamp 1704896540
transform 1 0 18308 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_195
timestamp 1704896540
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_197
timestamp 1704896540
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_209
timestamp 1704896540
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_221
timestamp 1704896540
transform 1 0 21436 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_233
timestamp 1704896540
transform 1 0 22540 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_245
timestamp 1704896540
transform 1 0 23644 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_251
timestamp 1704896540
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_253
timestamp 1704896540
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_265
timestamp 1704896540
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_277
timestamp 1704896540
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_289
timestamp 1704896540
transform 1 0 27692 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_301
timestamp 1704896540
transform 1 0 28796 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_307
timestamp 1704896540
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_309
timestamp 1704896540
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_321
timestamp 1704896540
transform 1 0 30636 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_333
timestamp 1704896540
transform 1 0 31740 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_341
timestamp 1704896540
transform 1 0 32476 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_365
timestamp 1704896540
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_377
timestamp 1704896540
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_389
timestamp 1704896540
transform 1 0 36892 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_393
timestamp 1704896540
transform 1 0 37260 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_406
timestamp 1704896540
transform 1 0 38456 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_418
timestamp 1704896540
transform 1 0 39560 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_421
timestamp 1704896540
transform 1 0 39836 0 1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_10
timestamp 1704896540
transform 1 0 2024 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_22
timestamp 1704896540
transform 1 0 3128 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_34
timestamp 1704896540
transform 1 0 4232 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_46
timestamp 1704896540
transform 1 0 5336 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_54
timestamp 1704896540
transform 1 0 6072 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_57
timestamp 1704896540
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_69
timestamp 1704896540
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_81
timestamp 1704896540
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_93
timestamp 1704896540
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_105
timestamp 1704896540
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_111
timestamp 1704896540
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_113
timestamp 1704896540
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_125
timestamp 1704896540
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_137
timestamp 1704896540
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_149
timestamp 1704896540
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_161
timestamp 1704896540
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_167
timestamp 1704896540
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_169
timestamp 1704896540
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_181
timestamp 1704896540
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_193
timestamp 1704896540
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_205
timestamp 1704896540
transform 1 0 19964 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_217
timestamp 1704896540
transform 1 0 21068 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_223
timestamp 1704896540
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_225
timestamp 1704896540
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_237
timestamp 1704896540
transform 1 0 22908 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_249
timestamp 1704896540
transform 1 0 24012 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_270
timestamp 1704896540
transform 1 0 25944 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_278
timestamp 1704896540
transform 1 0 26680 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_281
timestamp 1704896540
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_293
timestamp 1704896540
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_305
timestamp 1704896540
transform 1 0 29164 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_317
timestamp 1704896540
transform 1 0 30268 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_329
timestamp 1704896540
transform 1 0 31372 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_335
timestamp 1704896540
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_337
timestamp 1704896540
transform 1 0 32108 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_345
timestamp 1704896540
transform 1 0 32844 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_352
timestamp 1704896540
transform 1 0 33488 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_364
timestamp 1704896540
transform 1 0 34592 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_376
timestamp 1704896540
transform 1 0 35696 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_388
timestamp 1704896540
transform 1 0 36800 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_393
timestamp 1704896540
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_405
timestamp 1704896540
transform 1 0 38364 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_417
timestamp 1704896540
transform 1 0 39468 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_3
timestamp 1704896540
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_15
timestamp 1704896540
transform 1 0 2484 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_27
timestamp 1704896540
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_29
timestamp 1704896540
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_41
timestamp 1704896540
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_53
timestamp 1704896540
transform 1 0 5980 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_61
timestamp 1704896540
transform 1 0 6716 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_76
timestamp 1704896540
transform 1 0 8096 0 1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_85
timestamp 1704896540
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_97
timestamp 1704896540
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_109
timestamp 1704896540
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_121
timestamp 1704896540
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_133
timestamp 1704896540
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_139
timestamp 1704896540
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_141
timestamp 1704896540
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_153
timestamp 1704896540
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_165
timestamp 1704896540
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_177
timestamp 1704896540
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_189
timestamp 1704896540
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_195
timestamp 1704896540
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_197
timestamp 1704896540
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_209
timestamp 1704896540
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_221
timestamp 1704896540
transform 1 0 21436 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_239
timestamp 1704896540
transform 1 0 23092 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_251
timestamp 1704896540
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_253
timestamp 1704896540
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_265
timestamp 1704896540
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_277
timestamp 1704896540
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_289
timestamp 1704896540
transform 1 0 27692 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_301
timestamp 1704896540
transform 1 0 28796 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_307
timestamp 1704896540
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_309
timestamp 1704896540
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_321
timestamp 1704896540
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_333
timestamp 1704896540
transform 1 0 31740 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_345
timestamp 1704896540
transform 1 0 32844 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_357
timestamp 1704896540
transform 1 0 33948 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_363
timestamp 1704896540
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_365
timestamp 1704896540
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_377
timestamp 1704896540
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_389
timestamp 1704896540
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_401
timestamp 1704896540
transform 1 0 37996 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_413
timestamp 1704896540
transform 1 0 39100 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_419
timestamp 1704896540
transform 1 0 39652 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_421
timestamp 1704896540
transform 1 0 39836 0 1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_3
timestamp 1704896540
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_15
timestamp 1704896540
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_27
timestamp 1704896540
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_39
timestamp 1704896540
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_51
timestamp 1704896540
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_55
timestamp 1704896540
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_57
timestamp 1704896540
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_69
timestamp 1704896540
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_81
timestamp 1704896540
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_93
timestamp 1704896540
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_105
timestamp 1704896540
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_111
timestamp 1704896540
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_113
timestamp 1704896540
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_125
timestamp 1704896540
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_137
timestamp 1704896540
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_149
timestamp 1704896540
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_161
timestamp 1704896540
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_167
timestamp 1704896540
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_169
timestamp 1704896540
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_181
timestamp 1704896540
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_193
timestamp 1704896540
transform 1 0 18860 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_205
timestamp 1704896540
transform 1 0 19964 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_217
timestamp 1704896540
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_223
timestamp 1704896540
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_225
timestamp 1704896540
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_237
timestamp 1704896540
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_249
timestamp 1704896540
transform 1 0 24012 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_261
timestamp 1704896540
transform 1 0 25116 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_273
timestamp 1704896540
transform 1 0 26220 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_279
timestamp 1704896540
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_281
timestamp 1704896540
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_293
timestamp 1704896540
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_305
timestamp 1704896540
transform 1 0 29164 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_317
timestamp 1704896540
transform 1 0 30268 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_329
timestamp 1704896540
transform 1 0 31372 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_335
timestamp 1704896540
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_337
timestamp 1704896540
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_349
timestamp 1704896540
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_361
timestamp 1704896540
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_373
timestamp 1704896540
transform 1 0 35420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_385
timestamp 1704896540
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_391
timestamp 1704896540
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_393
timestamp 1704896540
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_405
timestamp 1704896540
transform 1 0 38364 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_417
timestamp 1704896540
transform 1 0 39468 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_3
timestamp 1704896540
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_15
timestamp 1704896540
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_27
timestamp 1704896540
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_29
timestamp 1704896540
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_41
timestamp 1704896540
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_53
timestamp 1704896540
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_65
timestamp 1704896540
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_77
timestamp 1704896540
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_83
timestamp 1704896540
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_85
timestamp 1704896540
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_97
timestamp 1704896540
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_109
timestamp 1704896540
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_121
timestamp 1704896540
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_133
timestamp 1704896540
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_139
timestamp 1704896540
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_141
timestamp 1704896540
transform 1 0 14076 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_147
timestamp 1704896540
transform 1 0 14628 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_156
timestamp 1704896540
transform 1 0 15456 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_168
timestamp 1704896540
transform 1 0 16560 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_180
timestamp 1704896540
transform 1 0 17664 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_192
timestamp 1704896540
transform 1 0 18768 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_197
timestamp 1704896540
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_209
timestamp 1704896540
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_221
timestamp 1704896540
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_233
timestamp 1704896540
transform 1 0 22540 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_245
timestamp 1704896540
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_251
timestamp 1704896540
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_253
timestamp 1704896540
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_265
timestamp 1704896540
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_277
timestamp 1704896540
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_289
timestamp 1704896540
transform 1 0 27692 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_301
timestamp 1704896540
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_307
timestamp 1704896540
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_309
timestamp 1704896540
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_321
timestamp 1704896540
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_333
timestamp 1704896540
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_345
timestamp 1704896540
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_357
timestamp 1704896540
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_363
timestamp 1704896540
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_365
timestamp 1704896540
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_377
timestamp 1704896540
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_389
timestamp 1704896540
transform 1 0 36892 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_401
timestamp 1704896540
transform 1 0 37996 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_413
timestamp 1704896540
transform 1 0 39100 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_419
timestamp 1704896540
transform 1 0 39652 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_421
timestamp 1704896540
transform 1 0 39836 0 1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_9
timestamp 1704896540
transform 1 0 1932 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_21
timestamp 1704896540
transform 1 0 3036 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_33
timestamp 1704896540
transform 1 0 4140 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_45
timestamp 1704896540
transform 1 0 5244 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_53
timestamp 1704896540
transform 1 0 5980 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_57
timestamp 1704896540
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_69
timestamp 1704896540
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_81
timestamp 1704896540
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_93
timestamp 1704896540
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_105
timestamp 1704896540
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_111
timestamp 1704896540
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_122
timestamp 1704896540
transform 1 0 12328 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_134
timestamp 1704896540
transform 1 0 13432 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_142
timestamp 1704896540
transform 1 0 14168 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_152
timestamp 1704896540
transform 1 0 15088 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_164
timestamp 1704896540
transform 1 0 16192 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_200
timestamp 1704896540
transform 1 0 19504 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_212
timestamp 1704896540
transform 1 0 20608 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_225
timestamp 1704896540
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_237
timestamp 1704896540
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_249
timestamp 1704896540
transform 1 0 24012 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_261
timestamp 1704896540
transform 1 0 25116 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_273
timestamp 1704896540
transform 1 0 26220 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_279
timestamp 1704896540
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_281
timestamp 1704896540
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_293
timestamp 1704896540
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_305
timestamp 1704896540
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_317
timestamp 1704896540
transform 1 0 30268 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_329
timestamp 1704896540
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_335
timestamp 1704896540
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_337
timestamp 1704896540
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_349
timestamp 1704896540
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_361
timestamp 1704896540
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_373
timestamp 1704896540
transform 1 0 35420 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_385
timestamp 1704896540
transform 1 0 36524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_391
timestamp 1704896540
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_393
timestamp 1704896540
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_405
timestamp 1704896540
transform 1 0 38364 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_3
timestamp 1704896540
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_15
timestamp 1704896540
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_27
timestamp 1704896540
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_29
timestamp 1704896540
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_41
timestamp 1704896540
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_53
timestamp 1704896540
transform 1 0 5980 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_57
timestamp 1704896540
transform 1 0 6348 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_70
timestamp 1704896540
transform 1 0 7544 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_81
timestamp 1704896540
transform 1 0 8556 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_85
timestamp 1704896540
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_97
timestamp 1704896540
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_109
timestamp 1704896540
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_121
timestamp 1704896540
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_133
timestamp 1704896540
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_139
timestamp 1704896540
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_141
timestamp 1704896540
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_153
timestamp 1704896540
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_165
timestamp 1704896540
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_177
timestamp 1704896540
transform 1 0 17388 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_189
timestamp 1704896540
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_195
timestamp 1704896540
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_197
timestamp 1704896540
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_209
timestamp 1704896540
transform 1 0 20332 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_220
timestamp 1704896540
transform 1 0 21344 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_232
timestamp 1704896540
transform 1 0 22448 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_244
timestamp 1704896540
transform 1 0 23552 0 1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_253
timestamp 1704896540
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_265
timestamp 1704896540
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_277
timestamp 1704896540
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_289
timestamp 1704896540
transform 1 0 27692 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_301
timestamp 1704896540
transform 1 0 28796 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_307
timestamp 1704896540
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_309
timestamp 1704896540
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_321
timestamp 1704896540
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_333
timestamp 1704896540
transform 1 0 31740 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_345
timestamp 1704896540
transform 1 0 32844 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_357
timestamp 1704896540
transform 1 0 33948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_363
timestamp 1704896540
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_365
timestamp 1704896540
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_377
timestamp 1704896540
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_389
timestamp 1704896540
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_401
timestamp 1704896540
transform 1 0 37996 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_413
timestamp 1704896540
transform 1 0 39100 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_419
timestamp 1704896540
transform 1 0 39652 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_421
timestamp 1704896540
transform 1 0 39836 0 1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_3
timestamp 1704896540
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_15
timestamp 1704896540
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_27
timestamp 1704896540
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_39
timestamp 1704896540
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_51
timestamp 1704896540
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_55
timestamp 1704896540
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_57
timestamp 1704896540
transform 1 0 6348 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_68
timestamp 1704896540
transform 1 0 7360 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_79
timestamp 1704896540
transform 1 0 8372 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_91
timestamp 1704896540
transform 1 0 9476 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_103
timestamp 1704896540
transform 1 0 10580 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_111
timestamp 1704896540
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_113
timestamp 1704896540
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_125
timestamp 1704896540
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_137
timestamp 1704896540
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_149
timestamp 1704896540
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_161
timestamp 1704896540
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_167
timestamp 1704896540
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_169
timestamp 1704896540
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_181
timestamp 1704896540
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_193
timestamp 1704896540
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_205
timestamp 1704896540
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_217
timestamp 1704896540
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_223
timestamp 1704896540
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_225
timestamp 1704896540
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_237
timestamp 1704896540
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_249
timestamp 1704896540
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_261
timestamp 1704896540
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_273
timestamp 1704896540
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_279
timestamp 1704896540
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_281
timestamp 1704896540
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_293
timestamp 1704896540
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_305
timestamp 1704896540
transform 1 0 29164 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_317
timestamp 1704896540
transform 1 0 30268 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_329
timestamp 1704896540
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_335
timestamp 1704896540
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_337
timestamp 1704896540
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_349
timestamp 1704896540
transform 1 0 33212 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_353
timestamp 1704896540
transform 1 0 33580 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_368
timestamp 1704896540
transform 1 0 34960 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_380
timestamp 1704896540
transform 1 0 36064 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_393
timestamp 1704896540
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_405
timestamp 1704896540
transform 1 0 38364 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_417
timestamp 1704896540
transform 1 0 39468 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_3
timestamp 1704896540
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_15
timestamp 1704896540
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_27
timestamp 1704896540
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_29
timestamp 1704896540
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_41
timestamp 1704896540
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_53
timestamp 1704896540
transform 1 0 5980 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_61
timestamp 1704896540
transform 1 0 6716 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_80
timestamp 1704896540
transform 1 0 8464 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_85
timestamp 1704896540
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_97
timestamp 1704896540
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_109
timestamp 1704896540
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_121
timestamp 1704896540
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_133
timestamp 1704896540
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_139
timestamp 1704896540
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_141
timestamp 1704896540
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_153
timestamp 1704896540
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_165
timestamp 1704896540
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_177
timestamp 1704896540
transform 1 0 17388 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_195
timestamp 1704896540
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_197
timestamp 1704896540
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_209
timestamp 1704896540
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_221
timestamp 1704896540
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_233
timestamp 1704896540
transform 1 0 22540 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_245
timestamp 1704896540
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_251
timestamp 1704896540
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_253
timestamp 1704896540
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_265
timestamp 1704896540
transform 1 0 25484 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_278
timestamp 1704896540
transform 1 0 26680 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_290
timestamp 1704896540
transform 1 0 27784 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_302
timestamp 1704896540
transform 1 0 28888 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_309
timestamp 1704896540
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_321
timestamp 1704896540
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_333
timestamp 1704896540
transform 1 0 31740 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_345
timestamp 1704896540
transform 1 0 32844 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_355
timestamp 1704896540
transform 1 0 33764 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_363
timestamp 1704896540
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_365
timestamp 1704896540
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_377
timestamp 1704896540
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_389
timestamp 1704896540
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_401
timestamp 1704896540
transform 1 0 37996 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_413
timestamp 1704896540
transform 1 0 39100 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_419
timestamp 1704896540
transform 1 0 39652 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_421
timestamp 1704896540
transform 1 0 39836 0 1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_3
timestamp 1704896540
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_15
timestamp 1704896540
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_27
timestamp 1704896540
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_39
timestamp 1704896540
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_51
timestamp 1704896540
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_55
timestamp 1704896540
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_57
timestamp 1704896540
transform 1 0 6348 0 -1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_72
timestamp 1704896540
transform 1 0 7728 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_84
timestamp 1704896540
transform 1 0 8832 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_96
timestamp 1704896540
transform 1 0 9936 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_113
timestamp 1704896540
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_125
timestamp 1704896540
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_137
timestamp 1704896540
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_149
timestamp 1704896540
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_161
timestamp 1704896540
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_167
timestamp 1704896540
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_169
timestamp 1704896540
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_181
timestamp 1704896540
transform 1 0 17756 0 -1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_207
timestamp 1704896540
transform 1 0 20148 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_219
timestamp 1704896540
transform 1 0 21252 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_223
timestamp 1704896540
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_225
timestamp 1704896540
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_237
timestamp 1704896540
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_249
timestamp 1704896540
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_261
timestamp 1704896540
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_273
timestamp 1704896540
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_279
timestamp 1704896540
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_281
timestamp 1704896540
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_293
timestamp 1704896540
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_305
timestamp 1704896540
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_317
timestamp 1704896540
transform 1 0 30268 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_329
timestamp 1704896540
transform 1 0 31372 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_335
timestamp 1704896540
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_337
timestamp 1704896540
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_349
timestamp 1704896540
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_361
timestamp 1704896540
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_373
timestamp 1704896540
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_385
timestamp 1704896540
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_391
timestamp 1704896540
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_393
timestamp 1704896540
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_405
timestamp 1704896540
transform 1 0 38364 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_417
timestamp 1704896540
transform 1 0 39468 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_3
timestamp 1704896540
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_15
timestamp 1704896540
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_27
timestamp 1704896540
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_29
timestamp 1704896540
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_41
timestamp 1704896540
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_53
timestamp 1704896540
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_65
timestamp 1704896540
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_77
timestamp 1704896540
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_83
timestamp 1704896540
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_85
timestamp 1704896540
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_97
timestamp 1704896540
transform 1 0 10028 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_106
timestamp 1704896540
transform 1 0 10856 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_118
timestamp 1704896540
transform 1 0 11960 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_130
timestamp 1704896540
transform 1 0 13064 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_138
timestamp 1704896540
transform 1 0 13800 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_141
timestamp 1704896540
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_153
timestamp 1704896540
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_165
timestamp 1704896540
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_177
timestamp 1704896540
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_189
timestamp 1704896540
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_195
timestamp 1704896540
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_197
timestamp 1704896540
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_209
timestamp 1704896540
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_221
timestamp 1704896540
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_233
timestamp 1704896540
transform 1 0 22540 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_245
timestamp 1704896540
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_251
timestamp 1704896540
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_253
timestamp 1704896540
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_265
timestamp 1704896540
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_277
timestamp 1704896540
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_289
timestamp 1704896540
transform 1 0 27692 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_301
timestamp 1704896540
transform 1 0 28796 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_307
timestamp 1704896540
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_309
timestamp 1704896540
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_321
timestamp 1704896540
transform 1 0 30636 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_333
timestamp 1704896540
transform 1 0 31740 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_345
timestamp 1704896540
transform 1 0 32844 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_357
timestamp 1704896540
transform 1 0 33948 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_363
timestamp 1704896540
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_365
timestamp 1704896540
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_377
timestamp 1704896540
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_389
timestamp 1704896540
transform 1 0 36892 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_395
timestamp 1704896540
transform 1 0 37444 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_408
timestamp 1704896540
transform 1 0 38640 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_421
timestamp 1704896540
transform 1 0 39836 0 1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_3
timestamp 1704896540
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_15
timestamp 1704896540
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_27
timestamp 1704896540
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_39
timestamp 1704896540
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_51
timestamp 1704896540
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_55
timestamp 1704896540
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_57
timestamp 1704896540
transform 1 0 6348 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_77
timestamp 1704896540
transform 1 0 8188 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_89
timestamp 1704896540
transform 1 0 9292 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_101
timestamp 1704896540
transform 1 0 10396 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_109
timestamp 1704896540
transform 1 0 11132 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_113
timestamp 1704896540
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_125
timestamp 1704896540
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_137
timestamp 1704896540
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_149
timestamp 1704896540
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_161
timestamp 1704896540
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_167
timestamp 1704896540
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_169
timestamp 1704896540
transform 1 0 16652 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_177
timestamp 1704896540
transform 1 0 17388 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_185
timestamp 1704896540
transform 1 0 18124 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_197
timestamp 1704896540
transform 1 0 19228 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_209
timestamp 1704896540
transform 1 0 20332 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_221
timestamp 1704896540
transform 1 0 21436 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_225
timestamp 1704896540
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_237
timestamp 1704896540
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_249
timestamp 1704896540
transform 1 0 24012 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_255
timestamp 1704896540
transform 1 0 24564 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_263
timestamp 1704896540
transform 1 0 25300 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_275
timestamp 1704896540
transform 1 0 26404 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_279
timestamp 1704896540
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_281
timestamp 1704896540
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_293
timestamp 1704896540
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_305
timestamp 1704896540
transform 1 0 29164 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_317
timestamp 1704896540
transform 1 0 30268 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_329
timestamp 1704896540
transform 1 0 31372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_335
timestamp 1704896540
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_337
timestamp 1704896540
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_349
timestamp 1704896540
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_361
timestamp 1704896540
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_373
timestamp 1704896540
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_385
timestamp 1704896540
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_391
timestamp 1704896540
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_393
timestamp 1704896540
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_405
timestamp 1704896540
transform 1 0 38364 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_417
timestamp 1704896540
transform 1 0 39468 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_3
timestamp 1704896540
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_15
timestamp 1704896540
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_27
timestamp 1704896540
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_29
timestamp 1704896540
transform 1 0 3772 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_39
timestamp 1704896540
transform 1 0 4692 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_51
timestamp 1704896540
transform 1 0 5796 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_63
timestamp 1704896540
transform 1 0 6900 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_75
timestamp 1704896540
transform 1 0 8004 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_83
timestamp 1704896540
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_85
timestamp 1704896540
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_97
timestamp 1704896540
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_109
timestamp 1704896540
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_121
timestamp 1704896540
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_133
timestamp 1704896540
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_139
timestamp 1704896540
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_141
timestamp 1704896540
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_153
timestamp 1704896540
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_165
timestamp 1704896540
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_177
timestamp 1704896540
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_189
timestamp 1704896540
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_195
timestamp 1704896540
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_197
timestamp 1704896540
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_209
timestamp 1704896540
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_221
timestamp 1704896540
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_233
timestamp 1704896540
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_245
timestamp 1704896540
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_251
timestamp 1704896540
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_253
timestamp 1704896540
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_265
timestamp 1704896540
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_277
timestamp 1704896540
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_289
timestamp 1704896540
transform 1 0 27692 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_301
timestamp 1704896540
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_307
timestamp 1704896540
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_309
timestamp 1704896540
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_321
timestamp 1704896540
transform 1 0 30636 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_325
timestamp 1704896540
transform 1 0 31004 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_329
timestamp 1704896540
transform 1 0 31372 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_339
timestamp 1704896540
transform 1 0 32292 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_343
timestamp 1704896540
transform 1 0 32660 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_355
timestamp 1704896540
transform 1 0 33764 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_363
timestamp 1704896540
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_365
timestamp 1704896540
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_377
timestamp 1704896540
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_389
timestamp 1704896540
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_401
timestamp 1704896540
transform 1 0 37996 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_413
timestamp 1704896540
transform 1 0 39100 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_419
timestamp 1704896540
transform 1 0 39652 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_421
timestamp 1704896540
transform 1 0 39836 0 1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_3
timestamp 1704896540
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_15
timestamp 1704896540
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_27
timestamp 1704896540
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_39
timestamp 1704896540
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_51
timestamp 1704896540
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_55
timestamp 1704896540
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_57
timestamp 1704896540
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_69
timestamp 1704896540
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_81
timestamp 1704896540
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_93
timestamp 1704896540
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_105
timestamp 1704896540
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_111
timestamp 1704896540
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_113
timestamp 1704896540
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_125
timestamp 1704896540
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_137
timestamp 1704896540
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_149
timestamp 1704896540
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_161
timestamp 1704896540
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_167
timestamp 1704896540
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_169
timestamp 1704896540
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_181
timestamp 1704896540
transform 1 0 17756 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_192
timestamp 1704896540
transform 1 0 18768 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_204
timestamp 1704896540
transform 1 0 19872 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_216
timestamp 1704896540
transform 1 0 20976 0 -1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_225
timestamp 1704896540
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_237
timestamp 1704896540
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_249
timestamp 1704896540
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_261
timestamp 1704896540
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_273
timestamp 1704896540
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_279
timestamp 1704896540
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_281
timestamp 1704896540
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_293
timestamp 1704896540
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_305
timestamp 1704896540
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_317
timestamp 1704896540
transform 1 0 30268 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_329
timestamp 1704896540
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_335
timestamp 1704896540
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_337
timestamp 1704896540
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_349
timestamp 1704896540
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_361
timestamp 1704896540
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_373
timestamp 1704896540
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_385
timestamp 1704896540
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_391
timestamp 1704896540
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_393
timestamp 1704896540
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_405
timestamp 1704896540
transform 1 0 38364 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_417
timestamp 1704896540
transform 1 0 39468 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_3
timestamp 1704896540
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_15
timestamp 1704896540
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_27
timestamp 1704896540
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_29
timestamp 1704896540
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_41
timestamp 1704896540
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_53
timestamp 1704896540
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_65
timestamp 1704896540
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_77
timestamp 1704896540
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_83
timestamp 1704896540
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_85
timestamp 1704896540
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_97
timestamp 1704896540
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_109
timestamp 1704896540
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_121
timestamp 1704896540
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_133
timestamp 1704896540
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_139
timestamp 1704896540
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_141
timestamp 1704896540
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_153
timestamp 1704896540
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_165
timestamp 1704896540
transform 1 0 16284 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_177
timestamp 1704896540
transform 1 0 17388 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_189
timestamp 1704896540
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_195
timestamp 1704896540
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_197
timestamp 1704896540
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_209
timestamp 1704896540
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_221
timestamp 1704896540
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_233
timestamp 1704896540
transform 1 0 22540 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_245
timestamp 1704896540
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_251
timestamp 1704896540
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_253
timestamp 1704896540
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_265
timestamp 1704896540
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_277
timestamp 1704896540
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_289
timestamp 1704896540
transform 1 0 27692 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_301
timestamp 1704896540
transform 1 0 28796 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_307
timestamp 1704896540
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_309
timestamp 1704896540
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_321
timestamp 1704896540
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_333
timestamp 1704896540
transform 1 0 31740 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_345
timestamp 1704896540
transform 1 0 32844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_357
timestamp 1704896540
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_363
timestamp 1704896540
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_379
timestamp 1704896540
transform 1 0 35972 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_391
timestamp 1704896540
transform 1 0 37076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_403
timestamp 1704896540
transform 1 0 38180 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_415
timestamp 1704896540
transform 1 0 39284 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_419
timestamp 1704896540
transform 1 0 39652 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_421
timestamp 1704896540
transform 1 0 39836 0 1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_3
timestamp 1704896540
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_15
timestamp 1704896540
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_27
timestamp 1704896540
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_39
timestamp 1704896540
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_51
timestamp 1704896540
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_55
timestamp 1704896540
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_57
timestamp 1704896540
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_69
timestamp 1704896540
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_81
timestamp 1704896540
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_93
timestamp 1704896540
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_105
timestamp 1704896540
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_111
timestamp 1704896540
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_113
timestamp 1704896540
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_125
timestamp 1704896540
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_137
timestamp 1704896540
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_149
timestamp 1704896540
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_161
timestamp 1704896540
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_167
timestamp 1704896540
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_169
timestamp 1704896540
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_181
timestamp 1704896540
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_193
timestamp 1704896540
transform 1 0 18860 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_205
timestamp 1704896540
transform 1 0 19964 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_217
timestamp 1704896540
transform 1 0 21068 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_223
timestamp 1704896540
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_225
timestamp 1704896540
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_237
timestamp 1704896540
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_249
timestamp 1704896540
transform 1 0 24012 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_262
timestamp 1704896540
transform 1 0 25208 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_274
timestamp 1704896540
transform 1 0 26312 0 -1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_281
timestamp 1704896540
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_293
timestamp 1704896540
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_305
timestamp 1704896540
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_317
timestamp 1704896540
transform 1 0 30268 0 -1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_337
timestamp 1704896540
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_349
timestamp 1704896540
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_361
timestamp 1704896540
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_373
timestamp 1704896540
transform 1 0 35420 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_385
timestamp 1704896540
transform 1 0 36524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_391
timestamp 1704896540
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_393
timestamp 1704896540
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_405
timestamp 1704896540
transform 1 0 38364 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_417
timestamp 1704896540
transform 1 0 39468 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_3
timestamp 1704896540
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_15
timestamp 1704896540
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_27
timestamp 1704896540
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_29
timestamp 1704896540
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_41
timestamp 1704896540
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_53
timestamp 1704896540
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_65
timestamp 1704896540
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_77
timestamp 1704896540
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_83
timestamp 1704896540
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_85
timestamp 1704896540
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_97
timestamp 1704896540
transform 1 0 10028 0 1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_108
timestamp 1704896540
transform 1 0 11040 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_120
timestamp 1704896540
transform 1 0 12144 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_132
timestamp 1704896540
transform 1 0 13248 0 1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_141
timestamp 1704896540
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_153
timestamp 1704896540
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_182
timestamp 1704896540
transform 1 0 17848 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_194
timestamp 1704896540
transform 1 0 18952 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_197
timestamp 1704896540
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_209
timestamp 1704896540
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_221
timestamp 1704896540
transform 1 0 21436 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_233
timestamp 1704896540
transform 1 0 22540 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_245
timestamp 1704896540
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_251
timestamp 1704896540
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_253
timestamp 1704896540
transform 1 0 24380 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_264
timestamp 1704896540
transform 1 0 25392 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_276
timestamp 1704896540
transform 1 0 26496 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_288
timestamp 1704896540
transform 1 0 27600 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_300
timestamp 1704896540
transform 1 0 28704 0 1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_309
timestamp 1704896540
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_321
timestamp 1704896540
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_333
timestamp 1704896540
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_345
timestamp 1704896540
transform 1 0 32844 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_357
timestamp 1704896540
transform 1 0 33948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_363
timestamp 1704896540
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_365
timestamp 1704896540
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_377
timestamp 1704896540
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_389
timestamp 1704896540
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_401
timestamp 1704896540
transform 1 0 37996 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_413
timestamp 1704896540
transform 1 0 39100 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_419
timestamp 1704896540
transform 1 0 39652 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_421
timestamp 1704896540
transform 1 0 39836 0 1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_3
timestamp 1704896540
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_15
timestamp 1704896540
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_27
timestamp 1704896540
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_39
timestamp 1704896540
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_51
timestamp 1704896540
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_55
timestamp 1704896540
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_57
timestamp 1704896540
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_69
timestamp 1704896540
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_81
timestamp 1704896540
transform 1 0 8556 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_85
timestamp 1704896540
transform 1 0 8924 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_94
timestamp 1704896540
transform 1 0 9752 0 -1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_125
timestamp 1704896540
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_137
timestamp 1704896540
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_149
timestamp 1704896540
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_161
timestamp 1704896540
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_167
timestamp 1704896540
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_169
timestamp 1704896540
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_181
timestamp 1704896540
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_193
timestamp 1704896540
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_205
timestamp 1704896540
transform 1 0 19964 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_217
timestamp 1704896540
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_223
timestamp 1704896540
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_225
timestamp 1704896540
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_237
timestamp 1704896540
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_249
timestamp 1704896540
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_261
timestamp 1704896540
transform 1 0 25116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_273
timestamp 1704896540
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_279
timestamp 1704896540
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_281
timestamp 1704896540
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_293
timestamp 1704896540
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_305
timestamp 1704896540
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_317
timestamp 1704896540
transform 1 0 30268 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_329
timestamp 1704896540
transform 1 0 31372 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_335
timestamp 1704896540
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_337
timestamp 1704896540
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_349
timestamp 1704896540
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_361
timestamp 1704896540
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_373
timestamp 1704896540
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_385
timestamp 1704896540
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_391
timestamp 1704896540
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_393
timestamp 1704896540
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_405
timestamp 1704896540
transform 1 0 38364 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_415
timestamp 1704896540
transform 1 0 39284 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_427
timestamp 1704896540
transform 1 0 40388 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_3
timestamp 1704896540
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_15
timestamp 1704896540
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_27
timestamp 1704896540
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_29
timestamp 1704896540
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_41
timestamp 1704896540
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_53
timestamp 1704896540
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_65
timestamp 1704896540
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_77
timestamp 1704896540
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_83
timestamp 1704896540
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_85
timestamp 1704896540
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_97
timestamp 1704896540
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_109
timestamp 1704896540
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_121
timestamp 1704896540
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_133
timestamp 1704896540
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_139
timestamp 1704896540
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_141
timestamp 1704896540
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_153
timestamp 1704896540
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_165
timestamp 1704896540
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_177
timestamp 1704896540
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_189
timestamp 1704896540
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_195
timestamp 1704896540
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_197
timestamp 1704896540
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_216
timestamp 1704896540
transform 1 0 20976 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_222
timestamp 1704896540
transform 1 0 21528 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_231
timestamp 1704896540
transform 1 0 22356 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_243
timestamp 1704896540
transform 1 0 23460 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_251
timestamp 1704896540
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_253
timestamp 1704896540
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_265
timestamp 1704896540
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_277
timestamp 1704896540
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_289
timestamp 1704896540
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_301
timestamp 1704896540
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_307
timestamp 1704896540
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_309
timestamp 1704896540
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_321
timestamp 1704896540
transform 1 0 30636 0 1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_343
timestamp 1704896540
transform 1 0 32660 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_355
timestamp 1704896540
transform 1 0 33764 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_363
timestamp 1704896540
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_365
timestamp 1704896540
transform 1 0 34684 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_373
timestamp 1704896540
transform 1 0 35420 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_377
timestamp 1704896540
transform 1 0 35788 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_386
timestamp 1704896540
transform 1 0 36616 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_390
timestamp 1704896540
transform 1 0 36984 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_402
timestamp 1704896540
transform 1 0 38088 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_414
timestamp 1704896540
transform 1 0 39192 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_421
timestamp 1704896540
transform 1 0 39836 0 1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_3
timestamp 1704896540
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_15
timestamp 1704896540
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_27
timestamp 1704896540
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_39
timestamp 1704896540
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_51
timestamp 1704896540
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_55
timestamp 1704896540
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_57
timestamp 1704896540
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_69
timestamp 1704896540
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_81
timestamp 1704896540
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_93
timestamp 1704896540
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_105
timestamp 1704896540
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_111
timestamp 1704896540
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_113
timestamp 1704896540
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_125
timestamp 1704896540
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_137
timestamp 1704896540
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_149
timestamp 1704896540
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_161
timestamp 1704896540
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_167
timestamp 1704896540
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_169
timestamp 1704896540
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_181
timestamp 1704896540
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_193
timestamp 1704896540
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_205
timestamp 1704896540
transform 1 0 19964 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_217
timestamp 1704896540
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_223
timestamp 1704896540
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_225
timestamp 1704896540
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_237
timestamp 1704896540
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_249
timestamp 1704896540
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_261
timestamp 1704896540
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_273
timestamp 1704896540
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_279
timestamp 1704896540
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_281
timestamp 1704896540
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_293
timestamp 1704896540
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_305
timestamp 1704896540
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_330
timestamp 1704896540
transform 1 0 31464 0 -1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_337
timestamp 1704896540
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_349
timestamp 1704896540
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_361
timestamp 1704896540
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_373
timestamp 1704896540
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_385
timestamp 1704896540
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_391
timestamp 1704896540
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_393
timestamp 1704896540
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_405
timestamp 1704896540
transform 1 0 38364 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_417
timestamp 1704896540
transform 1 0 39468 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_3
timestamp 1704896540
transform 1 0 1380 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_7
timestamp 1704896540
transform 1 0 1748 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_15
timestamp 1704896540
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_27
timestamp 1704896540
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_29
timestamp 1704896540
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_41
timestamp 1704896540
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_53
timestamp 1704896540
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_65
timestamp 1704896540
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_77
timestamp 1704896540
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_83
timestamp 1704896540
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_85
timestamp 1704896540
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_97
timestamp 1704896540
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_109
timestamp 1704896540
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_121
timestamp 1704896540
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_133
timestamp 1704896540
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_139
timestamp 1704896540
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_141
timestamp 1704896540
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_153
timestamp 1704896540
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_165
timestamp 1704896540
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_177
timestamp 1704896540
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_189
timestamp 1704896540
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_195
timestamp 1704896540
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_197
timestamp 1704896540
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_209
timestamp 1704896540
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_221
timestamp 1704896540
transform 1 0 21436 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_233
timestamp 1704896540
transform 1 0 22540 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_245
timestamp 1704896540
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_251
timestamp 1704896540
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_253
timestamp 1704896540
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_265
timestamp 1704896540
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_277
timestamp 1704896540
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_289
timestamp 1704896540
transform 1 0 27692 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_301
timestamp 1704896540
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_307
timestamp 1704896540
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_309
timestamp 1704896540
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_321
timestamp 1704896540
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_333
timestamp 1704896540
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_345
timestamp 1704896540
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_357
timestamp 1704896540
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_363
timestamp 1704896540
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_365
timestamp 1704896540
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_377
timestamp 1704896540
transform 1 0 35788 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_390
timestamp 1704896540
transform 1 0 36984 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_402
timestamp 1704896540
transform 1 0 38088 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_414
timestamp 1704896540
transform 1 0 39192 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_421
timestamp 1704896540
transform 1 0 39836 0 1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_3
timestamp 1704896540
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_15
timestamp 1704896540
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_27
timestamp 1704896540
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_39
timestamp 1704896540
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_51
timestamp 1704896540
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_55
timestamp 1704896540
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_57
timestamp 1704896540
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_69
timestamp 1704896540
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_81
timestamp 1704896540
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_93
timestamp 1704896540
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_105
timestamp 1704896540
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_111
timestamp 1704896540
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_113
timestamp 1704896540
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_125
timestamp 1704896540
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_137
timestamp 1704896540
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_149
timestamp 1704896540
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_161
timestamp 1704896540
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_167
timestamp 1704896540
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_174
timestamp 1704896540
transform 1 0 17112 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_186
timestamp 1704896540
transform 1 0 18216 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_198
timestamp 1704896540
transform 1 0 19320 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_210
timestamp 1704896540
transform 1 0 20424 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_222
timestamp 1704896540
transform 1 0 21528 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_225
timestamp 1704896540
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_237
timestamp 1704896540
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_249
timestamp 1704896540
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_261
timestamp 1704896540
transform 1 0 25116 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_273
timestamp 1704896540
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_279
timestamp 1704896540
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_281
timestamp 1704896540
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_293
timestamp 1704896540
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_305
timestamp 1704896540
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_317
timestamp 1704896540
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_329
timestamp 1704896540
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_335
timestamp 1704896540
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_337
timestamp 1704896540
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_349
timestamp 1704896540
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_361
timestamp 1704896540
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_373
timestamp 1704896540
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_385
timestamp 1704896540
transform 1 0 36524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_391
timestamp 1704896540
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_393
timestamp 1704896540
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_405
timestamp 1704896540
transform 1 0 38364 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_9
timestamp 1704896540
transform 1 0 1932 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_21
timestamp 1704896540
transform 1 0 3036 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_27
timestamp 1704896540
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_29
timestamp 1704896540
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_41
timestamp 1704896540
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_53
timestamp 1704896540
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_65
timestamp 1704896540
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_77
timestamp 1704896540
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_83
timestamp 1704896540
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_85
timestamp 1704896540
transform 1 0 8924 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_102
timestamp 1704896540
transform 1 0 10488 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_114
timestamp 1704896540
transform 1 0 11592 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_126
timestamp 1704896540
transform 1 0 12696 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_138
timestamp 1704896540
transform 1 0 13800 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_141
timestamp 1704896540
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_153
timestamp 1704896540
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_165
timestamp 1704896540
transform 1 0 16284 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_178
timestamp 1704896540
transform 1 0 17480 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_186
timestamp 1704896540
transform 1 0 18216 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_195
timestamp 1704896540
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_197
timestamp 1704896540
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_209
timestamp 1704896540
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_221
timestamp 1704896540
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_233
timestamp 1704896540
transform 1 0 22540 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_245
timestamp 1704896540
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_251
timestamp 1704896540
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_253
timestamp 1704896540
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_265
timestamp 1704896540
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_277
timestamp 1704896540
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_289
timestamp 1704896540
transform 1 0 27692 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_301
timestamp 1704896540
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_307
timestamp 1704896540
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_309
timestamp 1704896540
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_321
timestamp 1704896540
transform 1 0 30636 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_329
timestamp 1704896540
transform 1 0 31372 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_341
timestamp 1704896540
transform 1 0 32476 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_353
timestamp 1704896540
transform 1 0 33580 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_361
timestamp 1704896540
transform 1 0 34316 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_365
timestamp 1704896540
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_377
timestamp 1704896540
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_389
timestamp 1704896540
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_401
timestamp 1704896540
transform 1 0 37996 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_413
timestamp 1704896540
transform 1 0 39100 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_419
timestamp 1704896540
transform 1 0 39652 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_421
timestamp 1704896540
transform 1 0 39836 0 1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_3
timestamp 1704896540
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_15
timestamp 1704896540
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_27
timestamp 1704896540
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_39
timestamp 1704896540
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_51
timestamp 1704896540
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_55
timestamp 1704896540
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_64
timestamp 1704896540
transform 1 0 6992 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_76
timestamp 1704896540
transform 1 0 8096 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_88
timestamp 1704896540
transform 1 0 9200 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_100
timestamp 1704896540
transform 1 0 10304 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_113
timestamp 1704896540
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_125
timestamp 1704896540
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_137
timestamp 1704896540
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_149
timestamp 1704896540
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_161
timestamp 1704896540
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_167
timestamp 1704896540
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_169
timestamp 1704896540
transform 1 0 16652 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_176
timestamp 1704896540
transform 1 0 17296 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_188
timestamp 1704896540
transform 1 0 18400 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_200
timestamp 1704896540
transform 1 0 19504 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_208
timestamp 1704896540
transform 1 0 20240 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_220
timestamp 1704896540
transform 1 0 21344 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_225
timestamp 1704896540
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_237
timestamp 1704896540
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_249
timestamp 1704896540
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_261
timestamp 1704896540
transform 1 0 25116 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_273
timestamp 1704896540
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_279
timestamp 1704896540
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_281
timestamp 1704896540
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_293
timestamp 1704896540
transform 1 0 28060 0 -1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_307
timestamp 1704896540
transform 1 0 29348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_319
timestamp 1704896540
transform 1 0 30452 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_331
timestamp 1704896540
transform 1 0 31556 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_335
timestamp 1704896540
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_337
timestamp 1704896540
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_349
timestamp 1704896540
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_361
timestamp 1704896540
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_373
timestamp 1704896540
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_385
timestamp 1704896540
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_391
timestamp 1704896540
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_393
timestamp 1704896540
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_405
timestamp 1704896540
transform 1 0 38364 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_417
timestamp 1704896540
transform 1 0 39468 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_3
timestamp 1704896540
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_15
timestamp 1704896540
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_27
timestamp 1704896540
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_29
timestamp 1704896540
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_41
timestamp 1704896540
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_53
timestamp 1704896540
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_65
timestamp 1704896540
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_77
timestamp 1704896540
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_83
timestamp 1704896540
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_85
timestamp 1704896540
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_97
timestamp 1704896540
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_109
timestamp 1704896540
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_121
timestamp 1704896540
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_133
timestamp 1704896540
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_139
timestamp 1704896540
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_141
timestamp 1704896540
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_153
timestamp 1704896540
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_56_165
timestamp 1704896540
transform 1 0 16284 0 1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_172
timestamp 1704896540
transform 1 0 16928 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_184
timestamp 1704896540
transform 1 0 18032 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_197
timestamp 1704896540
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_209
timestamp 1704896540
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_221
timestamp 1704896540
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_233
timestamp 1704896540
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_245
timestamp 1704896540
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_251
timestamp 1704896540
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_253
timestamp 1704896540
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_265
timestamp 1704896540
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_277
timestamp 1704896540
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_289
timestamp 1704896540
transform 1 0 27692 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_301
timestamp 1704896540
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_307
timestamp 1704896540
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_309
timestamp 1704896540
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_321
timestamp 1704896540
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_333
timestamp 1704896540
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_345
timestamp 1704896540
transform 1 0 32844 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_359
timestamp 1704896540
transform 1 0 34132 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_363
timestamp 1704896540
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_365
timestamp 1704896540
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_377
timestamp 1704896540
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_389
timestamp 1704896540
transform 1 0 36892 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_416
timestamp 1704896540
transform 1 0 39376 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_421
timestamp 1704896540
transform 1 0 39836 0 1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_3
timestamp 1704896540
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_15
timestamp 1704896540
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_27
timestamp 1704896540
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_39
timestamp 1704896540
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_51
timestamp 1704896540
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_55
timestamp 1704896540
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_62
timestamp 1704896540
transform 1 0 6808 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_74
timestamp 1704896540
transform 1 0 7912 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_86
timestamp 1704896540
transform 1 0 9016 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_98
timestamp 1704896540
transform 1 0 10120 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_110
timestamp 1704896540
transform 1 0 11224 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_113
timestamp 1704896540
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_125
timestamp 1704896540
transform 1 0 12604 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57_133
timestamp 1704896540
transform 1 0 13340 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_153
timestamp 1704896540
transform 1 0 15180 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57_165
timestamp 1704896540
transform 1 0 16284 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_169
timestamp 1704896540
transform 1 0 16652 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57_177
timestamp 1704896540
transform 1 0 17388 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_183
timestamp 1704896540
transform 1 0 17940 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_187
timestamp 1704896540
transform 1 0 18308 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_193
timestamp 1704896540
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_205
timestamp 1704896540
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_217
timestamp 1704896540
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_223
timestamp 1704896540
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_225
timestamp 1704896540
transform 1 0 21804 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_249
timestamp 1704896540
transform 1 0 24012 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_257
timestamp 1704896540
transform 1 0 24748 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_281
timestamp 1704896540
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_293
timestamp 1704896540
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_305
timestamp 1704896540
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_317
timestamp 1704896540
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_329
timestamp 1704896540
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_335
timestamp 1704896540
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_337
timestamp 1704896540
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_349
timestamp 1704896540
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_361
timestamp 1704896540
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_373
timestamp 1704896540
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_385
timestamp 1704896540
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_391
timestamp 1704896540
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_393
timestamp 1704896540
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_405
timestamp 1704896540
transform 1 0 38364 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_417
timestamp 1704896540
transform 1 0 39468 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_3
timestamp 1704896540
transform 1 0 1380 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_16
timestamp 1704896540
transform 1 0 2576 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_29
timestamp 1704896540
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_41
timestamp 1704896540
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_53
timestamp 1704896540
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_65
timestamp 1704896540
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_77
timestamp 1704896540
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_83
timestamp 1704896540
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_85
timestamp 1704896540
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_97
timestamp 1704896540
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_109
timestamp 1704896540
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_121
timestamp 1704896540
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_133
timestamp 1704896540
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_139
timestamp 1704896540
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_141
timestamp 1704896540
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_153
timestamp 1704896540
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_165
timestamp 1704896540
transform 1 0 16284 0 1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_177
timestamp 1704896540
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_189
timestamp 1704896540
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_195
timestamp 1704896540
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_197
timestamp 1704896540
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_209
timestamp 1704896540
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_221
timestamp 1704896540
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_233
timestamp 1704896540
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_245
timestamp 1704896540
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_251
timestamp 1704896540
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_253
timestamp 1704896540
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_265
timestamp 1704896540
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_277
timestamp 1704896540
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_289
timestamp 1704896540
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_301
timestamp 1704896540
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_307
timestamp 1704896540
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_309
timestamp 1704896540
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_321
timestamp 1704896540
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_333
timestamp 1704896540
transform 1 0 31740 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_341
timestamp 1704896540
transform 1 0 32476 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_353
timestamp 1704896540
transform 1 0 33580 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_58_361
timestamp 1704896540
transform 1 0 34316 0 1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_365
timestamp 1704896540
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_377
timestamp 1704896540
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_389
timestamp 1704896540
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_401
timestamp 1704896540
transform 1 0 37996 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_413
timestamp 1704896540
transform 1 0 39100 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_419
timestamp 1704896540
transform 1 0 39652 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_421
timestamp 1704896540
transform 1 0 39836 0 1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_3
timestamp 1704896540
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_15
timestamp 1704896540
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_27
timestamp 1704896540
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_39
timestamp 1704896540
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_51
timestamp 1704896540
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_55
timestamp 1704896540
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_57
timestamp 1704896540
transform 1 0 6348 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_63
timestamp 1704896540
transform 1 0 6900 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_71
timestamp 1704896540
transform 1 0 7636 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_83
timestamp 1704896540
transform 1 0 8740 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_95
timestamp 1704896540
transform 1 0 9844 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_107
timestamp 1704896540
transform 1 0 10948 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_111
timestamp 1704896540
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_113
timestamp 1704896540
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_125
timestamp 1704896540
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_137
timestamp 1704896540
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_149
timestamp 1704896540
transform 1 0 14812 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_162
timestamp 1704896540
transform 1 0 16008 0 -1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_169
timestamp 1704896540
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_181
timestamp 1704896540
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_193
timestamp 1704896540
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_205
timestamp 1704896540
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_217
timestamp 1704896540
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_223
timestamp 1704896540
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_241
timestamp 1704896540
transform 1 0 23276 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_253
timestamp 1704896540
transform 1 0 24380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_265
timestamp 1704896540
transform 1 0 25484 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59_277
timestamp 1704896540
transform 1 0 26588 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_281
timestamp 1704896540
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_293
timestamp 1704896540
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_305
timestamp 1704896540
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_317
timestamp 1704896540
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_329
timestamp 1704896540
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_335
timestamp 1704896540
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_337
timestamp 1704896540
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_349
timestamp 1704896540
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_361
timestamp 1704896540
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_373
timestamp 1704896540
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_385
timestamp 1704896540
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_391
timestamp 1704896540
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_393
timestamp 1704896540
transform 1 0 37260 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_401
timestamp 1704896540
transform 1 0 37996 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_409
timestamp 1704896540
transform 1 0 38732 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_421
timestamp 1704896540
transform 1 0 39836 0 -1 34816
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_3
timestamp 1704896540
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_15
timestamp 1704896540
transform 1 0 2484 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_27
timestamp 1704896540
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_35
timestamp 1704896540
transform 1 0 4324 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_47
timestamp 1704896540
transform 1 0 5428 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_59
timestamp 1704896540
transform 1 0 6532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_71
timestamp 1704896540
transform 1 0 7636 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_83
timestamp 1704896540
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_85
timestamp 1704896540
transform 1 0 8924 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_93
timestamp 1704896540
transform 1 0 9660 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_102
timestamp 1704896540
transform 1 0 10488 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_114
timestamp 1704896540
transform 1 0 11592 0 1 34816
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_141
timestamp 1704896540
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_153
timestamp 1704896540
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_174
timestamp 1704896540
transform 1 0 17112 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_186
timestamp 1704896540
transform 1 0 18216 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_194
timestamp 1704896540
transform 1 0 18952 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_197
timestamp 1704896540
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_209
timestamp 1704896540
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_221
timestamp 1704896540
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_233
timestamp 1704896540
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_245
timestamp 1704896540
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_251
timestamp 1704896540
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_253
timestamp 1704896540
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_265
timestamp 1704896540
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_284
timestamp 1704896540
transform 1 0 27232 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_296
timestamp 1704896540
transform 1 0 28336 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_309
timestamp 1704896540
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_321
timestamp 1704896540
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_333
timestamp 1704896540
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_345
timestamp 1704896540
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_357
timestamp 1704896540
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_363
timestamp 1704896540
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_365
timestamp 1704896540
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_377
timestamp 1704896540
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_389
timestamp 1704896540
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_401
timestamp 1704896540
transform 1 0 37996 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_413
timestamp 1704896540
transform 1 0 39100 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_419
timestamp 1704896540
transform 1 0 39652 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_421
timestamp 1704896540
transform 1 0 39836 0 1 34816
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_3
timestamp 1704896540
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_15
timestamp 1704896540
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_61_27
timestamp 1704896540
transform 1 0 3588 0 -1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_37
timestamp 1704896540
transform 1 0 4508 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_49
timestamp 1704896540
transform 1 0 5612 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_55
timestamp 1704896540
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_57
timestamp 1704896540
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_69
timestamp 1704896540
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_81
timestamp 1704896540
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_93
timestamp 1704896540
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_105
timestamp 1704896540
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_111
timestamp 1704896540
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_113
timestamp 1704896540
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_125
timestamp 1704896540
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_137
timestamp 1704896540
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_149
timestamp 1704896540
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_161
timestamp 1704896540
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_167
timestamp 1704896540
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_169
timestamp 1704896540
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_181
timestamp 1704896540
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_193
timestamp 1704896540
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_205
timestamp 1704896540
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_217
timestamp 1704896540
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_223
timestamp 1704896540
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_225
timestamp 1704896540
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_237
timestamp 1704896540
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_249
timestamp 1704896540
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_261
timestamp 1704896540
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_273
timestamp 1704896540
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_279
timestamp 1704896540
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_281
timestamp 1704896540
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_293
timestamp 1704896540
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_305
timestamp 1704896540
transform 1 0 29164 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_321
timestamp 1704896540
transform 1 0 30636 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_61_333
timestamp 1704896540
transform 1 0 31740 0 -1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_337
timestamp 1704896540
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_349
timestamp 1704896540
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_361
timestamp 1704896540
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_373
timestamp 1704896540
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_385
timestamp 1704896540
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_391
timestamp 1704896540
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_393
timestamp 1704896540
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_405
timestamp 1704896540
transform 1 0 38364 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_417
timestamp 1704896540
transform 1 0 39468 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_3
timestamp 1704896540
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_15
timestamp 1704896540
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_27
timestamp 1704896540
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_29
timestamp 1704896540
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_41
timestamp 1704896540
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_53
timestamp 1704896540
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_65
timestamp 1704896540
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_77
timestamp 1704896540
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_83
timestamp 1704896540
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62_85
timestamp 1704896540
transform 1 0 8924 0 1 35904
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_96
timestamp 1704896540
transform 1 0 9936 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_108
timestamp 1704896540
transform 1 0 11040 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_120
timestamp 1704896540
transform 1 0 12144 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62_132
timestamp 1704896540
transform 1 0 13248 0 1 35904
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_141
timestamp 1704896540
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_153
timestamp 1704896540
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_165
timestamp 1704896540
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_177
timestamp 1704896540
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_189
timestamp 1704896540
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_195
timestamp 1704896540
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_197
timestamp 1704896540
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_209
timestamp 1704896540
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_221
timestamp 1704896540
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_233
timestamp 1704896540
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_245
timestamp 1704896540
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_251
timestamp 1704896540
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_253
timestamp 1704896540
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_265
timestamp 1704896540
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_277
timestamp 1704896540
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_289
timestamp 1704896540
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_301
timestamp 1704896540
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_307
timestamp 1704896540
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_309
timestamp 1704896540
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_321
timestamp 1704896540
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_333
timestamp 1704896540
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_345
timestamp 1704896540
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_357
timestamp 1704896540
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_363
timestamp 1704896540
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_377
timestamp 1704896540
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_389
timestamp 1704896540
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_401
timestamp 1704896540
transform 1 0 37996 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_413
timestamp 1704896540
transform 1 0 39100 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_419
timestamp 1704896540
transform 1 0 39652 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62_421
timestamp 1704896540
transform 1 0 39836 0 1 35904
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_3
timestamp 1704896540
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_15
timestamp 1704896540
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_27
timestamp 1704896540
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_39
timestamp 1704896540
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_51
timestamp 1704896540
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_55
timestamp 1704896540
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_57
timestamp 1704896540
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_69
timestamp 1704896540
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_81
timestamp 1704896540
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_93
timestamp 1704896540
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_105
timestamp 1704896540
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_111
timestamp 1704896540
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_113
timestamp 1704896540
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_125
timestamp 1704896540
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_137
timestamp 1704896540
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_149
timestamp 1704896540
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_161
timestamp 1704896540
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_167
timestamp 1704896540
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_169
timestamp 1704896540
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_181
timestamp 1704896540
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_193
timestamp 1704896540
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_205
timestamp 1704896540
transform 1 0 19964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_217
timestamp 1704896540
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_223
timestamp 1704896540
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_225
timestamp 1704896540
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_237
timestamp 1704896540
transform 1 0 22908 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_260
timestamp 1704896540
transform 1 0 25024 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63_272
timestamp 1704896540
transform 1 0 26128 0 -1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_281
timestamp 1704896540
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_293
timestamp 1704896540
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_305
timestamp 1704896540
transform 1 0 29164 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_317
timestamp 1704896540
transform 1 0 30268 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_329
timestamp 1704896540
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_335
timestamp 1704896540
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_337
timestamp 1704896540
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_349
timestamp 1704896540
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_361
timestamp 1704896540
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_373
timestamp 1704896540
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_385
timestamp 1704896540
transform 1 0 36524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_391
timestamp 1704896540
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_393
timestamp 1704896540
transform 1 0 37260 0 -1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_404
timestamp 1704896540
transform 1 0 38272 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_416
timestamp 1704896540
transform 1 0 39376 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_428
timestamp 1704896540
transform 1 0 40480 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_3
timestamp 1704896540
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_15
timestamp 1704896540
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_27
timestamp 1704896540
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_29
timestamp 1704896540
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_41
timestamp 1704896540
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_53
timestamp 1704896540
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_65
timestamp 1704896540
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_77
timestamp 1704896540
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_83
timestamp 1704896540
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_85
timestamp 1704896540
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_97
timestamp 1704896540
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_109
timestamp 1704896540
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_121
timestamp 1704896540
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_133
timestamp 1704896540
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_139
timestamp 1704896540
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_141
timestamp 1704896540
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_153
timestamp 1704896540
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_165
timestamp 1704896540
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64_177
timestamp 1704896540
transform 1 0 17388 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64_181
timestamp 1704896540
transform 1 0 17756 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_190
timestamp 1704896540
transform 1 0 18584 0 1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_197
timestamp 1704896540
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_209
timestamp 1704896540
transform 1 0 20332 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_221
timestamp 1704896540
transform 1 0 21436 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_233
timestamp 1704896540
transform 1 0 22540 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_245
timestamp 1704896540
transform 1 0 23644 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_251
timestamp 1704896540
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_253
timestamp 1704896540
transform 1 0 24380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_265
timestamp 1704896540
transform 1 0 25484 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_277
timestamp 1704896540
transform 1 0 26588 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_289
timestamp 1704896540
transform 1 0 27692 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_301
timestamp 1704896540
transform 1 0 28796 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_307
timestamp 1704896540
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_309
timestamp 1704896540
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_321
timestamp 1704896540
transform 1 0 30636 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_333
timestamp 1704896540
transform 1 0 31740 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_345
timestamp 1704896540
transform 1 0 32844 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_357
timestamp 1704896540
transform 1 0 33948 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_363
timestamp 1704896540
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_365
timestamp 1704896540
transform 1 0 34684 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_369
timestamp 1704896540
transform 1 0 35052 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_377
timestamp 1704896540
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_389
timestamp 1704896540
transform 1 0 36892 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_401
timestamp 1704896540
transform 1 0 37996 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_407
timestamp 1704896540
transform 1 0 38548 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_421
timestamp 1704896540
transform 1 0 39836 0 1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_3
timestamp 1704896540
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_15
timestamp 1704896540
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_27
timestamp 1704896540
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_39
timestamp 1704896540
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65_51
timestamp 1704896540
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_55
timestamp 1704896540
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_57
timestamp 1704896540
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_69
timestamp 1704896540
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_81
timestamp 1704896540
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_93
timestamp 1704896540
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_105
timestamp 1704896540
transform 1 0 10764 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_111
timestamp 1704896540
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_113
timestamp 1704896540
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_65_125
timestamp 1704896540
transform 1 0 12604 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_147
timestamp 1704896540
transform 1 0 14628 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_65_159
timestamp 1704896540
transform 1 0 15732 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_167
timestamp 1704896540
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_169
timestamp 1704896540
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_181
timestamp 1704896540
transform 1 0 17756 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_193
timestamp 1704896540
transform 1 0 18860 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_205
timestamp 1704896540
transform 1 0 19964 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_217
timestamp 1704896540
transform 1 0 21068 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_223
timestamp 1704896540
transform 1 0 21620 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_225
timestamp 1704896540
transform 1 0 21804 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_237
timestamp 1704896540
transform 1 0 22908 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_249
timestamp 1704896540
transform 1 0 24012 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_261
timestamp 1704896540
transform 1 0 25116 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_65_271
timestamp 1704896540
transform 1 0 26036 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_279
timestamp 1704896540
transform 1 0 26772 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_286
timestamp 1704896540
transform 1 0 27416 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_298
timestamp 1704896540
transform 1 0 28520 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_310
timestamp 1704896540
transform 1 0 29624 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_322
timestamp 1704896540
transform 1 0 30728 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_65_334
timestamp 1704896540
transform 1 0 31832 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_337
timestamp 1704896540
transform 1 0 32108 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_349
timestamp 1704896540
transform 1 0 33212 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_361
timestamp 1704896540
transform 1 0 34316 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_373
timestamp 1704896540
transform 1 0 35420 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_385
timestamp 1704896540
transform 1 0 36524 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_391
timestamp 1704896540
transform 1 0 37076 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_401
timestamp 1704896540
transform 1 0 37996 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_413
timestamp 1704896540
transform 1 0 39100 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65_425
timestamp 1704896540
transform 1 0 40204 0 -1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_3
timestamp 1704896540
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_15
timestamp 1704896540
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_27
timestamp 1704896540
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_29
timestamp 1704896540
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_41
timestamp 1704896540
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_53
timestamp 1704896540
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_65
timestamp 1704896540
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_77
timestamp 1704896540
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_83
timestamp 1704896540
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_85
timestamp 1704896540
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_97
timestamp 1704896540
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_109
timestamp 1704896540
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_121
timestamp 1704896540
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_133
timestamp 1704896540
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_139
timestamp 1704896540
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_141
timestamp 1704896540
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_153
timestamp 1704896540
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_165
timestamp 1704896540
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_177
timestamp 1704896540
transform 1 0 17388 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_189
timestamp 1704896540
transform 1 0 18492 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_195
timestamp 1704896540
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_197
timestamp 1704896540
transform 1 0 19228 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_204
timestamp 1704896540
transform 1 0 19872 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_216
timestamp 1704896540
transform 1 0 20976 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_228
timestamp 1704896540
transform 1 0 22080 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_240
timestamp 1704896540
transform 1 0 23184 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_262
timestamp 1704896540
transform 1 0 25208 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_274
timestamp 1704896540
transform 1 0 26312 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_286
timestamp 1704896540
transform 1 0 27416 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_66_298
timestamp 1704896540
transform 1 0 28520 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_66_306
timestamp 1704896540
transform 1 0 29256 0 1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_309
timestamp 1704896540
transform 1 0 29532 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_321
timestamp 1704896540
transform 1 0 30636 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_333
timestamp 1704896540
transform 1 0 31740 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_345
timestamp 1704896540
transform 1 0 32844 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_357
timestamp 1704896540
transform 1 0 33948 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_363
timestamp 1704896540
transform 1 0 34500 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_365
timestamp 1704896540
transform 1 0 34684 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_377
timestamp 1704896540
transform 1 0 35788 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_389
timestamp 1704896540
transform 1 0 36892 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_401
timestamp 1704896540
transform 1 0 37996 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_413
timestamp 1704896540
transform 1 0 39100 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_419
timestamp 1704896540
transform 1 0 39652 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_66_421
timestamp 1704896540
transform 1 0 39836 0 1 38080
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_3
timestamp 1704896540
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_15
timestamp 1704896540
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_27
timestamp 1704896540
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_39
timestamp 1704896540
transform 1 0 4692 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67_51
timestamp 1704896540
transform 1 0 5796 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_55
timestamp 1704896540
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_57
timestamp 1704896540
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_69
timestamp 1704896540
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_81
timestamp 1704896540
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_93
timestamp 1704896540
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_105
timestamp 1704896540
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_111
timestamp 1704896540
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_113
timestamp 1704896540
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_125
timestamp 1704896540
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_137
timestamp 1704896540
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_149
timestamp 1704896540
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_161
timestamp 1704896540
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_167
timestamp 1704896540
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_169
timestamp 1704896540
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_181
timestamp 1704896540
transform 1 0 17756 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_193
timestamp 1704896540
transform 1 0 18860 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_67_205
timestamp 1704896540
transform 1 0 19964 0 -1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_225
timestamp 1704896540
transform 1 0 21804 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67_237
timestamp 1704896540
transform 1 0 22908 0 -1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_248
timestamp 1704896540
transform 1 0 23920 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_260
timestamp 1704896540
transform 1 0 25024 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_67_272
timestamp 1704896540
transform 1 0 26128 0 -1 39168
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_281
timestamp 1704896540
transform 1 0 26956 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_67_293
timestamp 1704896540
transform 1 0 28060 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_67_301
timestamp 1704896540
transform 1 0 28796 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_67_325
timestamp 1704896540
transform 1 0 31004 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_67_333
timestamp 1704896540
transform 1 0 31740 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_67_342
timestamp 1704896540
transform 1 0 32568 0 -1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_346
timestamp 1704896540
transform 1 0 32936 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_358
timestamp 1704896540
transform 1 0 34040 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_370
timestamp 1704896540
transform 1 0 35144 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_67_382
timestamp 1704896540
transform 1 0 36248 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_67_390
timestamp 1704896540
transform 1 0 36984 0 -1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_393
timestamp 1704896540
transform 1 0 37260 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_405
timestamp 1704896540
transform 1 0 38364 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_417
timestamp 1704896540
transform 1 0 39468 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_3
timestamp 1704896540
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_15
timestamp 1704896540
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_27
timestamp 1704896540
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_29
timestamp 1704896540
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_41
timestamp 1704896540
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_53
timestamp 1704896540
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_65
timestamp 1704896540
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_77
timestamp 1704896540
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_83
timestamp 1704896540
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_85
timestamp 1704896540
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_97
timestamp 1704896540
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_109
timestamp 1704896540
transform 1 0 11132 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_68_121
timestamp 1704896540
transform 1 0 12236 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_125
timestamp 1704896540
transform 1 0 12604 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_134
timestamp 1704896540
transform 1 0 13432 0 1 39168
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_141
timestamp 1704896540
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_153
timestamp 1704896540
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_165
timestamp 1704896540
transform 1 0 16284 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_177
timestamp 1704896540
transform 1 0 17388 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_189
timestamp 1704896540
transform 1 0 18492 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_195
timestamp 1704896540
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_197
timestamp 1704896540
transform 1 0 19228 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_209
timestamp 1704896540
transform 1 0 20332 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_221
timestamp 1704896540
transform 1 0 21436 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_68_233
timestamp 1704896540
transform 1 0 22540 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_246
timestamp 1704896540
transform 1 0 23736 0 1 39168
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_253
timestamp 1704896540
transform 1 0 24380 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_265
timestamp 1704896540
transform 1 0 25484 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_273
timestamp 1704896540
transform 1 0 26220 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_285
timestamp 1704896540
transform 1 0 27324 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_68_297
timestamp 1704896540
transform 1 0 28428 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_68_303
timestamp 1704896540
transform 1 0 28980 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_307
timestamp 1704896540
transform 1 0 29348 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_68_309
timestamp 1704896540
transform 1 0 29532 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_313
timestamp 1704896540
transform 1 0 29900 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_330
timestamp 1704896540
transform 1 0 31464 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_349
timestamp 1704896540
transform 1 0 33212 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_68_361
timestamp 1704896540
transform 1 0 34316 0 1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_365
timestamp 1704896540
transform 1 0 34684 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_377
timestamp 1704896540
transform 1 0 35788 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_389
timestamp 1704896540
transform 1 0 36892 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_401
timestamp 1704896540
transform 1 0 37996 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_413
timestamp 1704896540
transform 1 0 39100 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_419
timestamp 1704896540
transform 1 0 39652 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_68_421
timestamp 1704896540
transform 1 0 39836 0 1 39168
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_14
timestamp 1704896540
transform 1 0 2392 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_26
timestamp 1704896540
transform 1 0 3496 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_38
timestamp 1704896540
transform 1 0 4600 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_50
timestamp 1704896540
transform 1 0 5704 0 -1 40256
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_57
timestamp 1704896540
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_69
timestamp 1704896540
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_81
timestamp 1704896540
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_93
timestamp 1704896540
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_105
timestamp 1704896540
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_111
timestamp 1704896540
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_113
timestamp 1704896540
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_125
timestamp 1704896540
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_137
timestamp 1704896540
transform 1 0 13708 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_149
timestamp 1704896540
transform 1 0 14812 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_161
timestamp 1704896540
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_167
timestamp 1704896540
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_169
timestamp 1704896540
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_181
timestamp 1704896540
transform 1 0 17756 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_193
timestamp 1704896540
transform 1 0 18860 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_205
timestamp 1704896540
transform 1 0 19964 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_217
timestamp 1704896540
transform 1 0 21068 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_223
timestamp 1704896540
transform 1 0 21620 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_225
timestamp 1704896540
transform 1 0 21804 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_237
timestamp 1704896540
transform 1 0 22908 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_249
timestamp 1704896540
transform 1 0 24012 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_261
timestamp 1704896540
transform 1 0 25116 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_273
timestamp 1704896540
transform 1 0 26220 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_279
timestamp 1704896540
transform 1 0 26772 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_281
timestamp 1704896540
transform 1 0 26956 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_293
timestamp 1704896540
transform 1 0 28060 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_305
timestamp 1704896540
transform 1 0 29164 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_317
timestamp 1704896540
transform 1 0 30268 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_329
timestamp 1704896540
transform 1 0 31372 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_335
timestamp 1704896540
transform 1 0 31924 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_337
timestamp 1704896540
transform 1 0 32108 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_349
timestamp 1704896540
transform 1 0 33212 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_361
timestamp 1704896540
transform 1 0 34316 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_373
timestamp 1704896540
transform 1 0 35420 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_385
timestamp 1704896540
transform 1 0 36524 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_391
timestamp 1704896540
transform 1 0 37076 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_393
timestamp 1704896540
transform 1 0 37260 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_69_405
timestamp 1704896540
transform 1 0 38364 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_70_3
timestamp 1704896540
transform 1 0 1380 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_11
timestamp 1704896540
transform 1 0 2116 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_27
timestamp 1704896540
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_29
timestamp 1704896540
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_41
timestamp 1704896540
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_53
timestamp 1704896540
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_65
timestamp 1704896540
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_77
timestamp 1704896540
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_83
timestamp 1704896540
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_85
timestamp 1704896540
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_97
timestamp 1704896540
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_109
timestamp 1704896540
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_121
timestamp 1704896540
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_133
timestamp 1704896540
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_139
timestamp 1704896540
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_141
timestamp 1704896540
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_153
timestamp 1704896540
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_70_165
timestamp 1704896540
transform 1 0 16284 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_169
timestamp 1704896540
transform 1 0 16652 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_176
timestamp 1704896540
transform 1 0 17296 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_70_188
timestamp 1704896540
transform 1 0 18400 0 1 40256
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_197
timestamp 1704896540
transform 1 0 19228 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_209
timestamp 1704896540
transform 1 0 20332 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_70_221
timestamp 1704896540
transform 1 0 21436 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_229
timestamp 1704896540
transform 1 0 22172 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_245
timestamp 1704896540
transform 1 0 23644 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_251
timestamp 1704896540
transform 1 0 24196 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_253
timestamp 1704896540
transform 1 0 24380 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_263
timestamp 1704896540
transform 1 0 25300 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_275
timestamp 1704896540
transform 1 0 26404 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_287
timestamp 1704896540
transform 1 0 27508 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_70_299
timestamp 1704896540
transform 1 0 28612 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_307
timestamp 1704896540
transform 1 0 29348 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_309
timestamp 1704896540
transform 1 0 29532 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_70_321
timestamp 1704896540
transform 1 0 30636 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_70_329
timestamp 1704896540
transform 1 0 31372 0 1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_338
timestamp 1704896540
transform 1 0 32200 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_350
timestamp 1704896540
transform 1 0 33304 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_70_362
timestamp 1704896540
transform 1 0 34408 0 1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_365
timestamp 1704896540
transform 1 0 34684 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_377
timestamp 1704896540
transform 1 0 35788 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_389
timestamp 1704896540
transform 1 0 36892 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_70_401
timestamp 1704896540
transform 1 0 37996 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_70_415
timestamp 1704896540
transform 1 0 39284 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_419
timestamp 1704896540
transform 1 0 39652 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_70_421
timestamp 1704896540
transform 1 0 39836 0 1 40256
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_3
timestamp 1704896540
transform 1 0 1380 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_15
timestamp 1704896540
transform 1 0 2484 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_28
timestamp 1704896540
transform 1 0 3680 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_40
timestamp 1704896540
transform 1 0 4784 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_71_52
timestamp 1704896540
transform 1 0 5888 0 -1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_57
timestamp 1704896540
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_69
timestamp 1704896540
transform 1 0 7452 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_82
timestamp 1704896540
transform 1 0 8648 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_94
timestamp 1704896540
transform 1 0 9752 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_106
timestamp 1704896540
transform 1 0 10856 0 -1 41344
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_113
timestamp 1704896540
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_125
timestamp 1704896540
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_137
timestamp 1704896540
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_149
timestamp 1704896540
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_161
timestamp 1704896540
transform 1 0 15916 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_167
timestamp 1704896540
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_169
timestamp 1704896540
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_181
timestamp 1704896540
transform 1 0 17756 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_193
timestamp 1704896540
transform 1 0 18860 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_205
timestamp 1704896540
transform 1 0 19964 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_217
timestamp 1704896540
transform 1 0 21068 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_223
timestamp 1704896540
transform 1 0 21620 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_225
timestamp 1704896540
transform 1 0 21804 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_237
timestamp 1704896540
transform 1 0 22908 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_249
timestamp 1704896540
transform 1 0 24012 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_71_261
timestamp 1704896540
transform 1 0 25116 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_265
timestamp 1704896540
transform 1 0 25484 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_71_270
timestamp 1704896540
transform 1 0 25944 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_71_278
timestamp 1704896540
transform 1 0 26680 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_281
timestamp 1704896540
transform 1 0 26956 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_71_293
timestamp 1704896540
transform 1 0 28060 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_297
timestamp 1704896540
transform 1 0 28428 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_71_327
timestamp 1704896540
transform 1 0 31188 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_335
timestamp 1704896540
transform 1 0 31924 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_337
timestamp 1704896540
transform 1 0 32108 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_349
timestamp 1704896540
transform 1 0 33212 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_361
timestamp 1704896540
transform 1 0 34316 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_373
timestamp 1704896540
transform 1 0 35420 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_385
timestamp 1704896540
transform 1 0 36524 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_391
timestamp 1704896540
transform 1 0 37076 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_393
timestamp 1704896540
transform 1 0 37260 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_405
timestamp 1704896540
transform 1 0 38364 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_417
timestamp 1704896540
transform 1 0 39468 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_3
timestamp 1704896540
transform 1 0 1380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_15
timestamp 1704896540
transform 1 0 2484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_27
timestamp 1704896540
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_29
timestamp 1704896540
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_41
timestamp 1704896540
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_53
timestamp 1704896540
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_65
timestamp 1704896540
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_77
timestamp 1704896540
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_83
timestamp 1704896540
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_85
timestamp 1704896540
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_97
timestamp 1704896540
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_109
timestamp 1704896540
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_121
timestamp 1704896540
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_133
timestamp 1704896540
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_139
timestamp 1704896540
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_141
timestamp 1704896540
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_153
timestamp 1704896540
transform 1 0 15180 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_165
timestamp 1704896540
transform 1 0 16284 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_177
timestamp 1704896540
transform 1 0 17388 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_189
timestamp 1704896540
transform 1 0 18492 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_195
timestamp 1704896540
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_197
timestamp 1704896540
transform 1 0 19228 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_209
timestamp 1704896540
transform 1 0 20332 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_221
timestamp 1704896540
transform 1 0 21436 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_233
timestamp 1704896540
transform 1 0 22540 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_245
timestamp 1704896540
transform 1 0 23644 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_251
timestamp 1704896540
transform 1 0 24196 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_253
timestamp 1704896540
transform 1 0 24380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_265
timestamp 1704896540
transform 1 0 25484 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_277
timestamp 1704896540
transform 1 0 26588 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_289
timestamp 1704896540
transform 1 0 27692 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_301
timestamp 1704896540
transform 1 0 28796 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_307
timestamp 1704896540
transform 1 0 29348 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_309
timestamp 1704896540
transform 1 0 29532 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_321
timestamp 1704896540
transform 1 0 30636 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_72_333
timestamp 1704896540
transform 1 0 31740 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_357
timestamp 1704896540
transform 1 0 33948 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_363
timestamp 1704896540
transform 1 0 34500 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_365
timestamp 1704896540
transform 1 0 34684 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_377
timestamp 1704896540
transform 1 0 35788 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_389
timestamp 1704896540
transform 1 0 36892 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_401
timestamp 1704896540
transform 1 0 37996 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_413
timestamp 1704896540
transform 1 0 39100 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_419
timestamp 1704896540
transform 1 0 39652 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_72_421
timestamp 1704896540
transform 1 0 39836 0 1 41344
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_3
timestamp 1704896540
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_15
timestamp 1704896540
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_27
timestamp 1704896540
transform 1 0 3588 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_39
timestamp 1704896540
transform 1 0 4692 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_73_51
timestamp 1704896540
transform 1 0 5796 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_55
timestamp 1704896540
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_57
timestamp 1704896540
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_69
timestamp 1704896540
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_81
timestamp 1704896540
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_93
timestamp 1704896540
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_105
timestamp 1704896540
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_111
timestamp 1704896540
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_113
timestamp 1704896540
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_125
timestamp 1704896540
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_137
timestamp 1704896540
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_149
timestamp 1704896540
transform 1 0 14812 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_161
timestamp 1704896540
transform 1 0 15916 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_167
timestamp 1704896540
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_169
timestamp 1704896540
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_181
timestamp 1704896540
transform 1 0 17756 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_193
timestamp 1704896540
transform 1 0 18860 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_205
timestamp 1704896540
transform 1 0 19964 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_217
timestamp 1704896540
transform 1 0 21068 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_223
timestamp 1704896540
transform 1 0 21620 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_225
timestamp 1704896540
transform 1 0 21804 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_251
timestamp 1704896540
transform 1 0 24196 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_263
timestamp 1704896540
transform 1 0 25300 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_73_275
timestamp 1704896540
transform 1 0 26404 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_279
timestamp 1704896540
transform 1 0 26772 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_293
timestamp 1704896540
transform 1 0 28060 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_305
timestamp 1704896540
transform 1 0 29164 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_317
timestamp 1704896540
transform 1 0 30268 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_329
timestamp 1704896540
transform 1 0 31372 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_335
timestamp 1704896540
transform 1 0 31924 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_362
timestamp 1704896540
transform 1 0 34408 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_374
timestamp 1704896540
transform 1 0 35512 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_386
timestamp 1704896540
transform 1 0 36616 0 -1 42432
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_393
timestamp 1704896540
transform 1 0 37260 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_405
timestamp 1704896540
transform 1 0 38364 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_417
timestamp 1704896540
transform 1 0 39468 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_3
timestamp 1704896540
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_15
timestamp 1704896540
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_27
timestamp 1704896540
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_29
timestamp 1704896540
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_41
timestamp 1704896540
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_53
timestamp 1704896540
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_65
timestamp 1704896540
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_77
timestamp 1704896540
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_83
timestamp 1704896540
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_85
timestamp 1704896540
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_97
timestamp 1704896540
transform 1 0 10028 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_109
timestamp 1704896540
transform 1 0 11132 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_121
timestamp 1704896540
transform 1 0 12236 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_133
timestamp 1704896540
transform 1 0 13340 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_139
timestamp 1704896540
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_141
timestamp 1704896540
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_153
timestamp 1704896540
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_165
timestamp 1704896540
transform 1 0 16284 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_177
timestamp 1704896540
transform 1 0 17388 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_189
timestamp 1704896540
transform 1 0 18492 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_195
timestamp 1704896540
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_197
timestamp 1704896540
transform 1 0 19228 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_74_223
timestamp 1704896540
transform 1 0 21620 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_231
timestamp 1704896540
transform 1 0 22356 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_239
timestamp 1704896540
transform 1 0 23092 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_251
timestamp 1704896540
transform 1 0 24196 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_253
timestamp 1704896540
transform 1 0 24380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_265
timestamp 1704896540
transform 1 0 25484 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_277
timestamp 1704896540
transform 1 0 26588 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_289
timestamp 1704896540
transform 1 0 27692 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_301
timestamp 1704896540
transform 1 0 28796 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_307
timestamp 1704896540
transform 1 0 29348 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_309
timestamp 1704896540
transform 1 0 29532 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_321
timestamp 1704896540
transform 1 0 30636 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_333
timestamp 1704896540
transform 1 0 31740 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_345
timestamp 1704896540
transform 1 0 32844 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_357
timestamp 1704896540
transform 1 0 33948 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_363
timestamp 1704896540
transform 1 0 34500 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_365
timestamp 1704896540
transform 1 0 34684 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_377
timestamp 1704896540
transform 1 0 35788 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_389
timestamp 1704896540
transform 1 0 36892 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_401
timestamp 1704896540
transform 1 0 37996 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_413
timestamp 1704896540
transform 1 0 39100 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_419
timestamp 1704896540
transform 1 0 39652 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_74_421
timestamp 1704896540
transform 1 0 39836 0 1 42432
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_3
timestamp 1704896540
transform 1 0 1380 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_15
timestamp 1704896540
transform 1 0 2484 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_27
timestamp 1704896540
transform 1 0 3588 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_39
timestamp 1704896540
transform 1 0 4692 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_75_51
timestamp 1704896540
transform 1 0 5796 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_55
timestamp 1704896540
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_57
timestamp 1704896540
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_69
timestamp 1704896540
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_75_81
timestamp 1704896540
transform 1 0 8556 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_89
timestamp 1704896540
transform 1 0 9292 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_97
timestamp 1704896540
transform 1 0 10028 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_75_109
timestamp 1704896540
transform 1 0 11132 0 -1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_125
timestamp 1704896540
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_137
timestamp 1704896540
transform 1 0 13708 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_149
timestamp 1704896540
transform 1 0 14812 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_161
timestamp 1704896540
transform 1 0 15916 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_167
timestamp 1704896540
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_169
timestamp 1704896540
transform 1 0 16652 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_181
timestamp 1704896540
transform 1 0 17756 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_193
timestamp 1704896540
transform 1 0 18860 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_205
timestamp 1704896540
transform 1 0 19964 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_217
timestamp 1704896540
transform 1 0 21068 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_223
timestamp 1704896540
transform 1 0 21620 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_225
timestamp 1704896540
transform 1 0 21804 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_237
timestamp 1704896540
transform 1 0 22908 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_249
timestamp 1704896540
transform 1 0 24012 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_261
timestamp 1704896540
transform 1 0 25116 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_273
timestamp 1704896540
transform 1 0 26220 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_279
timestamp 1704896540
transform 1 0 26772 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_281
timestamp 1704896540
transform 1 0 26956 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_293
timestamp 1704896540
transform 1 0 28060 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_305
timestamp 1704896540
transform 1 0 29164 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_317
timestamp 1704896540
transform 1 0 30268 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_329
timestamp 1704896540
transform 1 0 31372 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_335
timestamp 1704896540
transform 1 0 31924 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_337
timestamp 1704896540
transform 1 0 32108 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_349
timestamp 1704896540
transform 1 0 33212 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_361
timestamp 1704896540
transform 1 0 34316 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_373
timestamp 1704896540
transform 1 0 35420 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_385
timestamp 1704896540
transform 1 0 36524 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_391
timestamp 1704896540
transform 1 0 37076 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_393
timestamp 1704896540
transform 1 0 37260 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_405
timestamp 1704896540
transform 1 0 38364 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_417
timestamp 1704896540
transform 1 0 39468 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_3
timestamp 1704896540
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_15
timestamp 1704896540
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_27
timestamp 1704896540
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_29
timestamp 1704896540
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_41
timestamp 1704896540
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_53
timestamp 1704896540
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_65
timestamp 1704896540
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_77
timestamp 1704896540
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_83
timestamp 1704896540
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_85
timestamp 1704896540
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_97
timestamp 1704896540
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_109
timestamp 1704896540
transform 1 0 11132 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_121
timestamp 1704896540
transform 1 0 12236 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_133
timestamp 1704896540
transform 1 0 13340 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_139
timestamp 1704896540
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_141
timestamp 1704896540
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_153
timestamp 1704896540
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_165
timestamp 1704896540
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_177
timestamp 1704896540
transform 1 0 17388 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_189
timestamp 1704896540
transform 1 0 18492 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_195
timestamp 1704896540
transform 1 0 19044 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_197
timestamp 1704896540
transform 1 0 19228 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_209
timestamp 1704896540
transform 1 0 20332 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_221
timestamp 1704896540
transform 1 0 21436 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_233
timestamp 1704896540
transform 1 0 22540 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_245
timestamp 1704896540
transform 1 0 23644 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_251
timestamp 1704896540
transform 1 0 24196 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_253
timestamp 1704896540
transform 1 0 24380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_265
timestamp 1704896540
transform 1 0 25484 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_277
timestamp 1704896540
transform 1 0 26588 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_289
timestamp 1704896540
transform 1 0 27692 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_301
timestamp 1704896540
transform 1 0 28796 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_307
timestamp 1704896540
transform 1 0 29348 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_309
timestamp 1704896540
transform 1 0 29532 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_321
timestamp 1704896540
transform 1 0 30636 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_333
timestamp 1704896540
transform 1 0 31740 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_345
timestamp 1704896540
transform 1 0 32844 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_357
timestamp 1704896540
transform 1 0 33948 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_363
timestamp 1704896540
transform 1 0 34500 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_365
timestamp 1704896540
transform 1 0 34684 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_377
timestamp 1704896540
transform 1 0 35788 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_389
timestamp 1704896540
transform 1 0 36892 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_401
timestamp 1704896540
transform 1 0 37996 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_413
timestamp 1704896540
transform 1 0 39100 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_419
timestamp 1704896540
transform 1 0 39652 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_76_421
timestamp 1704896540
transform 1 0 39836 0 1 43520
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_3
timestamp 1704896540
transform 1 0 1380 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_15
timestamp 1704896540
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_77_27
timestamp 1704896540
transform 1 0 3588 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77_35
timestamp 1704896540
transform 1 0 4324 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_77_45
timestamp 1704896540
transform 1 0 5244 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_77_53
timestamp 1704896540
transform 1 0 5980 0 -1 44608
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_57
timestamp 1704896540
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_69
timestamp 1704896540
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_81
timestamp 1704896540
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_93
timestamp 1704896540
transform 1 0 9660 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_77_103
timestamp 1704896540
transform 1 0 10580 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_111
timestamp 1704896540
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_113
timestamp 1704896540
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_125
timestamp 1704896540
transform 1 0 12604 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_137
timestamp 1704896540
transform 1 0 13708 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_149
timestamp 1704896540
transform 1 0 14812 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_161
timestamp 1704896540
transform 1 0 15916 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_167
timestamp 1704896540
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_169
timestamp 1704896540
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_77_181
timestamp 1704896540
transform 1 0 17756 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_189
timestamp 1704896540
transform 1 0 18492 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_199
timestamp 1704896540
transform 1 0 19412 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_211
timestamp 1704896540
transform 1 0 20516 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_223
timestamp 1704896540
transform 1 0 21620 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_225
timestamp 1704896540
transform 1 0 21804 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_237
timestamp 1704896540
transform 1 0 22908 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_249
timestamp 1704896540
transform 1 0 24012 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_261
timestamp 1704896540
transform 1 0 25116 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_273
timestamp 1704896540
transform 1 0 26220 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_279
timestamp 1704896540
transform 1 0 26772 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_281
timestamp 1704896540
transform 1 0 26956 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_293
timestamp 1704896540
transform 1 0 28060 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_305
timestamp 1704896540
transform 1 0 29164 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_317
timestamp 1704896540
transform 1 0 30268 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_329
timestamp 1704896540
transform 1 0 31372 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_335
timestamp 1704896540
transform 1 0 31924 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_337
timestamp 1704896540
transform 1 0 32108 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_349
timestamp 1704896540
transform 1 0 33212 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_361
timestamp 1704896540
transform 1 0 34316 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_373
timestamp 1704896540
transform 1 0 35420 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_385
timestamp 1704896540
transform 1 0 36524 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_391
timestamp 1704896540
transform 1 0 37076 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_409
timestamp 1704896540
transform 1 0 38732 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_77_421
timestamp 1704896540
transform 1 0 39836 0 -1 44608
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_3
timestamp 1704896540
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_15
timestamp 1704896540
transform 1 0 2484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_27
timestamp 1704896540
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_29
timestamp 1704896540
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_78_41
timestamp 1704896540
transform 1 0 4876 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_78_49
timestamp 1704896540
transform 1 0 5612 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_78_74
timestamp 1704896540
transform 1 0 7912 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_78_82
timestamp 1704896540
transform 1 0 8648 0 1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_85
timestamp 1704896540
transform 1 0 8924 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_97
timestamp 1704896540
transform 1 0 10028 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_109
timestamp 1704896540
transform 1 0 11132 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_121
timestamp 1704896540
transform 1 0 12236 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_133
timestamp 1704896540
transform 1 0 13340 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_139
timestamp 1704896540
transform 1 0 13892 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_141
timestamp 1704896540
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_153
timestamp 1704896540
transform 1 0 15180 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_165
timestamp 1704896540
transform 1 0 16284 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_177
timestamp 1704896540
transform 1 0 17388 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_189
timestamp 1704896540
transform 1 0 18492 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_195
timestamp 1704896540
transform 1 0 19044 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_197
timestamp 1704896540
transform 1 0 19228 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_204
timestamp 1704896540
transform 1 0 19872 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_216
timestamp 1704896540
transform 1 0 20976 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_228
timestamp 1704896540
transform 1 0 22080 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_240
timestamp 1704896540
transform 1 0 23184 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_253
timestamp 1704896540
transform 1 0 24380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_265
timestamp 1704896540
transform 1 0 25484 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_277
timestamp 1704896540
transform 1 0 26588 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_289
timestamp 1704896540
transform 1 0 27692 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_301
timestamp 1704896540
transform 1 0 28796 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_307
timestamp 1704896540
transform 1 0 29348 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_309
timestamp 1704896540
transform 1 0 29532 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_321
timestamp 1704896540
transform 1 0 30636 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_333
timestamp 1704896540
transform 1 0 31740 0 1 44608
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_346
timestamp 1704896540
transform 1 0 32936 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_358
timestamp 1704896540
transform 1 0 34040 0 1 44608
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_365
timestamp 1704896540
transform 1 0 34684 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_377
timestamp 1704896540
transform 1 0 35788 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_389
timestamp 1704896540
transform 1 0 36892 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_401
timestamp 1704896540
transform 1 0 37996 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_413
timestamp 1704896540
transform 1 0 39100 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_419
timestamp 1704896540
transform 1 0 39652 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_78_421
timestamp 1704896540
transform 1 0 39836 0 1 44608
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_3
timestamp 1704896540
transform 1 0 1380 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_15
timestamp 1704896540
transform 1 0 2484 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_27
timestamp 1704896540
transform 1 0 3588 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_39
timestamp 1704896540
transform 1 0 4692 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_79_51
timestamp 1704896540
transform 1 0 5796 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_55
timestamp 1704896540
transform 1 0 6164 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_79_62
timestamp 1704896540
transform 1 0 6808 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_68
timestamp 1704896540
transform 1 0 7360 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_80
timestamp 1704896540
transform 1 0 8464 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_92
timestamp 1704896540
transform 1 0 9568 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_79_104
timestamp 1704896540
transform 1 0 10672 0 -1 45696
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_113
timestamp 1704896540
transform 1 0 11500 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_125
timestamp 1704896540
transform 1 0 12604 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_137
timestamp 1704896540
transform 1 0 13708 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_149
timestamp 1704896540
transform 1 0 14812 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_79_161
timestamp 1704896540
transform 1 0 15916 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_167
timestamp 1704896540
transform 1 0 16468 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_169
timestamp 1704896540
transform 1 0 16652 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_181
timestamp 1704896540
transform 1 0 17756 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_193
timestamp 1704896540
transform 1 0 18860 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_205
timestamp 1704896540
transform 1 0 19964 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_79_217
timestamp 1704896540
transform 1 0 21068 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_223
timestamp 1704896540
transform 1 0 21620 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_225
timestamp 1704896540
transform 1 0 21804 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_79_237
timestamp 1704896540
transform 1 0 22908 0 -1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_260
timestamp 1704896540
transform 1 0 25024 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_79_272
timestamp 1704896540
transform 1 0 26128 0 -1 45696
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_281
timestamp 1704896540
transform 1 0 26956 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_293
timestamp 1704896540
transform 1 0 28060 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_305
timestamp 1704896540
transform 1 0 29164 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_317
timestamp 1704896540
transform 1 0 30268 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_79_329
timestamp 1704896540
transform 1 0 31372 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_335
timestamp 1704896540
transform 1 0 31924 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_337
timestamp 1704896540
transform 1 0 32108 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_349
timestamp 1704896540
transform 1 0 33212 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_361
timestamp 1704896540
transform 1 0 34316 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_373
timestamp 1704896540
transform 1 0 35420 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_79_385
timestamp 1704896540
transform 1 0 36524 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_391
timestamp 1704896540
transform 1 0 37076 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_393
timestamp 1704896540
transform 1 0 37260 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_405
timestamp 1704896540
transform 1 0 38364 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_417
timestamp 1704896540
transform 1 0 39468 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_3
timestamp 1704896540
transform 1 0 1380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_15
timestamp 1704896540
transform 1 0 2484 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_27
timestamp 1704896540
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_29
timestamp 1704896540
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_41
timestamp 1704896540
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_53
timestamp 1704896540
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_65
timestamp 1704896540
transform 1 0 7084 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80_77
timestamp 1704896540
transform 1 0 8188 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_83
timestamp 1704896540
transform 1 0 8740 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_85
timestamp 1704896540
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_97
timestamp 1704896540
transform 1 0 10028 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_109
timestamp 1704896540
transform 1 0 11132 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_121
timestamp 1704896540
transform 1 0 12236 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80_133
timestamp 1704896540
transform 1 0 13340 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_139
timestamp 1704896540
transform 1 0 13892 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_141
timestamp 1704896540
transform 1 0 14076 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_153
timestamp 1704896540
transform 1 0 15180 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_165
timestamp 1704896540
transform 1 0 16284 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_177
timestamp 1704896540
transform 1 0 17388 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80_189
timestamp 1704896540
transform 1 0 18492 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_195
timestamp 1704896540
transform 1 0 19044 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_197
timestamp 1704896540
transform 1 0 19228 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_209
timestamp 1704896540
transform 1 0 20332 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_221
timestamp 1704896540
transform 1 0 21436 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_233
timestamp 1704896540
transform 1 0 22540 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80_245
timestamp 1704896540
transform 1 0 23644 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_251
timestamp 1704896540
transform 1 0 24196 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_253
timestamp 1704896540
transform 1 0 24380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_265
timestamp 1704896540
transform 1 0 25484 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_277
timestamp 1704896540
transform 1 0 26588 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_289
timestamp 1704896540
transform 1 0 27692 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80_301
timestamp 1704896540
transform 1 0 28796 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_307
timestamp 1704896540
transform 1 0 29348 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_309
timestamp 1704896540
transform 1 0 29532 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_321
timestamp 1704896540
transform 1 0 30636 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_80_333
timestamp 1704896540
transform 1 0 31740 0 1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_346
timestamp 1704896540
transform 1 0 32936 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80_358
timestamp 1704896540
transform 1 0 34040 0 1 45696
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_365
timestamp 1704896540
transform 1 0 34684 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_377
timestamp 1704896540
transform 1 0 35788 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_389
timestamp 1704896540
transform 1 0 36892 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_401
timestamp 1704896540
transform 1 0 37996 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80_413
timestamp 1704896540
transform 1 0 39100 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_419
timestamp 1704896540
transform 1 0 39652 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_80_421
timestamp 1704896540
transform 1 0 39836 0 1 45696
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_3
timestamp 1704896540
transform 1 0 1380 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_15
timestamp 1704896540
transform 1 0 2484 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_27
timestamp 1704896540
transform 1 0 3588 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_39
timestamp 1704896540
transform 1 0 4692 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_81_51
timestamp 1704896540
transform 1 0 5796 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_55
timestamp 1704896540
transform 1 0 6164 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_57
timestamp 1704896540
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_69
timestamp 1704896540
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_81
timestamp 1704896540
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_93
timestamp 1704896540
transform 1 0 9660 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_81_105
timestamp 1704896540
transform 1 0 10764 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_111
timestamp 1704896540
transform 1 0 11316 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_113
timestamp 1704896540
transform 1 0 11500 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_125
timestamp 1704896540
transform 1 0 12604 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_137
timestamp 1704896540
transform 1 0 13708 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_149
timestamp 1704896540
transform 1 0 14812 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_81_161
timestamp 1704896540
transform 1 0 15916 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_167
timestamp 1704896540
transform 1 0 16468 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_169
timestamp 1704896540
transform 1 0 16652 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_181
timestamp 1704896540
transform 1 0 17756 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_193
timestamp 1704896540
transform 1 0 18860 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_205
timestamp 1704896540
transform 1 0 19964 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_81_217
timestamp 1704896540
transform 1 0 21068 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_223
timestamp 1704896540
transform 1 0 21620 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_225
timestamp 1704896540
transform 1 0 21804 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_237
timestamp 1704896540
transform 1 0 22908 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_249
timestamp 1704896540
transform 1 0 24012 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_261
timestamp 1704896540
transform 1 0 25116 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_81_273
timestamp 1704896540
transform 1 0 26220 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_279
timestamp 1704896540
transform 1 0 26772 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_281
timestamp 1704896540
transform 1 0 26956 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_293
timestamp 1704896540
transform 1 0 28060 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_305
timestamp 1704896540
transform 1 0 29164 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_317
timestamp 1704896540
transform 1 0 30268 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_81_329
timestamp 1704896540
transform 1 0 31372 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_335
timestamp 1704896540
transform 1 0 31924 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_337
timestamp 1704896540
transform 1 0 32108 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_349
timestamp 1704896540
transform 1 0 33212 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_361
timestamp 1704896540
transform 1 0 34316 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_373
timestamp 1704896540
transform 1 0 35420 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_81_385
timestamp 1704896540
transform 1 0 36524 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_391
timestamp 1704896540
transform 1 0 37076 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_393
timestamp 1704896540
transform 1 0 37260 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_405
timestamp 1704896540
transform 1 0 38364 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_417
timestamp 1704896540
transform 1 0 39468 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_3
timestamp 1704896540
transform 1 0 1380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_15
timestamp 1704896540
transform 1 0 2484 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_27
timestamp 1704896540
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_29
timestamp 1704896540
transform 1 0 3772 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_41
timestamp 1704896540
transform 1 0 4876 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_53
timestamp 1704896540
transform 1 0 5980 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_65
timestamp 1704896540
transform 1 0 7084 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_82_77
timestamp 1704896540
transform 1 0 8188 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_83
timestamp 1704896540
transform 1 0 8740 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_85
timestamp 1704896540
transform 1 0 8924 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_97
timestamp 1704896540
transform 1 0 10028 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_109
timestamp 1704896540
transform 1 0 11132 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_121
timestamp 1704896540
transform 1 0 12236 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_82_133
timestamp 1704896540
transform 1 0 13340 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_139
timestamp 1704896540
transform 1 0 13892 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_141
timestamp 1704896540
transform 1 0 14076 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_153
timestamp 1704896540
transform 1 0 15180 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_165
timestamp 1704896540
transform 1 0 16284 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_177
timestamp 1704896540
transform 1 0 17388 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_82_189
timestamp 1704896540
transform 1 0 18492 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_195
timestamp 1704896540
transform 1 0 19044 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_197
timestamp 1704896540
transform 1 0 19228 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_209
timestamp 1704896540
transform 1 0 20332 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_221
timestamp 1704896540
transform 1 0 21436 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_233
timestamp 1704896540
transform 1 0 22540 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_82_245
timestamp 1704896540
transform 1 0 23644 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_251
timestamp 1704896540
transform 1 0 24196 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_253
timestamp 1704896540
transform 1 0 24380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_265
timestamp 1704896540
transform 1 0 25484 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_277
timestamp 1704896540
transform 1 0 26588 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_289
timestamp 1704896540
transform 1 0 27692 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_82_301
timestamp 1704896540
transform 1 0 28796 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_307
timestamp 1704896540
transform 1 0 29348 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_309
timestamp 1704896540
transform 1 0 29532 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_321
timestamp 1704896540
transform 1 0 30636 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_333
timestamp 1704896540
transform 1 0 31740 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_345
timestamp 1704896540
transform 1 0 32844 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_82_357
timestamp 1704896540
transform 1 0 33948 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_363
timestamp 1704896540
transform 1 0 34500 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_365
timestamp 1704896540
transform 1 0 34684 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_377
timestamp 1704896540
transform 1 0 35788 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_389
timestamp 1704896540
transform 1 0 36892 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_401
timestamp 1704896540
transform 1 0 37996 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_82_413
timestamp 1704896540
transform 1 0 39100 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_419
timestamp 1704896540
transform 1 0 39652 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_82_421
timestamp 1704896540
transform 1 0 39836 0 1 46784
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_3
timestamp 1704896540
transform 1 0 1380 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_15
timestamp 1704896540
transform 1 0 2484 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_27
timestamp 1704896540
transform 1 0 3588 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_39
timestamp 1704896540
transform 1 0 4692 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_83_51
timestamp 1704896540
transform 1 0 5796 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_55
timestamp 1704896540
transform 1 0 6164 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_57
timestamp 1704896540
transform 1 0 6348 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_69
timestamp 1704896540
transform 1 0 7452 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_81
timestamp 1704896540
transform 1 0 8556 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_93
timestamp 1704896540
transform 1 0 9660 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_83_105
timestamp 1704896540
transform 1 0 10764 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_111
timestamp 1704896540
transform 1 0 11316 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_113
timestamp 1704896540
transform 1 0 11500 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_125
timestamp 1704896540
transform 1 0 12604 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_137
timestamp 1704896540
transform 1 0 13708 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_149
timestamp 1704896540
transform 1 0 14812 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_83_161
timestamp 1704896540
transform 1 0 15916 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_167
timestamp 1704896540
transform 1 0 16468 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_169
timestamp 1704896540
transform 1 0 16652 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_181
timestamp 1704896540
transform 1 0 17756 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_193
timestamp 1704896540
transform 1 0 18860 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_205
timestamp 1704896540
transform 1 0 19964 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_83_217
timestamp 1704896540
transform 1 0 21068 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_223
timestamp 1704896540
transform 1 0 21620 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_225
timestamp 1704896540
transform 1 0 21804 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_237
timestamp 1704896540
transform 1 0 22908 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_249
timestamp 1704896540
transform 1 0 24012 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_261
timestamp 1704896540
transform 1 0 25116 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_83_273
timestamp 1704896540
transform 1 0 26220 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_279
timestamp 1704896540
transform 1 0 26772 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_281
timestamp 1704896540
transform 1 0 26956 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_293
timestamp 1704896540
transform 1 0 28060 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_305
timestamp 1704896540
transform 1 0 29164 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_83_317
timestamp 1704896540
transform 1 0 30268 0 -1 47872
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_337
timestamp 1704896540
transform 1 0 32108 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_349
timestamp 1704896540
transform 1 0 33212 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_361
timestamp 1704896540
transform 1 0 34316 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_373
timestamp 1704896540
transform 1 0 35420 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_83_385
timestamp 1704896540
transform 1 0 36524 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_391
timestamp 1704896540
transform 1 0 37076 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_393
timestamp 1704896540
transform 1 0 37260 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_405
timestamp 1704896540
transform 1 0 38364 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_417
timestamp 1704896540
transform 1 0 39468 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_3
timestamp 1704896540
transform 1 0 1380 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_15
timestamp 1704896540
transform 1 0 2484 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_27
timestamp 1704896540
transform 1 0 3588 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_29
timestamp 1704896540
transform 1 0 3772 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_41
timestamp 1704896540
transform 1 0 4876 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_53
timestamp 1704896540
transform 1 0 5980 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_65
timestamp 1704896540
transform 1 0 7084 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_77
timestamp 1704896540
transform 1 0 8188 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_83
timestamp 1704896540
transform 1 0 8740 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_85
timestamp 1704896540
transform 1 0 8924 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_97
timestamp 1704896540
transform 1 0 10028 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_109
timestamp 1704896540
transform 1 0 11132 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_121
timestamp 1704896540
transform 1 0 12236 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_133
timestamp 1704896540
transform 1 0 13340 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_139
timestamp 1704896540
transform 1 0 13892 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_141
timestamp 1704896540
transform 1 0 14076 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_153
timestamp 1704896540
transform 1 0 15180 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_165
timestamp 1704896540
transform 1 0 16284 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_177
timestamp 1704896540
transform 1 0 17388 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_189
timestamp 1704896540
transform 1 0 18492 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_195
timestamp 1704896540
transform 1 0 19044 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_197
timestamp 1704896540
transform 1 0 19228 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_209
timestamp 1704896540
transform 1 0 20332 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_221
timestamp 1704896540
transform 1 0 21436 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_233
timestamp 1704896540
transform 1 0 22540 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_245
timestamp 1704896540
transform 1 0 23644 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_251
timestamp 1704896540
transform 1 0 24196 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_253
timestamp 1704896540
transform 1 0 24380 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_265
timestamp 1704896540
transform 1 0 25484 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_277
timestamp 1704896540
transform 1 0 26588 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_289
timestamp 1704896540
transform 1 0 27692 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_301
timestamp 1704896540
transform 1 0 28796 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_307
timestamp 1704896540
transform 1 0 29348 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_309
timestamp 1704896540
transform 1 0 29532 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_321
timestamp 1704896540
transform 1 0 30636 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_333
timestamp 1704896540
transform 1 0 31740 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_345
timestamp 1704896540
transform 1 0 32844 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_357
timestamp 1704896540
transform 1 0 33948 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_363
timestamp 1704896540
transform 1 0 34500 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_365
timestamp 1704896540
transform 1 0 34684 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_377
timestamp 1704896540
transform 1 0 35788 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_389
timestamp 1704896540
transform 1 0 36892 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_401
timestamp 1704896540
transform 1 0 37996 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_413
timestamp 1704896540
transform 1 0 39100 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_419
timestamp 1704896540
transform 1 0 39652 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_84_421
timestamp 1704896540
transform 1 0 39836 0 1 47872
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_3
timestamp 1704896540
transform 1 0 1380 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_15
timestamp 1704896540
transform 1 0 2484 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_27
timestamp 1704896540
transform 1 0 3588 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_39
timestamp 1704896540
transform 1 0 4692 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_85_51
timestamp 1704896540
transform 1 0 5796 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_55
timestamp 1704896540
transform 1 0 6164 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_57
timestamp 1704896540
transform 1 0 6348 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_69
timestamp 1704896540
transform 1 0 7452 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_81
timestamp 1704896540
transform 1 0 8556 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85_93
timestamp 1704896540
transform 1 0 9660 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85_106
timestamp 1704896540
transform 1 0 10856 0 -1 48960
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_113
timestamp 1704896540
transform 1 0 11500 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_125
timestamp 1704896540
transform 1 0 12604 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_137
timestamp 1704896540
transform 1 0 13708 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_149
timestamp 1704896540
transform 1 0 14812 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85_161
timestamp 1704896540
transform 1 0 15916 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_167
timestamp 1704896540
transform 1 0 16468 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_169
timestamp 1704896540
transform 1 0 16652 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_177
timestamp 1704896540
transform 1 0 17388 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_189
timestamp 1704896540
transform 1 0 18492 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_201
timestamp 1704896540
transform 1 0 19596 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_85_213
timestamp 1704896540
transform 1 0 20700 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_85_221
timestamp 1704896540
transform 1 0 21436 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85_225
timestamp 1704896540
transform 1 0 21804 0 -1 48960
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_234
timestamp 1704896540
transform 1 0 22632 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_246
timestamp 1704896540
transform 1 0 23736 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_258
timestamp 1704896540
transform 1 0 24840 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_85_270
timestamp 1704896540
transform 1 0 25944 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85_278
timestamp 1704896540
transform 1 0 26680 0 -1 48960
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_281
timestamp 1704896540
transform 1 0 26956 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_293
timestamp 1704896540
transform 1 0 28060 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_305
timestamp 1704896540
transform 1 0 29164 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_317
timestamp 1704896540
transform 1 0 30268 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85_329
timestamp 1704896540
transform 1 0 31372 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_335
timestamp 1704896540
transform 1 0 31924 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_337
timestamp 1704896540
transform 1 0 32108 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_349
timestamp 1704896540
transform 1 0 33212 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_361
timestamp 1704896540
transform 1 0 34316 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_373
timestamp 1704896540
transform 1 0 35420 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85_385
timestamp 1704896540
transform 1 0 36524 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_391
timestamp 1704896540
transform 1 0 37076 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_402
timestamp 1704896540
transform 1 0 38088 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_414
timestamp 1704896540
transform 1 0 39192 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_85_426
timestamp 1704896540
transform 1 0 40296 0 -1 48960
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_3
timestamp 1704896540
transform 1 0 1380 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_15
timestamp 1704896540
transform 1 0 2484 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_27
timestamp 1704896540
transform 1 0 3588 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_29
timestamp 1704896540
transform 1 0 3772 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_41
timestamp 1704896540
transform 1 0 4876 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_53
timestamp 1704896540
transform 1 0 5980 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_65
timestamp 1704896540
transform 1 0 7084 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_86_77
timestamp 1704896540
transform 1 0 8188 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_83
timestamp 1704896540
transform 1 0 8740 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_85
timestamp 1704896540
transform 1 0 8924 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_97
timestamp 1704896540
transform 1 0 10028 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_109
timestamp 1704896540
transform 1 0 11132 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_121
timestamp 1704896540
transform 1 0 12236 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_86_133
timestamp 1704896540
transform 1 0 13340 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_139
timestamp 1704896540
transform 1 0 13892 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_141
timestamp 1704896540
transform 1 0 14076 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_153
timestamp 1704896540
transform 1 0 15180 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_165
timestamp 1704896540
transform 1 0 16284 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_177
timestamp 1704896540
transform 1 0 17388 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_86_189
timestamp 1704896540
transform 1 0 18492 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_195
timestamp 1704896540
transform 1 0 19044 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_197
timestamp 1704896540
transform 1 0 19228 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_209
timestamp 1704896540
transform 1 0 20332 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_221
timestamp 1704896540
transform 1 0 21436 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_233
timestamp 1704896540
transform 1 0 22540 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_86_245
timestamp 1704896540
transform 1 0 23644 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_251
timestamp 1704896540
transform 1 0 24196 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_260
timestamp 1704896540
transform 1 0 25024 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_272
timestamp 1704896540
transform 1 0 26128 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_284
timestamp 1704896540
transform 1 0 27232 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_296
timestamp 1704896540
transform 1 0 28336 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_309
timestamp 1704896540
transform 1 0 29532 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_321
timestamp 1704896540
transform 1 0 30636 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_333
timestamp 1704896540
transform 1 0 31740 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_345
timestamp 1704896540
transform 1 0 32844 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_86_357
timestamp 1704896540
transform 1 0 33948 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_363
timestamp 1704896540
transform 1 0 34500 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_365
timestamp 1704896540
transform 1 0 34684 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_377
timestamp 1704896540
transform 1 0 35788 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_389
timestamp 1704896540
transform 1 0 36892 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_401
timestamp 1704896540
transform 1 0 37996 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_86_413
timestamp 1704896540
transform 1 0 39100 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_419
timestamp 1704896540
transform 1 0 39652 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_86_421
timestamp 1704896540
transform 1 0 39836 0 1 48960
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_19
timestamp 1704896540
transform 1 0 2852 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_31
timestamp 1704896540
transform 1 0 3956 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_43
timestamp 1704896540
transform 1 0 5060 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_55
timestamp 1704896540
transform 1 0 6164 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_57
timestamp 1704896540
transform 1 0 6348 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_69
timestamp 1704896540
transform 1 0 7452 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_81
timestamp 1704896540
transform 1 0 8556 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_93
timestamp 1704896540
transform 1 0 9660 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87_105
timestamp 1704896540
transform 1 0 10764 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_111
timestamp 1704896540
transform 1 0 11316 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_113
timestamp 1704896540
transform 1 0 11500 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_125
timestamp 1704896540
transform 1 0 12604 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_146
timestamp 1704896540
transform 1 0 14536 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_87_158
timestamp 1704896540
transform 1 0 15640 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_87_166
timestamp 1704896540
transform 1 0 16376 0 -1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_169
timestamp 1704896540
transform 1 0 16652 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_181
timestamp 1704896540
transform 1 0 17756 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_193
timestamp 1704896540
transform 1 0 18860 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_205
timestamp 1704896540
transform 1 0 19964 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87_217
timestamp 1704896540
transform 1 0 21068 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_223
timestamp 1704896540
transform 1 0 21620 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_225
timestamp 1704896540
transform 1 0 21804 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87_237
timestamp 1704896540
transform 1 0 22908 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_243
timestamp 1704896540
transform 1 0 23460 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_261
timestamp 1704896540
transform 1 0 25116 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87_273
timestamp 1704896540
transform 1 0 26220 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_279
timestamp 1704896540
transform 1 0 26772 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_281
timestamp 1704896540
transform 1 0 26956 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_293
timestamp 1704896540
transform 1 0 28060 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_305
timestamp 1704896540
transform 1 0 29164 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_317
timestamp 1704896540
transform 1 0 30268 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87_329
timestamp 1704896540
transform 1 0 31372 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_335
timestamp 1704896540
transform 1 0 31924 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_337
timestamp 1704896540
transform 1 0 32108 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_349
timestamp 1704896540
transform 1 0 33212 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_361
timestamp 1704896540
transform 1 0 34316 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_87_373
timestamp 1704896540
transform 1 0 35420 0 -1 50048
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_393
timestamp 1704896540
transform 1 0 37260 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_405
timestamp 1704896540
transform 1 0 38364 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_417
timestamp 1704896540
transform 1 0 39468 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_88_3
timestamp 1704896540
transform 1 0 1380 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_88_24
timestamp 1704896540
transform 1 0 3312 0 1 50048
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_29
timestamp 1704896540
transform 1 0 3772 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_41
timestamp 1704896540
transform 1 0 4876 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_53
timestamp 1704896540
transform 1 0 5980 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_65
timestamp 1704896540
transform 1 0 7084 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_88_77
timestamp 1704896540
transform 1 0 8188 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_83
timestamp 1704896540
transform 1 0 8740 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_85
timestamp 1704896540
transform 1 0 8924 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_97
timestamp 1704896540
transform 1 0 10028 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_109
timestamp 1704896540
transform 1 0 11132 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_88_121
timestamp 1704896540
transform 1 0 12236 0 1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_127
timestamp 1704896540
transform 1 0 12788 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_139
timestamp 1704896540
transform 1 0 13892 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_141
timestamp 1704896540
transform 1 0 14076 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_153
timestamp 1704896540
transform 1 0 15180 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_165
timestamp 1704896540
transform 1 0 16284 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_177
timestamp 1704896540
transform 1 0 17388 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_88_189
timestamp 1704896540
transform 1 0 18492 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_195
timestamp 1704896540
transform 1 0 19044 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_197
timestamp 1704896540
transform 1 0 19228 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_209
timestamp 1704896540
transform 1 0 20332 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_221
timestamp 1704896540
transform 1 0 21436 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_233
timestamp 1704896540
transform 1 0 22540 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_88_245
timestamp 1704896540
transform 1 0 23644 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_251
timestamp 1704896540
transform 1 0 24196 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_253
timestamp 1704896540
transform 1 0 24380 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_265
timestamp 1704896540
transform 1 0 25484 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_277
timestamp 1704896540
transform 1 0 26588 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_289
timestamp 1704896540
transform 1 0 27692 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_88_301
timestamp 1704896540
transform 1 0 28796 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_307
timestamp 1704896540
transform 1 0 29348 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_309
timestamp 1704896540
transform 1 0 29532 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_321
timestamp 1704896540
transform 1 0 30636 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_333
timestamp 1704896540
transform 1 0 31740 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_345
timestamp 1704896540
transform 1 0 32844 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_88_357
timestamp 1704896540
transform 1 0 33948 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_363
timestamp 1704896540
transform 1 0 34500 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_365
timestamp 1704896540
transform 1 0 34684 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_377
timestamp 1704896540
transform 1 0 35788 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_389
timestamp 1704896540
transform 1 0 36892 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_401
timestamp 1704896540
transform 1 0 37996 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_88_413
timestamp 1704896540
transform 1 0 39100 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_419
timestamp 1704896540
transform 1 0 39652 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_88_421
timestamp 1704896540
transform 1 0 39836 0 1 50048
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_3
timestamp 1704896540
transform 1 0 1380 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_15
timestamp 1704896540
transform 1 0 2484 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_27
timestamp 1704896540
transform 1 0 3588 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_39
timestamp 1704896540
transform 1 0 4692 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_89_51
timestamp 1704896540
transform 1 0 5796 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_55
timestamp 1704896540
transform 1 0 6164 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_57
timestamp 1704896540
transform 1 0 6348 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_69
timestamp 1704896540
transform 1 0 7452 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_81
timestamp 1704896540
transform 1 0 8556 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_89_93
timestamp 1704896540
transform 1 0 9660 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_97
timestamp 1704896540
transform 1 0 10028 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_111
timestamp 1704896540
transform 1 0 11316 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_89_113
timestamp 1704896540
transform 1 0 11500 0 -1 51136
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_134
timestamp 1704896540
transform 1 0 13432 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_146
timestamp 1704896540
transform 1 0 14536 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_89_158
timestamp 1704896540
transform 1 0 15640 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_89_166
timestamp 1704896540
transform 1 0 16376 0 -1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_169
timestamp 1704896540
transform 1 0 16652 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_181
timestamp 1704896540
transform 1 0 17756 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_193
timestamp 1704896540
transform 1 0 18860 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_205
timestamp 1704896540
transform 1 0 19964 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_89_217
timestamp 1704896540
transform 1 0 21068 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_223
timestamp 1704896540
transform 1 0 21620 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_234
timestamp 1704896540
transform 1 0 22632 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_246
timestamp 1704896540
transform 1 0 23736 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_258
timestamp 1704896540
transform 1 0 24840 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_89_270
timestamp 1704896540
transform 1 0 25944 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_89_278
timestamp 1704896540
transform 1 0 26680 0 -1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_281
timestamp 1704896540
transform 1 0 26956 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_293
timestamp 1704896540
transform 1 0 28060 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_305
timestamp 1704896540
transform 1 0 29164 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_317
timestamp 1704896540
transform 1 0 30268 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_89_329
timestamp 1704896540
transform 1 0 31372 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_335
timestamp 1704896540
transform 1 0 31924 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_337
timestamp 1704896540
transform 1 0 32108 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_349
timestamp 1704896540
transform 1 0 33212 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_361
timestamp 1704896540
transform 1 0 34316 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_373
timestamp 1704896540
transform 1 0 35420 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_89_385
timestamp 1704896540
transform 1 0 36524 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_391
timestamp 1704896540
transform 1 0 37076 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_393
timestamp 1704896540
transform 1 0 37260 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_405
timestamp 1704896540
transform 1 0 38364 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_417
timestamp 1704896540
transform 1 0 39468 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_3
timestamp 1704896540
transform 1 0 1380 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_15
timestamp 1704896540
transform 1 0 2484 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_27
timestamp 1704896540
transform 1 0 3588 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_29
timestamp 1704896540
transform 1 0 3772 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_41
timestamp 1704896540
transform 1 0 4876 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_53
timestamp 1704896540
transform 1 0 5980 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_65
timestamp 1704896540
transform 1 0 7084 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_90_77
timestamp 1704896540
transform 1 0 8188 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_83
timestamp 1704896540
transform 1 0 8740 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_85
timestamp 1704896540
transform 1 0 8924 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_97
timestamp 1704896540
transform 1 0 10028 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_109
timestamp 1704896540
transform 1 0 11132 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_121
timestamp 1704896540
transform 1 0 12236 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_90_133
timestamp 1704896540
transform 1 0 13340 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_139
timestamp 1704896540
transform 1 0 13892 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_141
timestamp 1704896540
transform 1 0 14076 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_153
timestamp 1704896540
transform 1 0 15180 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_165
timestamp 1704896540
transform 1 0 16284 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_177
timestamp 1704896540
transform 1 0 17388 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_90_189
timestamp 1704896540
transform 1 0 18492 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_195
timestamp 1704896540
transform 1 0 19044 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_197
timestamp 1704896540
transform 1 0 19228 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_209
timestamp 1704896540
transform 1 0 20332 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_221
timestamp 1704896540
transform 1 0 21436 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_233
timestamp 1704896540
transform 1 0 22540 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_90_245
timestamp 1704896540
transform 1 0 23644 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_251
timestamp 1704896540
transform 1 0 24196 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_253
timestamp 1704896540
transform 1 0 24380 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_265
timestamp 1704896540
transform 1 0 25484 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_277
timestamp 1704896540
transform 1 0 26588 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_289
timestamp 1704896540
transform 1 0 27692 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_90_301
timestamp 1704896540
transform 1 0 28796 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_307
timestamp 1704896540
transform 1 0 29348 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_309
timestamp 1704896540
transform 1 0 29532 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_90_321
timestamp 1704896540
transform 1 0 30636 0 1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_345
timestamp 1704896540
transform 1 0 32844 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_90_357
timestamp 1704896540
transform 1 0 33948 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_363
timestamp 1704896540
transform 1 0 34500 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_365
timestamp 1704896540
transform 1 0 34684 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_377
timestamp 1704896540
transform 1 0 35788 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_389
timestamp 1704896540
transform 1 0 36892 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_401
timestamp 1704896540
transform 1 0 37996 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_90_413
timestamp 1704896540
transform 1 0 39100 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_419
timestamp 1704896540
transform 1 0 39652 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_90_421
timestamp 1704896540
transform 1 0 39836 0 1 51136
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_3
timestamp 1704896540
transform 1 0 1380 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_15
timestamp 1704896540
transform 1 0 2484 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_91_27
timestamp 1704896540
transform 1 0 3588 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_33
timestamp 1704896540
transform 1 0 4140 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_91_48
timestamp 1704896540
transform 1 0 5520 0 -1 52224
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_57
timestamp 1704896540
transform 1 0 6348 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_69
timestamp 1704896540
transform 1 0 7452 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_81
timestamp 1704896540
transform 1 0 8556 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_93
timestamp 1704896540
transform 1 0 9660 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_91_105
timestamp 1704896540
transform 1 0 10764 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_111
timestamp 1704896540
transform 1 0 11316 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_113
timestamp 1704896540
transform 1 0 11500 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_125
timestamp 1704896540
transform 1 0 12604 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_137
timestamp 1704896540
transform 1 0 13708 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_149
timestamp 1704896540
transform 1 0 14812 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_91_161
timestamp 1704896540
transform 1 0 15916 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_167
timestamp 1704896540
transform 1 0 16468 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_169
timestamp 1704896540
transform 1 0 16652 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_181
timestamp 1704896540
transform 1 0 17756 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_193
timestamp 1704896540
transform 1 0 18860 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_91_205
timestamp 1704896540
transform 1 0 19964 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_91_213
timestamp 1704896540
transform 1 0 20700 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_223
timestamp 1704896540
transform 1 0 21620 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_225
timestamp 1704896540
transform 1 0 21804 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_237
timestamp 1704896540
transform 1 0 22908 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_249
timestamp 1704896540
transform 1 0 24012 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_261
timestamp 1704896540
transform 1 0 25116 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_91_273
timestamp 1704896540
transform 1 0 26220 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_279
timestamp 1704896540
transform 1 0 26772 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_281
timestamp 1704896540
transform 1 0 26956 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_293
timestamp 1704896540
transform 1 0 28060 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_305
timestamp 1704896540
transform 1 0 29164 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_317
timestamp 1704896540
transform 1 0 30268 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_91_329
timestamp 1704896540
transform 1 0 31372 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_335
timestamp 1704896540
transform 1 0 31924 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_337
timestamp 1704896540
transform 1 0 32108 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_349
timestamp 1704896540
transform 1 0 33212 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_361
timestamp 1704896540
transform 1 0 34316 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_91_373
timestamp 1704896540
transform 1 0 35420 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_91_383
timestamp 1704896540
transform 1 0 36340 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_391
timestamp 1704896540
transform 1 0 37076 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_393
timestamp 1704896540
transform 1 0 37260 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_405
timestamp 1704896540
transform 1 0 38364 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_417
timestamp 1704896540
transform 1 0 39468 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_3
timestamp 1704896540
transform 1 0 1380 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_15
timestamp 1704896540
transform 1 0 2484 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_27
timestamp 1704896540
transform 1 0 3588 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_29
timestamp 1704896540
transform 1 0 3772 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_92_41
timestamp 1704896540
transform 1 0 4876 0 1 52224
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_69
timestamp 1704896540
transform 1 0 7452 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_92_81
timestamp 1704896540
transform 1 0 8556 0 1 52224
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_85
timestamp 1704896540
transform 1 0 8924 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_97
timestamp 1704896540
transform 1 0 10028 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_109
timestamp 1704896540
transform 1 0 11132 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_121
timestamp 1704896540
transform 1 0 12236 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_92_133
timestamp 1704896540
transform 1 0 13340 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_139
timestamp 1704896540
transform 1 0 13892 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_141
timestamp 1704896540
transform 1 0 14076 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_153
timestamp 1704896540
transform 1 0 15180 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_165
timestamp 1704896540
transform 1 0 16284 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_177
timestamp 1704896540
transform 1 0 17388 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_92_189
timestamp 1704896540
transform 1 0 18492 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_195
timestamp 1704896540
transform 1 0 19044 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_197
timestamp 1704896540
transform 1 0 19228 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_209
timestamp 1704896540
transform 1 0 20332 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_221
timestamp 1704896540
transform 1 0 21436 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_233
timestamp 1704896540
transform 1 0 22540 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_92_245
timestamp 1704896540
transform 1 0 23644 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_251
timestamp 1704896540
transform 1 0 24196 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_253
timestamp 1704896540
transform 1 0 24380 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_265
timestamp 1704896540
transform 1 0 25484 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_277
timestamp 1704896540
transform 1 0 26588 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_289
timestamp 1704896540
transform 1 0 27692 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_92_301
timestamp 1704896540
transform 1 0 28796 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_307
timestamp 1704896540
transform 1 0 29348 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_309
timestamp 1704896540
transform 1 0 29532 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_321
timestamp 1704896540
transform 1 0 30636 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_333
timestamp 1704896540
transform 1 0 31740 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_345
timestamp 1704896540
transform 1 0 32844 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_92_357
timestamp 1704896540
transform 1 0 33948 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_363
timestamp 1704896540
transform 1 0 34500 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_92_372
timestamp 1704896540
transform 1 0 35328 0 1 52224
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_388
timestamp 1704896540
transform 1 0 36800 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_92_400
timestamp 1704896540
transform 1 0 37904 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_92_408
timestamp 1704896540
transform 1 0 38640 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_92_417
timestamp 1704896540
transform 1 0 39468 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_92_421
timestamp 1704896540
transform 1 0 39836 0 1 52224
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_3
timestamp 1704896540
transform 1 0 1380 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_15
timestamp 1704896540
transform 1 0 2484 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_27
timestamp 1704896540
transform 1 0 3588 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_39
timestamp 1704896540
transform 1 0 4692 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_93_51
timestamp 1704896540
transform 1 0 5796 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_55
timestamp 1704896540
transform 1 0 6164 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_57
timestamp 1704896540
transform 1 0 6348 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_69
timestamp 1704896540
transform 1 0 7452 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_81
timestamp 1704896540
transform 1 0 8556 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_93
timestamp 1704896540
transform 1 0 9660 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_93_105
timestamp 1704896540
transform 1 0 10764 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_111
timestamp 1704896540
transform 1 0 11316 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_113
timestamp 1704896540
transform 1 0 11500 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_125
timestamp 1704896540
transform 1 0 12604 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_137
timestamp 1704896540
transform 1 0 13708 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_93_149
timestamp 1704896540
transform 1 0 14812 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_93_164
timestamp 1704896540
transform 1 0 16192 0 -1 53312
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_169
timestamp 1704896540
transform 1 0 16652 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_181
timestamp 1704896540
transform 1 0 17756 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_193
timestamp 1704896540
transform 1 0 18860 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_205
timestamp 1704896540
transform 1 0 19964 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_93_217
timestamp 1704896540
transform 1 0 21068 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_223
timestamp 1704896540
transform 1 0 21620 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_225
timestamp 1704896540
transform 1 0 21804 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_237
timestamp 1704896540
transform 1 0 22908 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_249
timestamp 1704896540
transform 1 0 24012 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_261
timestamp 1704896540
transform 1 0 25116 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_93_273
timestamp 1704896540
transform 1 0 26220 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_279
timestamp 1704896540
transform 1 0 26772 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_281
timestamp 1704896540
transform 1 0 26956 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_293
timestamp 1704896540
transform 1 0 28060 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_305
timestamp 1704896540
transform 1 0 29164 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_317
timestamp 1704896540
transform 1 0 30268 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_93_329
timestamp 1704896540
transform 1 0 31372 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_335
timestamp 1704896540
transform 1 0 31924 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_337
timestamp 1704896540
transform 1 0 32108 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_349
timestamp 1704896540
transform 1 0 33212 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_361
timestamp 1704896540
transform 1 0 34316 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_373
timestamp 1704896540
transform 1 0 35420 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_385
timestamp 1704896540
transform 1 0 36524 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_391
timestamp 1704896540
transform 1 0 37076 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_393
timestamp 1704896540
transform 1 0 37260 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_405
timestamp 1704896540
transform 1 0 38364 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_417
timestamp 1704896540
transform 1 0 39468 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_3
timestamp 1704896540
transform 1 0 1380 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_15
timestamp 1704896540
transform 1 0 2484 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_27
timestamp 1704896540
transform 1 0 3588 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_38
timestamp 1704896540
transform 1 0 4600 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_50
timestamp 1704896540
transform 1 0 5704 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_62
timestamp 1704896540
transform 1 0 6808 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_94_74
timestamp 1704896540
transform 1 0 7912 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_94_82
timestamp 1704896540
transform 1 0 8648 0 1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_85
timestamp 1704896540
transform 1 0 8924 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_97
timestamp 1704896540
transform 1 0 10028 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_109
timestamp 1704896540
transform 1 0 11132 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_121
timestamp 1704896540
transform 1 0 12236 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94_133
timestamp 1704896540
transform 1 0 13340 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_139
timestamp 1704896540
transform 1 0 13892 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_94_141
timestamp 1704896540
transform 1 0 14076 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_94_149
timestamp 1704896540
transform 1 0 14812 0 1 53312
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_161
timestamp 1704896540
transform 1 0 15916 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_173
timestamp 1704896540
transform 1 0 17020 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_94_185
timestamp 1704896540
transform 1 0 18124 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_94_193
timestamp 1704896540
transform 1 0 18860 0 1 53312
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_197
timestamp 1704896540
transform 1 0 19228 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_209
timestamp 1704896540
transform 1 0 20332 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_221
timestamp 1704896540
transform 1 0 21436 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_233
timestamp 1704896540
transform 1 0 22540 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94_245
timestamp 1704896540
transform 1 0 23644 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_251
timestamp 1704896540
transform 1 0 24196 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_253
timestamp 1704896540
transform 1 0 24380 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_265
timestamp 1704896540
transform 1 0 25484 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_277
timestamp 1704896540
transform 1 0 26588 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_289
timestamp 1704896540
transform 1 0 27692 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94_301
timestamp 1704896540
transform 1 0 28796 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_307
timestamp 1704896540
transform 1 0 29348 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_309
timestamp 1704896540
transform 1 0 29532 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_321
timestamp 1704896540
transform 1 0 30636 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_333
timestamp 1704896540
transform 1 0 31740 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_345
timestamp 1704896540
transform 1 0 32844 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94_357
timestamp 1704896540
transform 1 0 33948 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_363
timestamp 1704896540
transform 1 0 34500 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_365
timestamp 1704896540
transform 1 0 34684 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_377
timestamp 1704896540
transform 1 0 35788 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_389
timestamp 1704896540
transform 1 0 36892 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_94_401
timestamp 1704896540
transform 1 0 37996 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_94_421
timestamp 1704896540
transform 1 0 39836 0 1 53312
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_3
timestamp 1704896540
transform 1 0 1380 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_15
timestamp 1704896540
transform 1 0 2484 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_27
timestamp 1704896540
transform 1 0 3588 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_39
timestamp 1704896540
transform 1 0 4692 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_95_51
timestamp 1704896540
transform 1 0 5796 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_55
timestamp 1704896540
transform 1 0 6164 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_57
timestamp 1704896540
transform 1 0 6348 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_69
timestamp 1704896540
transform 1 0 7452 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_81
timestamp 1704896540
transform 1 0 8556 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_93
timestamp 1704896540
transform 1 0 9660 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_95_105
timestamp 1704896540
transform 1 0 10764 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_111
timestamp 1704896540
transform 1 0 11316 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_113
timestamp 1704896540
transform 1 0 11500 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_125
timestamp 1704896540
transform 1 0 12604 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_137
timestamp 1704896540
transform 1 0 13708 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_95_149
timestamp 1704896540
transform 1 0 14812 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_153
timestamp 1704896540
transform 1 0 15180 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_95_158
timestamp 1704896540
transform 1 0 15640 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_95_166
timestamp 1704896540
transform 1 0 16376 0 -1 54400
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_169
timestamp 1704896540
transform 1 0 16652 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_181
timestamp 1704896540
transform 1 0 17756 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_193
timestamp 1704896540
transform 1 0 18860 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_205
timestamp 1704896540
transform 1 0 19964 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_95_217
timestamp 1704896540
transform 1 0 21068 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_223
timestamp 1704896540
transform 1 0 21620 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_225
timestamp 1704896540
transform 1 0 21804 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_237
timestamp 1704896540
transform 1 0 22908 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_249
timestamp 1704896540
transform 1 0 24012 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_261
timestamp 1704896540
transform 1 0 25116 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_95_273
timestamp 1704896540
transform 1 0 26220 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_279
timestamp 1704896540
transform 1 0 26772 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_281
timestamp 1704896540
transform 1 0 26956 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_95_293
timestamp 1704896540
transform 1 0 28060 0 -1 54400
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_309
timestamp 1704896540
transform 1 0 29532 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_321
timestamp 1704896540
transform 1 0 30636 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_95_333
timestamp 1704896540
transform 1 0 31740 0 -1 54400
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_337
timestamp 1704896540
transform 1 0 32108 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_349
timestamp 1704896540
transform 1 0 33212 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_361
timestamp 1704896540
transform 1 0 34316 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_373
timestamp 1704896540
transform 1 0 35420 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_95_385
timestamp 1704896540
transform 1 0 36524 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_391
timestamp 1704896540
transform 1 0 37076 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_393
timestamp 1704896540
transform 1 0 37260 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_405
timestamp 1704896540
transform 1 0 38364 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_417
timestamp 1704896540
transform 1 0 39468 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_3
timestamp 1704896540
transform 1 0 1380 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_15
timestamp 1704896540
transform 1 0 2484 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_27
timestamp 1704896540
transform 1 0 3588 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_96_49
timestamp 1704896540
transform 1 0 5612 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_96_57
timestamp 1704896540
transform 1 0 6348 0 1 54400
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_67
timestamp 1704896540
transform 1 0 7268 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_96_79
timestamp 1704896540
transform 1 0 8372 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_83
timestamp 1704896540
transform 1 0 8740 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_85
timestamp 1704896540
transform 1 0 8924 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_97
timestamp 1704896540
transform 1 0 10028 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_109
timestamp 1704896540
transform 1 0 11132 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_121
timestamp 1704896540
transform 1 0 12236 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_96_133
timestamp 1704896540
transform 1 0 13340 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_139
timestamp 1704896540
transform 1 0 13892 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_141
timestamp 1704896540
transform 1 0 14076 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_96_153
timestamp 1704896540
transform 1 0 15180 0 1 54400
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_166
timestamp 1704896540
transform 1 0 16376 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_178
timestamp 1704896540
transform 1 0 17480 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_96_190
timestamp 1704896540
transform 1 0 18584 0 1 54400
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_197
timestamp 1704896540
transform 1 0 19228 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_209
timestamp 1704896540
transform 1 0 20332 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_221
timestamp 1704896540
transform 1 0 21436 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_233
timestamp 1704896540
transform 1 0 22540 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_96_245
timestamp 1704896540
transform 1 0 23644 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_251
timestamp 1704896540
transform 1 0 24196 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_253
timestamp 1704896540
transform 1 0 24380 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_265
timestamp 1704896540
transform 1 0 25484 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_277
timestamp 1704896540
transform 1 0 26588 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_289
timestamp 1704896540
transform 1 0 27692 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_96_301
timestamp 1704896540
transform 1 0 28796 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_307
timestamp 1704896540
transform 1 0 29348 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_309
timestamp 1704896540
transform 1 0 29532 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_321
timestamp 1704896540
transform 1 0 30636 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_333
timestamp 1704896540
transform 1 0 31740 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_96_345
timestamp 1704896540
transform 1 0 32844 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_96_353
timestamp 1704896540
transform 1 0 33580 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_96_362
timestamp 1704896540
transform 1 0 34408 0 1 54400
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_365
timestamp 1704896540
transform 1 0 34684 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_377
timestamp 1704896540
transform 1 0 35788 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_389
timestamp 1704896540
transform 1 0 36892 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_401
timestamp 1704896540
transform 1 0 37996 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_96_413
timestamp 1704896540
transform 1 0 39100 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_419
timestamp 1704896540
transform 1 0 39652 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_96_421
timestamp 1704896540
transform 1 0 39836 0 1 54400
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_3
timestamp 1704896540
transform 1 0 1380 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_15
timestamp 1704896540
transform 1 0 2484 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_97_27
timestamp 1704896540
transform 1 0 3588 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_97_52
timestamp 1704896540
transform 1 0 5888 0 -1 55488
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_57
timestamp 1704896540
transform 1 0 6348 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_69
timestamp 1704896540
transform 1 0 7452 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_81
timestamp 1704896540
transform 1 0 8556 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_93
timestamp 1704896540
transform 1 0 9660 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_97_105
timestamp 1704896540
transform 1 0 10764 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_111
timestamp 1704896540
transform 1 0 11316 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_113
timestamp 1704896540
transform 1 0 11500 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_125
timestamp 1704896540
transform 1 0 12604 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_137
timestamp 1704896540
transform 1 0 13708 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_149
timestamp 1704896540
transform 1 0 14812 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_97_161
timestamp 1704896540
transform 1 0 15916 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_167
timestamp 1704896540
transform 1 0 16468 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_169
timestamp 1704896540
transform 1 0 16652 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_181
timestamp 1704896540
transform 1 0 17756 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_193
timestamp 1704896540
transform 1 0 18860 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_205
timestamp 1704896540
transform 1 0 19964 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_97_217
timestamp 1704896540
transform 1 0 21068 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_223
timestamp 1704896540
transform 1 0 21620 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_225
timestamp 1704896540
transform 1 0 21804 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_237
timestamp 1704896540
transform 1 0 22908 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_249
timestamp 1704896540
transform 1 0 24012 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_261
timestamp 1704896540
transform 1 0 25116 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_97_273
timestamp 1704896540
transform 1 0 26220 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_279
timestamp 1704896540
transform 1 0 26772 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_281
timestamp 1704896540
transform 1 0 26956 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_293
timestamp 1704896540
transform 1 0 28060 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_305
timestamp 1704896540
transform 1 0 29164 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_317
timestamp 1704896540
transform 1 0 30268 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_97_329
timestamp 1704896540
transform 1 0 31372 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_335
timestamp 1704896540
transform 1 0 31924 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_337
timestamp 1704896540
transform 1 0 32108 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_349
timestamp 1704896540
transform 1 0 33212 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_361
timestamp 1704896540
transform 1 0 34316 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_373
timestamp 1704896540
transform 1 0 35420 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_97_385
timestamp 1704896540
transform 1 0 36524 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_391
timestamp 1704896540
transform 1 0 37076 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_393
timestamp 1704896540
transform 1 0 37260 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_405
timestamp 1704896540
transform 1 0 38364 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_417
timestamp 1704896540
transform 1 0 39468 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_3
timestamp 1704896540
transform 1 0 1380 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_15
timestamp 1704896540
transform 1 0 2484 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_27
timestamp 1704896540
transform 1 0 3588 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_29
timestamp 1704896540
transform 1 0 3772 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_41
timestamp 1704896540
transform 1 0 4876 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_53
timestamp 1704896540
transform 1 0 5980 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_65
timestamp 1704896540
transform 1 0 7084 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_98_77
timestamp 1704896540
transform 1 0 8188 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_83
timestamp 1704896540
transform 1 0 8740 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_98_85
timestamp 1704896540
transform 1 0 8924 0 1 55488
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_99
timestamp 1704896540
transform 1 0 10212 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_111
timestamp 1704896540
transform 1 0 11316 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_123
timestamp 1704896540
transform 1 0 12420 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_98_135
timestamp 1704896540
transform 1 0 13524 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_139
timestamp 1704896540
transform 1 0 13892 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_141
timestamp 1704896540
transform 1 0 14076 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_98_153
timestamp 1704896540
transform 1 0 15180 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_159
timestamp 1704896540
transform 1 0 15732 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_169
timestamp 1704896540
transform 1 0 16652 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_181
timestamp 1704896540
transform 1 0 17756 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_98_193
timestamp 1704896540
transform 1 0 18860 0 1 55488
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_197
timestamp 1704896540
transform 1 0 19228 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_209
timestamp 1704896540
transform 1 0 20332 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_221
timestamp 1704896540
transform 1 0 21436 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_233
timestamp 1704896540
transform 1 0 22540 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_98_245
timestamp 1704896540
transform 1 0 23644 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_251
timestamp 1704896540
transform 1 0 24196 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_253
timestamp 1704896540
transform 1 0 24380 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_265
timestamp 1704896540
transform 1 0 25484 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_277
timestamp 1704896540
transform 1 0 26588 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_289
timestamp 1704896540
transform 1 0 27692 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_98_301
timestamp 1704896540
transform 1 0 28796 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_307
timestamp 1704896540
transform 1 0 29348 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_309
timestamp 1704896540
transform 1 0 29532 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_321
timestamp 1704896540
transform 1 0 30636 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_333
timestamp 1704896540
transform 1 0 31740 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_345
timestamp 1704896540
transform 1 0 32844 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_98_357
timestamp 1704896540
transform 1 0 33948 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_363
timestamp 1704896540
transform 1 0 34500 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_365
timestamp 1704896540
transform 1 0 34684 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_377
timestamp 1704896540
transform 1 0 35788 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_389
timestamp 1704896540
transform 1 0 36892 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_401
timestamp 1704896540
transform 1 0 37996 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_98_413
timestamp 1704896540
transform 1 0 39100 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_419
timestamp 1704896540
transform 1 0 39652 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_98_421
timestamp 1704896540
transform 1 0 39836 0 1 55488
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_3
timestamp 1704896540
transform 1 0 1380 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_15
timestamp 1704896540
transform 1 0 2484 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_27
timestamp 1704896540
transform 1 0 3588 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_39
timestamp 1704896540
transform 1 0 4692 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_99_51
timestamp 1704896540
transform 1 0 5796 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_55
timestamp 1704896540
transform 1 0 6164 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_57
timestamp 1704896540
transform 1 0 6348 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_69
timestamp 1704896540
transform 1 0 7452 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_81
timestamp 1704896540
transform 1 0 8556 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_93
timestamp 1704896540
transform 1 0 9660 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_99_105
timestamp 1704896540
transform 1 0 10764 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_111
timestamp 1704896540
transform 1 0 11316 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_113
timestamp 1704896540
transform 1 0 11500 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_125
timestamp 1704896540
transform 1 0 12604 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_137
timestamp 1704896540
transform 1 0 13708 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_149
timestamp 1704896540
transform 1 0 14812 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_99_161
timestamp 1704896540
transform 1 0 15916 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_167
timestamp 1704896540
transform 1 0 16468 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_169
timestamp 1704896540
transform 1 0 16652 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_181
timestamp 1704896540
transform 1 0 17756 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_193
timestamp 1704896540
transform 1 0 18860 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_205
timestamp 1704896540
transform 1 0 19964 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_99_217
timestamp 1704896540
transform 1 0 21068 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_223
timestamp 1704896540
transform 1 0 21620 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_225
timestamp 1704896540
transform 1 0 21804 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_237
timestamp 1704896540
transform 1 0 22908 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_249
timestamp 1704896540
transform 1 0 24012 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_261
timestamp 1704896540
transform 1 0 25116 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_99_273
timestamp 1704896540
transform 1 0 26220 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_279
timestamp 1704896540
transform 1 0 26772 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_281
timestamp 1704896540
transform 1 0 26956 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_293
timestamp 1704896540
transform 1 0 28060 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_305
timestamp 1704896540
transform 1 0 29164 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_317
timestamp 1704896540
transform 1 0 30268 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_99_329
timestamp 1704896540
transform 1 0 31372 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_335
timestamp 1704896540
transform 1 0 31924 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_337
timestamp 1704896540
transform 1 0 32108 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_349
timestamp 1704896540
transform 1 0 33212 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_361
timestamp 1704896540
transform 1 0 34316 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_373
timestamp 1704896540
transform 1 0 35420 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_99_385
timestamp 1704896540
transform 1 0 36524 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_391
timestamp 1704896540
transform 1 0 37076 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_393
timestamp 1704896540
transform 1 0 37260 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_405
timestamp 1704896540
transform 1 0 38364 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_417
timestamp 1704896540
transform 1 0 39468 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_3
timestamp 1704896540
transform 1 0 1380 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_15
timestamp 1704896540
transform 1 0 2484 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_27
timestamp 1704896540
transform 1 0 3588 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_29
timestamp 1704896540
transform 1 0 3772 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_41
timestamp 1704896540
transform 1 0 4876 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_53
timestamp 1704896540
transform 1 0 5980 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_65
timestamp 1704896540
transform 1 0 7084 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_100_77
timestamp 1704896540
transform 1 0 8188 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_83
timestamp 1704896540
transform 1 0 8740 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_85
timestamp 1704896540
transform 1 0 8924 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_114
timestamp 1704896540
transform 1 0 11592 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_126
timestamp 1704896540
transform 1 0 12696 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_100_138
timestamp 1704896540
transform 1 0 13800 0 1 56576
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_141
timestamp 1704896540
transform 1 0 14076 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_153
timestamp 1704896540
transform 1 0 15180 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_165
timestamp 1704896540
transform 1 0 16284 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_177
timestamp 1704896540
transform 1 0 17388 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_100_189
timestamp 1704896540
transform 1 0 18492 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_195
timestamp 1704896540
transform 1 0 19044 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_197
timestamp 1704896540
transform 1 0 19228 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_209
timestamp 1704896540
transform 1 0 20332 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_221
timestamp 1704896540
transform 1 0 21436 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_233
timestamp 1704896540
transform 1 0 22540 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_100_245
timestamp 1704896540
transform 1 0 23644 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_251
timestamp 1704896540
transform 1 0 24196 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_253
timestamp 1704896540
transform 1 0 24380 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_100_265
timestamp 1704896540
transform 1 0 25484 0 1 56576
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_280
timestamp 1704896540
transform 1 0 26864 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_292
timestamp 1704896540
transform 1 0 27968 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_100_304
timestamp 1704896540
transform 1 0 29072 0 1 56576
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_309
timestamp 1704896540
transform 1 0 29532 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_321
timestamp 1704896540
transform 1 0 30636 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_333
timestamp 1704896540
transform 1 0 31740 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_345
timestamp 1704896540
transform 1 0 32844 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_100_357
timestamp 1704896540
transform 1 0 33948 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_363
timestamp 1704896540
transform 1 0 34500 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_365
timestamp 1704896540
transform 1 0 34684 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_377
timestamp 1704896540
transform 1 0 35788 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_389
timestamp 1704896540
transform 1 0 36892 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_401
timestamp 1704896540
transform 1 0 37996 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_100_413
timestamp 1704896540
transform 1 0 39100 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_419
timestamp 1704896540
transform 1 0 39652 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_100_421
timestamp 1704896540
transform 1 0 39836 0 1 56576
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_3
timestamp 1704896540
transform 1 0 1380 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_15
timestamp 1704896540
transform 1 0 2484 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_27
timestamp 1704896540
transform 1 0 3588 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_39
timestamp 1704896540
transform 1 0 4692 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_101_51
timestamp 1704896540
transform 1 0 5796 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_55
timestamp 1704896540
transform 1 0 6164 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_57
timestamp 1704896540
transform 1 0 6348 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_69
timestamp 1704896540
transform 1 0 7452 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_81
timestamp 1704896540
transform 1 0 8556 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_93
timestamp 1704896540
transform 1 0 9660 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_101_105
timestamp 1704896540
transform 1 0 10764 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_111
timestamp 1704896540
transform 1 0 11316 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_113
timestamp 1704896540
transform 1 0 11500 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_125
timestamp 1704896540
transform 1 0 12604 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_137
timestamp 1704896540
transform 1 0 13708 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_149
timestamp 1704896540
transform 1 0 14812 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_101_161
timestamp 1704896540
transform 1 0 15916 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_167
timestamp 1704896540
transform 1 0 16468 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_176
timestamp 1704896540
transform 1 0 17296 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_188
timestamp 1704896540
transform 1 0 18400 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_200
timestamp 1704896540
transform 1 0 19504 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_212
timestamp 1704896540
transform 1 0 20608 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_225
timestamp 1704896540
transform 1 0 21804 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_237
timestamp 1704896540
transform 1 0 22908 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_249
timestamp 1704896540
transform 1 0 24012 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_261
timestamp 1704896540
transform 1 0 25116 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_101_273
timestamp 1704896540
transform 1 0 26220 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_279
timestamp 1704896540
transform 1 0 26772 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_281
timestamp 1704896540
transform 1 0 26956 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_293
timestamp 1704896540
transform 1 0 28060 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_305
timestamp 1704896540
transform 1 0 29164 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_317
timestamp 1704896540
transform 1 0 30268 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_101_329
timestamp 1704896540
transform 1 0 31372 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_335
timestamp 1704896540
transform 1 0 31924 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_337
timestamp 1704896540
transform 1 0 32108 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_349
timestamp 1704896540
transform 1 0 33212 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_361
timestamp 1704896540
transform 1 0 34316 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_373
timestamp 1704896540
transform 1 0 35420 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_101_385
timestamp 1704896540
transform 1 0 36524 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_391
timestamp 1704896540
transform 1 0 37076 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_393
timestamp 1704896540
transform 1 0 37260 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_101_405
timestamp 1704896540
transform 1 0 38364 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_411
timestamp 1704896540
transform 1 0 38916 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_3
timestamp 1704896540
transform 1 0 1380 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_15
timestamp 1704896540
transform 1 0 2484 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_102_27
timestamp 1704896540
transform 1 0 3588 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_29
timestamp 1704896540
transform 1 0 3772 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_41
timestamp 1704896540
transform 1 0 4876 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_53
timestamp 1704896540
transform 1 0 5980 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_65
timestamp 1704896540
transform 1 0 7084 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_102_77
timestamp 1704896540
transform 1 0 8188 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_102_83
timestamp 1704896540
transform 1 0 8740 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_85
timestamp 1704896540
transform 1 0 8924 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_97
timestamp 1704896540
transform 1 0 10028 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_109
timestamp 1704896540
transform 1 0 11132 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_121
timestamp 1704896540
transform 1 0 12236 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_102_133
timestamp 1704896540
transform 1 0 13340 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_102_139
timestamp 1704896540
transform 1 0 13892 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_141
timestamp 1704896540
transform 1 0 14076 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_153
timestamp 1704896540
transform 1 0 15180 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_165
timestamp 1704896540
transform 1 0 16284 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_177
timestamp 1704896540
transform 1 0 17388 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_102_189
timestamp 1704896540
transform 1 0 18492 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_102_195
timestamp 1704896540
transform 1 0 19044 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_102_197
timestamp 1704896540
transform 1 0 19228 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_102_203
timestamp 1704896540
transform 1 0 19780 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_218
timestamp 1704896540
transform 1 0 21160 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_230
timestamp 1704896540
transform 1 0 22264 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_102_242
timestamp 1704896540
transform 1 0 23368 0 1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_102_250
timestamp 1704896540
transform 1 0 24104 0 1 57664
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_257
timestamp 1704896540
transform 1 0 24748 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_102_269
timestamp 1704896540
transform 1 0 25852 0 1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_102_277
timestamp 1704896540
transform 1 0 26588 0 1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_102_281
timestamp 1704896540
transform 1 0 26956 0 1 57664
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_291
timestamp 1704896540
transform 1 0 27876 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_102_303
timestamp 1704896540
transform 1 0 28980 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_102_307
timestamp 1704896540
transform 1 0 29348 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_309
timestamp 1704896540
transform 1 0 29532 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_321
timestamp 1704896540
transform 1 0 30636 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_333
timestamp 1704896540
transform 1 0 31740 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_345
timestamp 1704896540
transform 1 0 32844 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_102_357
timestamp 1704896540
transform 1 0 33948 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_102_363
timestamp 1704896540
transform 1 0 34500 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_365
timestamp 1704896540
transform 1 0 34684 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_377
timestamp 1704896540
transform 1 0 35788 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_389
timestamp 1704896540
transform 1 0 36892 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_401
timestamp 1704896540
transform 1 0 37996 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_102_413
timestamp 1704896540
transform 1 0 39100 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_102_419
timestamp 1704896540
transform 1 0 39652 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_102_421
timestamp 1704896540
transform 1 0 39836 0 1 57664
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_19
timestamp 1704896540
transform 1 0 2852 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_31
timestamp 1704896540
transform 1 0 3956 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_43
timestamp 1704896540
transform 1 0 5060 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_103_55
timestamp 1704896540
transform 1 0 6164 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_57
timestamp 1704896540
transform 1 0 6348 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_69
timestamp 1704896540
transform 1 0 7452 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_81
timestamp 1704896540
transform 1 0 8556 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_93
timestamp 1704896540
transform 1 0 9660 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_103_105
timestamp 1704896540
transform 1 0 10764 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_103_111
timestamp 1704896540
transform 1 0 11316 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_113
timestamp 1704896540
transform 1 0 11500 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_103_125
timestamp 1704896540
transform 1 0 12604 0 -1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_103_133
timestamp 1704896540
transform 1 0 13340 0 -1 58752
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_149
timestamp 1704896540
transform 1 0 14812 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_103_161
timestamp 1704896540
transform 1 0 15916 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_103_167
timestamp 1704896540
transform 1 0 16468 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_169
timestamp 1704896540
transform 1 0 16652 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_181
timestamp 1704896540
transform 1 0 17756 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_193
timestamp 1704896540
transform 1 0 18860 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_205
timestamp 1704896540
transform 1 0 19964 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_103_217
timestamp 1704896540
transform 1 0 21068 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_103_223
timestamp 1704896540
transform 1 0 21620 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_225
timestamp 1704896540
transform 1 0 21804 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_237
timestamp 1704896540
transform 1 0 22908 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_249
timestamp 1704896540
transform 1 0 24012 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_261
timestamp 1704896540
transform 1 0 25116 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_103_273
timestamp 1704896540
transform 1 0 26220 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_103_279
timestamp 1704896540
transform 1 0 26772 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_281
timestamp 1704896540
transform 1 0 26956 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_293
timestamp 1704896540
transform 1 0 28060 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_305
timestamp 1704896540
transform 1 0 29164 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_317
timestamp 1704896540
transform 1 0 30268 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_103_329
timestamp 1704896540
transform 1 0 31372 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_103_335
timestamp 1704896540
transform 1 0 31924 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_337
timestamp 1704896540
transform 1 0 32108 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_349
timestamp 1704896540
transform 1 0 33212 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_361
timestamp 1704896540
transform 1 0 34316 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_373
timestamp 1704896540
transform 1 0 35420 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_103_385
timestamp 1704896540
transform 1 0 36524 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_103_391
timestamp 1704896540
transform 1 0 37076 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_103_393
timestamp 1704896540
transform 1 0 37260 0 -1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_103_423
timestamp 1704896540
transform 1 0 40020 0 -1 58752
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_3
timestamp 1704896540
transform 1 0 1380 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_15
timestamp 1704896540
transform 1 0 2484 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_104_27
timestamp 1704896540
transform 1 0 3588 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_104_29
timestamp 1704896540
transform 1 0 3772 0 1 58752
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_40
timestamp 1704896540
transform 1 0 4784 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_104_52
timestamp 1704896540
transform 1 0 5888 0 1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_104_60
timestamp 1704896540
transform 1 0 6624 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_68
timestamp 1704896540
transform 1 0 7360 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_104_80
timestamp 1704896540
transform 1 0 8464 0 1 58752
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_85
timestamp 1704896540
transform 1 0 8924 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_97
timestamp 1704896540
transform 1 0 10028 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_109
timestamp 1704896540
transform 1 0 11132 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_121
timestamp 1704896540
transform 1 0 12236 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_104_133
timestamp 1704896540
transform 1 0 13340 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_104_139
timestamp 1704896540
transform 1 0 13892 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_141
timestamp 1704896540
transform 1 0 14076 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_153
timestamp 1704896540
transform 1 0 15180 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_165
timestamp 1704896540
transform 1 0 16284 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_177
timestamp 1704896540
transform 1 0 17388 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_104_189
timestamp 1704896540
transform 1 0 18492 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_104_195
timestamp 1704896540
transform 1 0 19044 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_197
timestamp 1704896540
transform 1 0 19228 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_209
timestamp 1704896540
transform 1 0 20332 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_221
timestamp 1704896540
transform 1 0 21436 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_104_233
timestamp 1704896540
transform 1 0 22540 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_104_246
timestamp 1704896540
transform 1 0 23736 0 1 58752
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_253
timestamp 1704896540
transform 1 0 24380 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_265
timestamp 1704896540
transform 1 0 25484 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_277
timestamp 1704896540
transform 1 0 26588 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_289
timestamp 1704896540
transform 1 0 27692 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_104_301
timestamp 1704896540
transform 1 0 28796 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_104_307
timestamp 1704896540
transform 1 0 29348 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_104_309
timestamp 1704896540
transform 1 0 29532 0 1 58752
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_326
timestamp 1704896540
transform 1 0 31096 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_338
timestamp 1704896540
transform 1 0 32200 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_350
timestamp 1704896540
transform 1 0 33304 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_104_362
timestamp 1704896540
transform 1 0 34408 0 1 58752
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_365
timestamp 1704896540
transform 1 0 34684 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_377
timestamp 1704896540
transform 1 0 35788 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_389
timestamp 1704896540
transform 1 0 36892 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_104_401
timestamp 1704896540
transform 1 0 37996 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_407
timestamp 1704896540
transform 1 0 38548 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_104_419
timestamp 1704896540
transform 1 0 39652 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_104_421
timestamp 1704896540
transform 1 0 39836 0 1 58752
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_3
timestamp 1704896540
transform 1 0 1380 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_15
timestamp 1704896540
transform 1 0 2484 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_27
timestamp 1704896540
transform 1 0 3588 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_39
timestamp 1704896540
transform 1 0 4692 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_105_51
timestamp 1704896540
transform 1 0 5796 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_105_55
timestamp 1704896540
transform 1 0 6164 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_57
timestamp 1704896540
transform 1 0 6348 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_69
timestamp 1704896540
transform 1 0 7452 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_81
timestamp 1704896540
transform 1 0 8556 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_93
timestamp 1704896540
transform 1 0 9660 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_105_105
timestamp 1704896540
transform 1 0 10764 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_105_111
timestamp 1704896540
transform 1 0 11316 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_113
timestamp 1704896540
transform 1 0 11500 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_125
timestamp 1704896540
transform 1 0 12604 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_137
timestamp 1704896540
transform 1 0 13708 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_149
timestamp 1704896540
transform 1 0 14812 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_105_161
timestamp 1704896540
transform 1 0 15916 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_105_167
timestamp 1704896540
transform 1 0 16468 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_169
timestamp 1704896540
transform 1 0 16652 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_181
timestamp 1704896540
transform 1 0 17756 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_105_193
timestamp 1704896540
transform 1 0 18860 0 -1 59840
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_199
timestamp 1704896540
transform 1 0 19412 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_211
timestamp 1704896540
transform 1 0 20516 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_105_223
timestamp 1704896540
transform 1 0 21620 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_225
timestamp 1704896540
transform 1 0 21804 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_237
timestamp 1704896540
transform 1 0 22908 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_249
timestamp 1704896540
transform 1 0 24012 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_261
timestamp 1704896540
transform 1 0 25116 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_105_273
timestamp 1704896540
transform 1 0 26220 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_105_279
timestamp 1704896540
transform 1 0 26772 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_281
timestamp 1704896540
transform 1 0 26956 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_293
timestamp 1704896540
transform 1 0 28060 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_305
timestamp 1704896540
transform 1 0 29164 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_317
timestamp 1704896540
transform 1 0 30268 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_105_329
timestamp 1704896540
transform 1 0 31372 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_105_335
timestamp 1704896540
transform 1 0 31924 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_337
timestamp 1704896540
transform 1 0 32108 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_349
timestamp 1704896540
transform 1 0 33212 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_361
timestamp 1704896540
transform 1 0 34316 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_373
timestamp 1704896540
transform 1 0 35420 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_105_385
timestamp 1704896540
transform 1 0 36524 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_105_391
timestamp 1704896540
transform 1 0 37076 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_393
timestamp 1704896540
transform 1 0 37260 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_405
timestamp 1704896540
transform 1 0 38364 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_3
timestamp 1704896540
transform 1 0 1380 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_15
timestamp 1704896540
transform 1 0 2484 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_106_27
timestamp 1704896540
transform 1 0 3588 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_29
timestamp 1704896540
transform 1 0 3772 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_41
timestamp 1704896540
transform 1 0 4876 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_53
timestamp 1704896540
transform 1 0 5980 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_65
timestamp 1704896540
transform 1 0 7084 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_106_77
timestamp 1704896540
transform 1 0 8188 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_106_83
timestamp 1704896540
transform 1 0 8740 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_85
timestamp 1704896540
transform 1 0 8924 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_97
timestamp 1704896540
transform 1 0 10028 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_109
timestamp 1704896540
transform 1 0 11132 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_121
timestamp 1704896540
transform 1 0 12236 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_106_133
timestamp 1704896540
transform 1 0 13340 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_106_139
timestamp 1704896540
transform 1 0 13892 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_141
timestamp 1704896540
transform 1 0 14076 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_153
timestamp 1704896540
transform 1 0 15180 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_165
timestamp 1704896540
transform 1 0 16284 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_177
timestamp 1704896540
transform 1 0 17388 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_106_189
timestamp 1704896540
transform 1 0 18492 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_106_195
timestamp 1704896540
transform 1 0 19044 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_204
timestamp 1704896540
transform 1 0 19872 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_106_216
timestamp 1704896540
transform 1 0 20976 0 1 59840
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_231
timestamp 1704896540
transform 1 0 22356 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_106_243
timestamp 1704896540
transform 1 0 23460 0 1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_106_251
timestamp 1704896540
transform 1 0 24196 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_253
timestamp 1704896540
transform 1 0 24380 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_265
timestamp 1704896540
transform 1 0 25484 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_277
timestamp 1704896540
transform 1 0 26588 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_289
timestamp 1704896540
transform 1 0 27692 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_106_301
timestamp 1704896540
transform 1 0 28796 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_106_307
timestamp 1704896540
transform 1 0 29348 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_318
timestamp 1704896540
transform 1 0 30360 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_330
timestamp 1704896540
transform 1 0 31464 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_369
timestamp 1704896540
transform 1 0 35052 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_381
timestamp 1704896540
transform 1 0 36156 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_393
timestamp 1704896540
transform 1 0 37260 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_405
timestamp 1704896540
transform 1 0 38364 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_106_417
timestamp 1704896540
transform 1 0 39468 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_106_421
timestamp 1704896540
transform 1 0 39836 0 1 59840
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_3
timestamp 1704896540
transform 1 0 1380 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_15
timestamp 1704896540
transform 1 0 2484 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_27
timestamp 1704896540
transform 1 0 3588 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_39
timestamp 1704896540
transform 1 0 4692 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_107_51
timestamp 1704896540
transform 1 0 5796 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_107_55
timestamp 1704896540
transform 1 0 6164 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_57
timestamp 1704896540
transform 1 0 6348 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_107_69
timestamp 1704896540
transform 1 0 7452 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_107_73
timestamp 1704896540
transform 1 0 7820 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_88
timestamp 1704896540
transform 1 0 9200 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_100
timestamp 1704896540
transform 1 0 10304 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_113
timestamp 1704896540
transform 1 0 11500 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_125
timestamp 1704896540
transform 1 0 12604 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_137
timestamp 1704896540
transform 1 0 13708 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_149
timestamp 1704896540
transform 1 0 14812 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_107_161
timestamp 1704896540
transform 1 0 15916 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_107_167
timestamp 1704896540
transform 1 0 16468 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_169
timestamp 1704896540
transform 1 0 16652 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_181
timestamp 1704896540
transform 1 0 17756 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_107_193
timestamp 1704896540
transform 1 0 18860 0 -1 60928
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_199
timestamp 1704896540
transform 1 0 19412 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_211
timestamp 1704896540
transform 1 0 20516 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_107_223
timestamp 1704896540
transform 1 0 21620 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_225
timestamp 1704896540
transform 1 0 21804 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_237
timestamp 1704896540
transform 1 0 22908 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_249
timestamp 1704896540
transform 1 0 24012 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_261
timestamp 1704896540
transform 1 0 25116 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_107_273
timestamp 1704896540
transform 1 0 26220 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_107_279
timestamp 1704896540
transform 1 0 26772 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_281
timestamp 1704896540
transform 1 0 26956 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_107_293
timestamp 1704896540
transform 1 0 28060 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_107_301
timestamp 1704896540
transform 1 0 28796 0 -1 60928
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_312
timestamp 1704896540
transform 1 0 29808 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_324
timestamp 1704896540
transform 1 0 30912 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_337
timestamp 1704896540
transform 1 0 32108 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_349
timestamp 1704896540
transform 1 0 33212 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_361
timestamp 1704896540
transform 1 0 34316 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_373
timestamp 1704896540
transform 1 0 35420 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_107_385
timestamp 1704896540
transform 1 0 36524 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_107_391
timestamp 1704896540
transform 1 0 37076 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_107_393
timestamp 1704896540
transform 1 0 37260 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_107_401
timestamp 1704896540
transform 1 0 37996 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_107_406
timestamp 1704896540
transform 1 0 38456 0 -1 60928
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_414
timestamp 1704896540
transform 1 0 39192 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_107_426
timestamp 1704896540
transform 1 0 40296 0 -1 60928
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_16
timestamp 1704896540
transform 1 0 2576 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_108_37
timestamp 1704896540
transform 1 0 4508 0 1 60928
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_41
timestamp 1704896540
transform 1 0 4876 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_53
timestamp 1704896540
transform 1 0 5980 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_65
timestamp 1704896540
transform 1 0 7084 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_108_77
timestamp 1704896540
transform 1 0 8188 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_108_83
timestamp 1704896540
transform 1 0 8740 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_94
timestamp 1704896540
transform 1 0 9752 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_106
timestamp 1704896540
transform 1 0 10856 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_118
timestamp 1704896540
transform 1 0 11960 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_108_130
timestamp 1704896540
transform 1 0 13064 0 1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_108_138
timestamp 1704896540
transform 1 0 13800 0 1 60928
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_141
timestamp 1704896540
transform 1 0 14076 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_153
timestamp 1704896540
transform 1 0 15180 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_165
timestamp 1704896540
transform 1 0 16284 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_177
timestamp 1704896540
transform 1 0 17388 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_108_189
timestamp 1704896540
transform 1 0 18492 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_108_195
timestamp 1704896540
transform 1 0 19044 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_197
timestamp 1704896540
transform 1 0 19228 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_209
timestamp 1704896540
transform 1 0 20332 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_221
timestamp 1704896540
transform 1 0 21436 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_233
timestamp 1704896540
transform 1 0 22540 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_108_245
timestamp 1704896540
transform 1 0 23644 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_108_251
timestamp 1704896540
transform 1 0 24196 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_253
timestamp 1704896540
transform 1 0 24380 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_265
timestamp 1704896540
transform 1 0 25484 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_277
timestamp 1704896540
transform 1 0 26588 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_289
timestamp 1704896540
transform 1 0 27692 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_108_301
timestamp 1704896540
transform 1 0 28796 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_108_307
timestamp 1704896540
transform 1 0 29348 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_309
timestamp 1704896540
transform 1 0 29532 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_321
timestamp 1704896540
transform 1 0 30636 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_333
timestamp 1704896540
transform 1 0 31740 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_345
timestamp 1704896540
transform 1 0 32844 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_108_357
timestamp 1704896540
transform 1 0 33948 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_108_363
timestamp 1704896540
transform 1 0 34500 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_365
timestamp 1704896540
transform 1 0 34684 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_377
timestamp 1704896540
transform 1 0 35788 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_389
timestamp 1704896540
transform 1 0 36892 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_401
timestamp 1704896540
transform 1 0 37996 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_108_413
timestamp 1704896540
transform 1 0 39100 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_108_419
timestamp 1704896540
transform 1 0 39652 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_108_421
timestamp 1704896540
transform 1 0 39836 0 1 60928
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_3
timestamp 1704896540
transform 1 0 1380 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_15
timestamp 1704896540
transform 1 0 2484 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_27
timestamp 1704896540
transform 1 0 3588 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_39
timestamp 1704896540
transform 1 0 4692 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_109_51
timestamp 1704896540
transform 1 0 5796 0 -1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_109_55
timestamp 1704896540
transform 1 0 6164 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_57
timestamp 1704896540
transform 1 0 6348 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_69
timestamp 1704896540
transform 1 0 7452 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_81
timestamp 1704896540
transform 1 0 8556 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_93
timestamp 1704896540
transform 1 0 9660 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_109_105
timestamp 1704896540
transform 1 0 10764 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_109_111
timestamp 1704896540
transform 1 0 11316 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_113
timestamp 1704896540
transform 1 0 11500 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_109_125
timestamp 1704896540
transform 1 0 12604 0 -1 62016
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_138
timestamp 1704896540
transform 1 0 13800 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_150
timestamp 1704896540
transform 1 0 14904 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_109_162
timestamp 1704896540
transform 1 0 16008 0 -1 62016
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_169
timestamp 1704896540
transform 1 0 16652 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_183
timestamp 1704896540
transform 1 0 17940 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_195
timestamp 1704896540
transform 1 0 19044 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_207
timestamp 1704896540
transform 1 0 20148 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_109_219
timestamp 1704896540
transform 1 0 21252 0 -1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_109_223
timestamp 1704896540
transform 1 0 21620 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_225
timestamp 1704896540
transform 1 0 21804 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_237
timestamp 1704896540
transform 1 0 22908 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_249
timestamp 1704896540
transform 1 0 24012 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_261
timestamp 1704896540
transform 1 0 25116 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_109_273
timestamp 1704896540
transform 1 0 26220 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_109_279
timestamp 1704896540
transform 1 0 26772 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_281
timestamp 1704896540
transform 1 0 26956 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_293
timestamp 1704896540
transform 1 0 28060 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_305
timestamp 1704896540
transform 1 0 29164 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_317
timestamp 1704896540
transform 1 0 30268 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_109_329
timestamp 1704896540
transform 1 0 31372 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_109_335
timestamp 1704896540
transform 1 0 31924 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_337
timestamp 1704896540
transform 1 0 32108 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_349
timestamp 1704896540
transform 1 0 33212 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_361
timestamp 1704896540
transform 1 0 34316 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_373
timestamp 1704896540
transform 1 0 35420 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_109_385
timestamp 1704896540
transform 1 0 36524 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_109_391
timestamp 1704896540
transform 1 0 37076 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_393
timestamp 1704896540
transform 1 0 37260 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_405
timestamp 1704896540
transform 1 0 38364 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_417
timestamp 1704896540
transform 1 0 39468 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_3
timestamp 1704896540
transform 1 0 1380 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_15
timestamp 1704896540
transform 1 0 2484 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_110_27
timestamp 1704896540
transform 1 0 3588 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_29
timestamp 1704896540
transform 1 0 3772 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_41
timestamp 1704896540
transform 1 0 4876 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_53
timestamp 1704896540
transform 1 0 5980 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_110_65
timestamp 1704896540
transform 1 0 7084 0 1 62016
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_71
timestamp 1704896540
transform 1 0 7636 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_110_83
timestamp 1704896540
transform 1 0 8740 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_85
timestamp 1704896540
transform 1 0 8924 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_97
timestamp 1704896540
transform 1 0 10028 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_110_109
timestamp 1704896540
transform 1 0 11132 0 1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_110_134
timestamp 1704896540
transform 1 0 13432 0 1 62016
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_141
timestamp 1704896540
transform 1 0 14076 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_153
timestamp 1704896540
transform 1 0 15180 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_165
timestamp 1704896540
transform 1 0 16284 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_110_177
timestamp 1704896540
transform 1 0 17388 0 1 62016
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_183
timestamp 1704896540
transform 1 0 17940 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_110_195
timestamp 1704896540
transform 1 0 19044 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_110_197
timestamp 1704896540
transform 1 0 19228 0 1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110_205
timestamp 1704896540
transform 1 0 19964 0 1 62016
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_216
timestamp 1704896540
transform 1 0 20976 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_228
timestamp 1704896540
transform 1 0 22080 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_240
timestamp 1704896540
transform 1 0 23184 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_253
timestamp 1704896540
transform 1 0 24380 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_265
timestamp 1704896540
transform 1 0 25484 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_277
timestamp 1704896540
transform 1 0 26588 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_289
timestamp 1704896540
transform 1 0 27692 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_110_301
timestamp 1704896540
transform 1 0 28796 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_110_307
timestamp 1704896540
transform 1 0 29348 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_309
timestamp 1704896540
transform 1 0 29532 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_321
timestamp 1704896540
transform 1 0 30636 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_333
timestamp 1704896540
transform 1 0 31740 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_345
timestamp 1704896540
transform 1 0 32844 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_110_357
timestamp 1704896540
transform 1 0 33948 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_110_363
timestamp 1704896540
transform 1 0 34500 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_378
timestamp 1704896540
transform 1 0 35880 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_390
timestamp 1704896540
transform 1 0 36984 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_402
timestamp 1704896540
transform 1 0 38088 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_110_414
timestamp 1704896540
transform 1 0 39192 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_110_421
timestamp 1704896540
transform 1 0 39836 0 1 62016
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_3
timestamp 1704896540
transform 1 0 1380 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_15
timestamp 1704896540
transform 1 0 2484 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_27
timestamp 1704896540
transform 1 0 3588 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_39
timestamp 1704896540
transform 1 0 4692 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_111_51
timestamp 1704896540
transform 1 0 5796 0 -1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111_55
timestamp 1704896540
transform 1 0 6164 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_57
timestamp 1704896540
transform 1 0 6348 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_111_69
timestamp 1704896540
transform 1 0 7452 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111_75
timestamp 1704896540
transform 1 0 8004 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_81
timestamp 1704896540
transform 1 0 8556 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_93
timestamp 1704896540
transform 1 0 9660 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_111_105
timestamp 1704896540
transform 1 0 10764 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111_111
timestamp 1704896540
transform 1 0 11316 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_113
timestamp 1704896540
transform 1 0 11500 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_125
timestamp 1704896540
transform 1 0 12604 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_137
timestamp 1704896540
transform 1 0 13708 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_149
timestamp 1704896540
transform 1 0 14812 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_111_161
timestamp 1704896540
transform 1 0 15916 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111_167
timestamp 1704896540
transform 1 0 16468 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_169
timestamp 1704896540
transform 1 0 16652 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_190
timestamp 1704896540
transform 1 0 18584 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_202
timestamp 1704896540
transform 1 0 19688 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_111_214
timestamp 1704896540
transform 1 0 20792 0 -1 63104
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_111_222
timestamp 1704896540
transform 1 0 21528 0 -1 63104
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_225
timestamp 1704896540
transform 1 0 21804 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_237
timestamp 1704896540
transform 1 0 22908 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_249
timestamp 1704896540
transform 1 0 24012 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_261
timestamp 1704896540
transform 1 0 25116 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_111_273
timestamp 1704896540
transform 1 0 26220 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111_279
timestamp 1704896540
transform 1 0 26772 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_281
timestamp 1704896540
transform 1 0 26956 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_293
timestamp 1704896540
transform 1 0 28060 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_305
timestamp 1704896540
transform 1 0 29164 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_317
timestamp 1704896540
transform 1 0 30268 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_111_329
timestamp 1704896540
transform 1 0 31372 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111_335
timestamp 1704896540
transform 1 0 31924 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_337
timestamp 1704896540
transform 1 0 32108 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_349
timestamp 1704896540
transform 1 0 33212 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_361
timestamp 1704896540
transform 1 0 34316 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_373
timestamp 1704896540
transform 1 0 35420 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_111_385
timestamp 1704896540
transform 1 0 36524 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111_391
timestamp 1704896540
transform 1 0 37076 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_393
timestamp 1704896540
transform 1 0 37260 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_405
timestamp 1704896540
transform 1 0 38364 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_417
timestamp 1704896540
transform 1 0 39468 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_3
timestamp 1704896540
transform 1 0 1380 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_15
timestamp 1704896540
transform 1 0 2484 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_112_27
timestamp 1704896540
transform 1 0 3588 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_29
timestamp 1704896540
transform 1 0 3772 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_41
timestamp 1704896540
transform 1 0 4876 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_53
timestamp 1704896540
transform 1 0 5980 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_65
timestamp 1704896540
transform 1 0 7084 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_112_77
timestamp 1704896540
transform 1 0 8188 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_112_83
timestamp 1704896540
transform 1 0 8740 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_85
timestamp 1704896540
transform 1 0 8924 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_97
timestamp 1704896540
transform 1 0 10028 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_109
timestamp 1704896540
transform 1 0 11132 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_121
timestamp 1704896540
transform 1 0 12236 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_112_133
timestamp 1704896540
transform 1 0 13340 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_112_139
timestamp 1704896540
transform 1 0 13892 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_141
timestamp 1704896540
transform 1 0 14076 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_153
timestamp 1704896540
transform 1 0 15180 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_165
timestamp 1704896540
transform 1 0 16284 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_112_177
timestamp 1704896540
transform 1 0 17388 0 1 63104
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_183
timestamp 1704896540
transform 1 0 17940 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_112_195
timestamp 1704896540
transform 1 0 19044 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_197
timestamp 1704896540
transform 1 0 19228 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_209
timestamp 1704896540
transform 1 0 20332 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_221
timestamp 1704896540
transform 1 0 21436 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_233
timestamp 1704896540
transform 1 0 22540 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_112_245
timestamp 1704896540
transform 1 0 23644 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_112_251
timestamp 1704896540
transform 1 0 24196 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_253
timestamp 1704896540
transform 1 0 24380 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_265
timestamp 1704896540
transform 1 0 25484 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_112_279
timestamp 1704896540
transform 1 0 26772 0 1 63104
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_112_283
timestamp 1704896540
transform 1 0 27140 0 1 63104
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_292
timestamp 1704896540
transform 1 0 27968 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_112_304
timestamp 1704896540
transform 1 0 29072 0 1 63104
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_309
timestamp 1704896540
transform 1 0 29532 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_321
timestamp 1704896540
transform 1 0 30636 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_333
timestamp 1704896540
transform 1 0 31740 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_345
timestamp 1704896540
transform 1 0 32844 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_112_357
timestamp 1704896540
transform 1 0 33948 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_112_363
timestamp 1704896540
transform 1 0 34500 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_365
timestamp 1704896540
transform 1 0 34684 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_377
timestamp 1704896540
transform 1 0 35788 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_389
timestamp 1704896540
transform 1 0 36892 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_401
timestamp 1704896540
transform 1 0 37996 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_112_413
timestamp 1704896540
transform 1 0 39100 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_112_419
timestamp 1704896540
transform 1 0 39652 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_112_421
timestamp 1704896540
transform 1 0 39836 0 1 63104
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_3
timestamp 1704896540
transform 1 0 1380 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_15
timestamp 1704896540
transform 1 0 2484 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_27
timestamp 1704896540
transform 1 0 3588 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_39
timestamp 1704896540
transform 1 0 4692 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_113_51
timestamp 1704896540
transform 1 0 5796 0 -1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_113_55
timestamp 1704896540
transform 1 0 6164 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_57
timestamp 1704896540
transform 1 0 6348 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_69
timestamp 1704896540
transform 1 0 7452 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_81
timestamp 1704896540
transform 1 0 8556 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_93
timestamp 1704896540
transform 1 0 9660 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_113_105
timestamp 1704896540
transform 1 0 10764 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_113_111
timestamp 1704896540
transform 1 0 11316 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_113
timestamp 1704896540
transform 1 0 11500 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_125
timestamp 1704896540
transform 1 0 12604 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_137
timestamp 1704896540
transform 1 0 13708 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_149
timestamp 1704896540
transform 1 0 14812 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_113_161
timestamp 1704896540
transform 1 0 15916 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_113_167
timestamp 1704896540
transform 1 0 16468 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_169
timestamp 1704896540
transform 1 0 16652 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_181
timestamp 1704896540
transform 1 0 17756 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_193
timestamp 1704896540
transform 1 0 18860 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_205
timestamp 1704896540
transform 1 0 19964 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_113_217
timestamp 1704896540
transform 1 0 21068 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_113_223
timestamp 1704896540
transform 1 0 21620 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_225
timestamp 1704896540
transform 1 0 21804 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_237
timestamp 1704896540
transform 1 0 22908 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_249
timestamp 1704896540
transform 1 0 24012 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_261
timestamp 1704896540
transform 1 0 25116 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_113_273
timestamp 1704896540
transform 1 0 26220 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_113_279
timestamp 1704896540
transform 1 0 26772 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_281
timestamp 1704896540
transform 1 0 26956 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_293
timestamp 1704896540
transform 1 0 28060 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_305
timestamp 1704896540
transform 1 0 29164 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_317
timestamp 1704896540
transform 1 0 30268 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_113_329
timestamp 1704896540
transform 1 0 31372 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_113_335
timestamp 1704896540
transform 1 0 31924 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_337
timestamp 1704896540
transform 1 0 32108 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_349
timestamp 1704896540
transform 1 0 33212 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_361
timestamp 1704896540
transform 1 0 34316 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_373
timestamp 1704896540
transform 1 0 35420 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_113_385
timestamp 1704896540
transform 1 0 36524 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_113_391
timestamp 1704896540
transform 1 0 37076 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_405
timestamp 1704896540
transform 1 0 38364 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_417
timestamp 1704896540
transform 1 0 39468 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_3
timestamp 1704896540
transform 1 0 1380 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_15
timestamp 1704896540
transform 1 0 2484 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_114_27
timestamp 1704896540
transform 1 0 3588 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_29
timestamp 1704896540
transform 1 0 3772 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_41
timestamp 1704896540
transform 1 0 4876 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_53
timestamp 1704896540
transform 1 0 5980 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_114_65
timestamp 1704896540
transform 1 0 7084 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_114_80
timestamp 1704896540
transform 1 0 8464 0 1 64192
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_85
timestamp 1704896540
transform 1 0 8924 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_97
timestamp 1704896540
transform 1 0 10028 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_109
timestamp 1704896540
transform 1 0 11132 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_121
timestamp 1704896540
transform 1 0 12236 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_114_133
timestamp 1704896540
transform 1 0 13340 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_114_139
timestamp 1704896540
transform 1 0 13892 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_141
timestamp 1704896540
transform 1 0 14076 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_153
timestamp 1704896540
transform 1 0 15180 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_165
timestamp 1704896540
transform 1 0 16284 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_177
timestamp 1704896540
transform 1 0 17388 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_114_189
timestamp 1704896540
transform 1 0 18492 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_114_195
timestamp 1704896540
transform 1 0 19044 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_114_197
timestamp 1704896540
transform 1 0 19228 0 1 64192
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_114_205
timestamp 1704896540
transform 1 0 19964 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_227
timestamp 1704896540
transform 1 0 21988 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_239
timestamp 1704896540
transform 1 0 23092 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_114_251
timestamp 1704896540
transform 1 0 24196 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_253
timestamp 1704896540
transform 1 0 24380 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_265
timestamp 1704896540
transform 1 0 25484 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_277
timestamp 1704896540
transform 1 0 26588 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_289
timestamp 1704896540
transform 1 0 27692 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_114_301
timestamp 1704896540
transform 1 0 28796 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_114_307
timestamp 1704896540
transform 1 0 29348 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_309
timestamp 1704896540
transform 1 0 29532 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_321
timestamp 1704896540
transform 1 0 30636 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_333
timestamp 1704896540
transform 1 0 31740 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_114_345
timestamp 1704896540
transform 1 0 32844 0 1 64192
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_114_358
timestamp 1704896540
transform 1 0 34040 0 1 64192
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_365
timestamp 1704896540
transform 1 0 34684 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_377
timestamp 1704896540
transform 1 0 35788 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_389
timestamp 1704896540
transform 1 0 36892 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_401
timestamp 1704896540
transform 1 0 37996 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_114_413
timestamp 1704896540
transform 1 0 39100 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_114_419
timestamp 1704896540
transform 1 0 39652 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_114_421
timestamp 1704896540
transform 1 0 39836 0 1 64192
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_3
timestamp 1704896540
transform 1 0 1380 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_15
timestamp 1704896540
transform 1 0 2484 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_27
timestamp 1704896540
transform 1 0 3588 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_39
timestamp 1704896540
transform 1 0 4692 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_115_51
timestamp 1704896540
transform 1 0 5796 0 -1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_115_55
timestamp 1704896540
transform 1 0 6164 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_57
timestamp 1704896540
transform 1 0 6348 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_69
timestamp 1704896540
transform 1 0 7452 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_81
timestamp 1704896540
transform 1 0 8556 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_93
timestamp 1704896540
transform 1 0 9660 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_115_105
timestamp 1704896540
transform 1 0 10764 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_115_111
timestamp 1704896540
transform 1 0 11316 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_113
timestamp 1704896540
transform 1 0 11500 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_125
timestamp 1704896540
transform 1 0 12604 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_137
timestamp 1704896540
transform 1 0 13708 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_149
timestamp 1704896540
transform 1 0 14812 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_115_161
timestamp 1704896540
transform 1 0 15916 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_115_167
timestamp 1704896540
transform 1 0 16468 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_169
timestamp 1704896540
transform 1 0 16652 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_181
timestamp 1704896540
transform 1 0 17756 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_193
timestamp 1704896540
transform 1 0 18860 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_205
timestamp 1704896540
transform 1 0 19964 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_115_217
timestamp 1704896540
transform 1 0 21068 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_115_223
timestamp 1704896540
transform 1 0 21620 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_225
timestamp 1704896540
transform 1 0 21804 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_237
timestamp 1704896540
transform 1 0 22908 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_249
timestamp 1704896540
transform 1 0 24012 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_261
timestamp 1704896540
transform 1 0 25116 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_115_273
timestamp 1704896540
transform 1 0 26220 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_115_279
timestamp 1704896540
transform 1 0 26772 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_281
timestamp 1704896540
transform 1 0 26956 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_293
timestamp 1704896540
transform 1 0 28060 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_305
timestamp 1704896540
transform 1 0 29164 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_317
timestamp 1704896540
transform 1 0 30268 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_115_329
timestamp 1704896540
transform 1 0 31372 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_115_335
timestamp 1704896540
transform 1 0 31924 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_337
timestamp 1704896540
transform 1 0 32108 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_349
timestamp 1704896540
transform 1 0 33212 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_361
timestamp 1704896540
transform 1 0 34316 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_373
timestamp 1704896540
transform 1 0 35420 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_115_385
timestamp 1704896540
transform 1 0 36524 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_115_391
timestamp 1704896540
transform 1 0 37076 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_393
timestamp 1704896540
transform 1 0 37260 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_405
timestamp 1704896540
transform 1 0 38364 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_417
timestamp 1704896540
transform 1 0 39468 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_116_3
timestamp 1704896540
transform 1 0 1380 0 1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_116_7
timestamp 1704896540
transform 1 0 1748 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_116_10
timestamp 1704896540
transform 1 0 2024 0 1 65280
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_116_20
timestamp 1704896540
transform 1 0 2944 0 1 65280
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_116_24
timestamp 1704896540
transform 1 0 3312 0 1 65280
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_29
timestamp 1704896540
transform 1 0 3772 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_41
timestamp 1704896540
transform 1 0 4876 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_53
timestamp 1704896540
transform 1 0 5980 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_65
timestamp 1704896540
transform 1 0 7084 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_116_77
timestamp 1704896540
transform 1 0 8188 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_116_83
timestamp 1704896540
transform 1 0 8740 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_85
timestamp 1704896540
transform 1 0 8924 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_97
timestamp 1704896540
transform 1 0 10028 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_116_109
timestamp 1704896540
transform 1 0 11132 0 1 65280
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_122
timestamp 1704896540
transform 1 0 12328 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_116_134
timestamp 1704896540
transform 1 0 13432 0 1 65280
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_141
timestamp 1704896540
transform 1 0 14076 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_153
timestamp 1704896540
transform 1 0 15180 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_165
timestamp 1704896540
transform 1 0 16284 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_177
timestamp 1704896540
transform 1 0 17388 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_116_189
timestamp 1704896540
transform 1 0 18492 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_116_195
timestamp 1704896540
transform 1 0 19044 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_197
timestamp 1704896540
transform 1 0 19228 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_209
timestamp 1704896540
transform 1 0 20332 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_221
timestamp 1704896540
transform 1 0 21436 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_233
timestamp 1704896540
transform 1 0 22540 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_116_245
timestamp 1704896540
transform 1 0 23644 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_116_251
timestamp 1704896540
transform 1 0 24196 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_253
timestamp 1704896540
transform 1 0 24380 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_265
timestamp 1704896540
transform 1 0 25484 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_277
timestamp 1704896540
transform 1 0 26588 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_289
timestamp 1704896540
transform 1 0 27692 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_116_301
timestamp 1704896540
transform 1 0 28796 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_116_307
timestamp 1704896540
transform 1 0 29348 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_309
timestamp 1704896540
transform 1 0 29532 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_321
timestamp 1704896540
transform 1 0 30636 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_333
timestamp 1704896540
transform 1 0 31740 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_345
timestamp 1704896540
transform 1 0 32844 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_116_357
timestamp 1704896540
transform 1 0 33948 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_116_363
timestamp 1704896540
transform 1 0 34500 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_365
timestamp 1704896540
transform 1 0 34684 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_377
timestamp 1704896540
transform 1 0 35788 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_389
timestamp 1704896540
transform 1 0 36892 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_401
timestamp 1704896540
transform 1 0 37996 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_116_413
timestamp 1704896540
transform 1 0 39100 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_116_419
timestamp 1704896540
transform 1 0 39652 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_116_421
timestamp 1704896540
transform 1 0 39836 0 1 65280
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_3
timestamp 1704896540
transform 1 0 1380 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_15
timestamp 1704896540
transform 1 0 2484 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_117_27
timestamp 1704896540
transform 1 0 3588 0 -1 66368
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_43
timestamp 1704896540
transform 1 0 5060 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_117_55
timestamp 1704896540
transform 1 0 6164 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_57
timestamp 1704896540
transform 1 0 6348 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_69
timestamp 1704896540
transform 1 0 7452 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_81
timestamp 1704896540
transform 1 0 8556 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_93
timestamp 1704896540
transform 1 0 9660 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_117_105
timestamp 1704896540
transform 1 0 10764 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_117_111
timestamp 1704896540
transform 1 0 11316 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_113
timestamp 1704896540
transform 1 0 11500 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_125
timestamp 1704896540
transform 1 0 12604 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_137
timestamp 1704896540
transform 1 0 13708 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_149
timestamp 1704896540
transform 1 0 14812 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_117_161
timestamp 1704896540
transform 1 0 15916 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_117_167
timestamp 1704896540
transform 1 0 16468 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_169
timestamp 1704896540
transform 1 0 16652 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_181
timestamp 1704896540
transform 1 0 17756 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_193
timestamp 1704896540
transform 1 0 18860 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_205
timestamp 1704896540
transform 1 0 19964 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_117_217
timestamp 1704896540
transform 1 0 21068 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_117_223
timestamp 1704896540
transform 1 0 21620 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_225
timestamp 1704896540
transform 1 0 21804 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_237
timestamp 1704896540
transform 1 0 22908 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_249
timestamp 1704896540
transform 1 0 24012 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_261
timestamp 1704896540
transform 1 0 25116 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_117_273
timestamp 1704896540
transform 1 0 26220 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_117_279
timestamp 1704896540
transform 1 0 26772 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_281
timestamp 1704896540
transform 1 0 26956 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_293
timestamp 1704896540
transform 1 0 28060 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_305
timestamp 1704896540
transform 1 0 29164 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_317
timestamp 1704896540
transform 1 0 30268 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_117_329
timestamp 1704896540
transform 1 0 31372 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_117_335
timestamp 1704896540
transform 1 0 31924 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_337
timestamp 1704896540
transform 1 0 32108 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_349
timestamp 1704896540
transform 1 0 33212 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_361
timestamp 1704896540
transform 1 0 34316 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_117_390
timestamp 1704896540
transform 1 0 36984 0 -1 66368
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_393
timestamp 1704896540
transform 1 0 37260 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_405
timestamp 1704896540
transform 1 0 38364 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_417
timestamp 1704896540
transform 1 0 39468 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_3
timestamp 1704896540
transform 1 0 1380 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_15
timestamp 1704896540
transform 1 0 2484 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_118_27
timestamp 1704896540
transform 1 0 3588 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_29
timestamp 1704896540
transform 1 0 3772 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_41
timestamp 1704896540
transform 1 0 4876 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_53
timestamp 1704896540
transform 1 0 5980 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_118_65
timestamp 1704896540
transform 1 0 7084 0 1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118_78
timestamp 1704896540
transform 1 0 8280 0 1 66368
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_85
timestamp 1704896540
transform 1 0 8924 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_97
timestamp 1704896540
transform 1 0 10028 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_109
timestamp 1704896540
transform 1 0 11132 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_121
timestamp 1704896540
transform 1 0 12236 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118_133
timestamp 1704896540
transform 1 0 13340 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_118_139
timestamp 1704896540
transform 1 0 13892 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_141
timestamp 1704896540
transform 1 0 14076 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_153
timestamp 1704896540
transform 1 0 15180 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_165
timestamp 1704896540
transform 1 0 16284 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_177
timestamp 1704896540
transform 1 0 17388 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118_189
timestamp 1704896540
transform 1 0 18492 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_118_195
timestamp 1704896540
transform 1 0 19044 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_197
timestamp 1704896540
transform 1 0 19228 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_209
timestamp 1704896540
transform 1 0 20332 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_221
timestamp 1704896540
transform 1 0 21436 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_233
timestamp 1704896540
transform 1 0 22540 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118_245
timestamp 1704896540
transform 1 0 23644 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_118_251
timestamp 1704896540
transform 1 0 24196 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_253
timestamp 1704896540
transform 1 0 24380 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118_265
timestamp 1704896540
transform 1 0 25484 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_118_271
timestamp 1704896540
transform 1 0 26036 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_281
timestamp 1704896540
transform 1 0 26956 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_293
timestamp 1704896540
transform 1 0 28060 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_118_305
timestamp 1704896540
transform 1 0 29164 0 1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_322
timestamp 1704896540
transform 1 0 30728 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_334
timestamp 1704896540
transform 1 0 31832 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_346
timestamp 1704896540
transform 1 0 32936 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118_358
timestamp 1704896540
transform 1 0 34040 0 1 66368
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_365
timestamp 1704896540
transform 1 0 34684 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_377
timestamp 1704896540
transform 1 0 35788 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_389
timestamp 1704896540
transform 1 0 36892 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_401
timestamp 1704896540
transform 1 0 37996 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118_413
timestamp 1704896540
transform 1 0 39100 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_118_419
timestamp 1704896540
transform 1 0 39652 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_118_421
timestamp 1704896540
transform 1 0 39836 0 1 66368
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_3
timestamp 1704896540
transform 1 0 1380 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_15
timestamp 1704896540
transform 1 0 2484 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_27
timestamp 1704896540
transform 1 0 3588 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_39
timestamp 1704896540
transform 1 0 4692 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_119_51
timestamp 1704896540
transform 1 0 5796 0 -1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_119_55
timestamp 1704896540
transform 1 0 6164 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_57
timestamp 1704896540
transform 1 0 6348 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_69
timestamp 1704896540
transform 1 0 7452 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_81
timestamp 1704896540
transform 1 0 8556 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_119_106
timestamp 1704896540
transform 1 0 10856 0 -1 67456
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_113
timestamp 1704896540
transform 1 0 11500 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_125
timestamp 1704896540
transform 1 0 12604 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_137
timestamp 1704896540
transform 1 0 13708 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_149
timestamp 1704896540
transform 1 0 14812 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_119_161
timestamp 1704896540
transform 1 0 15916 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_119_167
timestamp 1704896540
transform 1 0 16468 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_169
timestamp 1704896540
transform 1 0 16652 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_119_181
timestamp 1704896540
transform 1 0 17756 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_195
timestamp 1704896540
transform 1 0 19044 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_207
timestamp 1704896540
transform 1 0 20148 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_119_219
timestamp 1704896540
transform 1 0 21252 0 -1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_119_223
timestamp 1704896540
transform 1 0 21620 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_225
timestamp 1704896540
transform 1 0 21804 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_237
timestamp 1704896540
transform 1 0 22908 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_249
timestamp 1704896540
transform 1 0 24012 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_261
timestamp 1704896540
transform 1 0 25116 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_119_273
timestamp 1704896540
transform 1 0 26220 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_119_279
timestamp 1704896540
transform 1 0 26772 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_281
timestamp 1704896540
transform 1 0 26956 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_293
timestamp 1704896540
transform 1 0 28060 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_305
timestamp 1704896540
transform 1 0 29164 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_317
timestamp 1704896540
transform 1 0 30268 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_119_329
timestamp 1704896540
transform 1 0 31372 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_119_335
timestamp 1704896540
transform 1 0 31924 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_337
timestamp 1704896540
transform 1 0 32108 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_349
timestamp 1704896540
transform 1 0 33212 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_361
timestamp 1704896540
transform 1 0 34316 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_373
timestamp 1704896540
transform 1 0 35420 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_119_385
timestamp 1704896540
transform 1 0 36524 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_119_391
timestamp 1704896540
transform 1 0 37076 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_119_415
timestamp 1704896540
transform 1 0 39284 0 -1 67456
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_120_15
timestamp 1704896540
transform 1 0 2484 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_120_27
timestamp 1704896540
transform 1 0 3588 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_120_29
timestamp 1704896540
transform 1 0 3772 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_120_41
timestamp 1704896540
transform 1 0 4876 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_120_53
timestamp 1704896540
transform 1 0 5980 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_120_65
timestamp 1704896540
transform 1 0 7084 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_120_77
timestamp 1704896540
transform 1 0 8188 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_120_83
timestamp 1704896540
transform 1 0 8740 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_120_85
timestamp 1704896540
transform 1 0 8924 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_120_97
timestamp 1704896540
transform 1 0 10028 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_120_109
timestamp 1704896540
transform 1 0 11132 0 1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_120_117
timestamp 1704896540
transform 1 0 11868 0 1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_120_121
timestamp 1704896540
transform 1 0 12236 0 1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_120_136
timestamp 1704896540
transform 1 0 13616 0 1 67456
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_120_141
timestamp 1704896540
transform 1 0 14076 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_120_153
timestamp 1704896540
transform 1 0 15180 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_120_165
timestamp 1704896540
transform 1 0 16284 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_120_177
timestamp 1704896540
transform 1 0 17388 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_120_189
timestamp 1704896540
transform 1 0 18492 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_120_195
timestamp 1704896540
transform 1 0 19044 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_120_197
timestamp 1704896540
transform 1 0 19228 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_120_209
timestamp 1704896540
transform 1 0 20332 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_120_221
timestamp 1704896540
transform 1 0 21436 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_120_233
timestamp 1704896540
transform 1 0 22540 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_120_245
timestamp 1704896540
transform 1 0 23644 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_120_251
timestamp 1704896540
transform 1 0 24196 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_120_253
timestamp 1704896540
transform 1 0 24380 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_120_265
timestamp 1704896540
transform 1 0 25484 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_120_277
timestamp 1704896540
transform 1 0 26588 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_120_289
timestamp 1704896540
transform 1 0 27692 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_120_301
timestamp 1704896540
transform 1 0 28796 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_120_307
timestamp 1704896540
transform 1 0 29348 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_120_309
timestamp 1704896540
transform 1 0 29532 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_120_321
timestamp 1704896540
transform 1 0 30636 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_120_333
timestamp 1704896540
transform 1 0 31740 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_120_345
timestamp 1704896540
transform 1 0 32844 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_120_357
timestamp 1704896540
transform 1 0 33948 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_120_363
timestamp 1704896540
transform 1 0 34500 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_120_365
timestamp 1704896540
transform 1 0 34684 0 1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_120_369
timestamp 1704896540
transform 1 0 35052 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_120_383
timestamp 1704896540
transform 1 0 36340 0 1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_120_393
timestamp 1704896540
transform 1 0 37260 0 1 67456
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_120_402
timestamp 1704896540
transform 1 0 38088 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_120_414
timestamp 1704896540
transform 1 0 39192 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_120_421
timestamp 1704896540
transform 1 0 39836 0 1 67456
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_121_3
timestamp 1704896540
transform 1 0 1380 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_121_15
timestamp 1704896540
transform 1 0 2484 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_121_27
timestamp 1704896540
transform 1 0 3588 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_121_39
timestamp 1704896540
transform 1 0 4692 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_121_51
timestamp 1704896540
transform 1 0 5796 0 -1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_121_55
timestamp 1704896540
transform 1 0 6164 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_121_57
timestamp 1704896540
transform 1 0 6348 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_121_69
timestamp 1704896540
transform 1 0 7452 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_121_81
timestamp 1704896540
transform 1 0 8556 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_121_93
timestamp 1704896540
transform 1 0 9660 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_121_105
timestamp 1704896540
transform 1 0 10764 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_121_111
timestamp 1704896540
transform 1 0 11316 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_121_113
timestamp 1704896540
transform 1 0 11500 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_121_125
timestamp 1704896540
transform 1 0 12604 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_121_137
timestamp 1704896540
transform 1 0 13708 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_121_149
timestamp 1704896540
transform 1 0 14812 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_121_161
timestamp 1704896540
transform 1 0 15916 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_121_167
timestamp 1704896540
transform 1 0 16468 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_121_169
timestamp 1704896540
transform 1 0 16652 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_121_181
timestamp 1704896540
transform 1 0 17756 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_121_193
timestamp 1704896540
transform 1 0 18860 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_121_205
timestamp 1704896540
transform 1 0 19964 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_121_217
timestamp 1704896540
transform 1 0 21068 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_121_223
timestamp 1704896540
transform 1 0 21620 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_121_225
timestamp 1704896540
transform 1 0 21804 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_121_259
timestamp 1704896540
transform 1 0 24932 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_121_271
timestamp 1704896540
transform 1 0 26036 0 -1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_121_279
timestamp 1704896540
transform 1 0 26772 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_121_281
timestamp 1704896540
transform 1 0 26956 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_121_293
timestamp 1704896540
transform 1 0 28060 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_121_305
timestamp 1704896540
transform 1 0 29164 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_121_317
timestamp 1704896540
transform 1 0 30268 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_121_329
timestamp 1704896540
transform 1 0 31372 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_121_335
timestamp 1704896540
transform 1 0 31924 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_121_337
timestamp 1704896540
transform 1 0 32108 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_121_349
timestamp 1704896540
transform 1 0 33212 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_121_361
timestamp 1704896540
transform 1 0 34316 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_121_373
timestamp 1704896540
transform 1 0 35420 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_121_385
timestamp 1704896540
transform 1 0 36524 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_121_391
timestamp 1704896540
transform 1 0 37076 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_121_393
timestamp 1704896540
transform 1 0 37260 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_121_405
timestamp 1704896540
transform 1 0 38364 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_121_417
timestamp 1704896540
transform 1 0 39468 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_122_3
timestamp 1704896540
transform 1 0 1380 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_122_15
timestamp 1704896540
transform 1 0 2484 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_122_27
timestamp 1704896540
transform 1 0 3588 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_122_29
timestamp 1704896540
transform 1 0 3772 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_122_41
timestamp 1704896540
transform 1 0 4876 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_122_53
timestamp 1704896540
transform 1 0 5980 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_122_65
timestamp 1704896540
transform 1 0 7084 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_122_77
timestamp 1704896540
transform 1 0 8188 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_122_83
timestamp 1704896540
transform 1 0 8740 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_122_85
timestamp 1704896540
transform 1 0 8924 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_122_97
timestamp 1704896540
transform 1 0 10028 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_122_109
timestamp 1704896540
transform 1 0 11132 0 1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_122_117
timestamp 1704896540
transform 1 0 11868 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_122_135
timestamp 1704896540
transform 1 0 13524 0 1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_122_139
timestamp 1704896540
transform 1 0 13892 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_122_141
timestamp 1704896540
transform 1 0 14076 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_122_153
timestamp 1704896540
transform 1 0 15180 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_122_165
timestamp 1704896540
transform 1 0 16284 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_122_177
timestamp 1704896540
transform 1 0 17388 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_122_189
timestamp 1704896540
transform 1 0 18492 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_122_195
timestamp 1704896540
transform 1 0 19044 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_122_197
timestamp 1704896540
transform 1 0 19228 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_122_209
timestamp 1704896540
transform 1 0 20332 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_122_221
timestamp 1704896540
transform 1 0 21436 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_122_233
timestamp 1704896540
transform 1 0 22540 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_122_245
timestamp 1704896540
transform 1 0 23644 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_122_251
timestamp 1704896540
transform 1 0 24196 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_122_253
timestamp 1704896540
transform 1 0 24380 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_122_265
timestamp 1704896540
transform 1 0 25484 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_122_277
timestamp 1704896540
transform 1 0 26588 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_122_289
timestamp 1704896540
transform 1 0 27692 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_122_301
timestamp 1704896540
transform 1 0 28796 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_122_307
timestamp 1704896540
transform 1 0 29348 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_122_309
timestamp 1704896540
transform 1 0 29532 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_122_321
timestamp 1704896540
transform 1 0 30636 0 1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_122_325
timestamp 1704896540
transform 1 0 31004 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_122_331
timestamp 1704896540
transform 1 0 31556 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_122_343
timestamp 1704896540
transform 1 0 32660 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_122_355
timestamp 1704896540
transform 1 0 33764 0 1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_122_363
timestamp 1704896540
transform 1 0 34500 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_122_365
timestamp 1704896540
transform 1 0 34684 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_122_377
timestamp 1704896540
transform 1 0 35788 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_122_389
timestamp 1704896540
transform 1 0 36892 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_122_401
timestamp 1704896540
transform 1 0 37996 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_122_413
timestamp 1704896540
transform 1 0 39100 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_122_419
timestamp 1704896540
transform 1 0 39652 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_122_421
timestamp 1704896540
transform 1 0 39836 0 1 68544
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_123_3
timestamp 1704896540
transform 1 0 1380 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_123_15
timestamp 1704896540
transform 1 0 2484 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_123_27
timestamp 1704896540
transform 1 0 3588 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_123_29
timestamp 1704896540
transform 1 0 3772 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_123_41
timestamp 1704896540
transform 1 0 4876 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_123_53
timestamp 1704896540
transform 1 0 5980 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_123_57
timestamp 1704896540
transform 1 0 6348 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_123_63
timestamp 1704896540
transform 1 0 6900 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_123_73
timestamp 1704896540
transform 1 0 7820 0 -1 69632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_123_81
timestamp 1704896540
transform 1 0 8556 0 -1 69632
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_123_85
timestamp 1704896540
transform 1 0 8924 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_123_97
timestamp 1704896540
transform 1 0 10028 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_123_109
timestamp 1704896540
transform 1 0 11132 0 -1 69632
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_123_113
timestamp 1704896540
transform 1 0 11500 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_123_125
timestamp 1704896540
transform 1 0 12604 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_123_137
timestamp 1704896540
transform 1 0 13708 0 -1 69632
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_123_141
timestamp 1704896540
transform 1 0 14076 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_123_153
timestamp 1704896540
transform 1 0 15180 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_123_165
timestamp 1704896540
transform 1 0 16284 0 -1 69632
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_123_169
timestamp 1704896540
transform 1 0 16652 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_123_181
timestamp 1704896540
transform 1 0 17756 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_123_193
timestamp 1704896540
transform 1 0 18860 0 -1 69632
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_123_197
timestamp 1704896540
transform 1 0 19228 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_123_209
timestamp 1704896540
transform 1 0 20332 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_123_221
timestamp 1704896540
transform 1 0 21436 0 -1 69632
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_123_234
timestamp 1704896540
transform 1 0 22632 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_123_246
timestamp 1704896540
transform 1 0 23736 0 -1 69632
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_123_253
timestamp 1704896540
transform 1 0 24380 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_123_265
timestamp 1704896540
transform 1 0 25484 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_123_277
timestamp 1704896540
transform 1 0 26588 0 -1 69632
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_123_281
timestamp 1704896540
transform 1 0 26956 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_123_293
timestamp 1704896540
transform 1 0 28060 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_123_305
timestamp 1704896540
transform 1 0 29164 0 -1 69632
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_123_309
timestamp 1704896540
transform 1 0 29532 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_123_321
timestamp 1704896540
transform 1 0 30636 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_123_333
timestamp 1704896540
transform 1 0 31740 0 -1 69632
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_123_337
timestamp 1704896540
transform 1 0 32108 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_123_349
timestamp 1704896540
transform 1 0 33212 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_123_361
timestamp 1704896540
transform 1 0 34316 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_123_365
timestamp 1704896540
transform 1 0 34684 0 -1 69632
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_123_379
timestamp 1704896540
transform 1 0 35972 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_123_391
timestamp 1704896540
transform 1 0 37076 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_123_393
timestamp 1704896540
transform 1 0 37260 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_123_405
timestamp 1704896540
transform 1 0 38364 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_123_417
timestamp 1704896540
transform 1 0 39468 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_123_421
timestamp 1704896540
transform 1 0 39836 0 -1 69632
box -38 -48 774 592
use sky130_fd_sc_hd__buf_8  input1
timestamp 1704896540
transform 1 0 1380 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_12  input2
timestamp 1704896540
transform 1 0 1380 0 -1 58752
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  input3
timestamp 1704896540
transform 1 0 1380 0 -1 50048
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_8  input4
timestamp 1704896540
transform 1 0 1380 0 -1 40256
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_4  input5 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 1380 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input6
timestamp 1704896540
transform 1 0 1380 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_16  input7
timestamp 1704896540
transform 1 0 1380 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_8  input8
timestamp 1704896540
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  input9
timestamp 1704896540
transform -1 0 40572 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  input10
timestamp 1704896540
transform -1 0 40572 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_8  input11
timestamp 1704896540
transform -1 0 40572 0 -1 50048
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_12  input12
timestamp 1704896540
transform -1 0 40572 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_8  input13
timestamp 1704896540
transform -1 0 40572 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  input14
timestamp 1704896540
transform -1 0 40572 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  input15
timestamp 1704896540
transform -1 0 40572 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_8  input16
timestamp 1704896540
transform -1 0 40572 0 -1 4352
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  input17
timestamp 1704896540
transform 1 0 34960 0 -1 69632
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_6  input18 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 21804 0 -1 69632
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  input19
timestamp 1704896540
transform 1 0 6992 0 -1 69632
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  max_cap30 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 16928 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  max_cap31
timestamp 1704896540
transform 1 0 18676 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  max_cap32
timestamp 1704896540
transform 1 0 33580 0 -1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  output20 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 39376 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output21
timestamp 1704896540
transform 1 0 34132 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output22
timestamp 1704896540
transform 1 0 28980 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output23
timestamp 1704896540
transform 1 0 23644 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output24
timestamp 1704896540
transform -1 0 18768 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output25
timestamp 1704896540
transform -1 0 13524 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  output26
timestamp 1704896540
transform -1 0 8280 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_8  output27
timestamp 1704896540
transform -1 0 3036 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_124
timestamp 1704896540
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1704896540
transform -1 0 40848 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_125
timestamp 1704896540
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1704896540
transform -1 0 40848 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_126
timestamp 1704896540
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1704896540
transform -1 0 40848 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_127
timestamp 1704896540
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1704896540
transform -1 0 40848 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_128
timestamp 1704896540
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1704896540
transform -1 0 40848 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_129
timestamp 1704896540
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1704896540
transform -1 0 40848 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_130
timestamp 1704896540
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1704896540
transform -1 0 40848 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_131
timestamp 1704896540
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1704896540
transform -1 0 40848 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_132
timestamp 1704896540
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1704896540
transform -1 0 40848 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_133
timestamp 1704896540
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1704896540
transform -1 0 40848 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_134
timestamp 1704896540
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1704896540
transform -1 0 40848 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_135
timestamp 1704896540
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1704896540
transform -1 0 40848 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_136
timestamp 1704896540
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1704896540
transform -1 0 40848 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_137
timestamp 1704896540
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1704896540
transform -1 0 40848 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_138
timestamp 1704896540
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1704896540
transform -1 0 40848 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_139
timestamp 1704896540
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1704896540
transform -1 0 40848 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_140
timestamp 1704896540
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1704896540
transform -1 0 40848 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_141
timestamp 1704896540
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1704896540
transform -1 0 40848 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_142
timestamp 1704896540
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1704896540
transform -1 0 40848 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_143
timestamp 1704896540
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1704896540
transform -1 0 40848 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_144
timestamp 1704896540
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1704896540
transform -1 0 40848 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_145
timestamp 1704896540
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1704896540
transform -1 0 40848 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_146
timestamp 1704896540
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1704896540
transform -1 0 40848 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_147
timestamp 1704896540
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 1704896540
transform -1 0 40848 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_148
timestamp 1704896540
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 1704896540
transform -1 0 40848 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_149
timestamp 1704896540
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 1704896540
transform -1 0 40848 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_150
timestamp 1704896540
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 1704896540
transform -1 0 40848 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_151
timestamp 1704896540
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 1704896540
transform -1 0 40848 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_152
timestamp 1704896540
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 1704896540
transform -1 0 40848 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_153
timestamp 1704896540
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 1704896540
transform -1 0 40848 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_154
timestamp 1704896540
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 1704896540
transform -1 0 40848 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_155
timestamp 1704896540
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp 1704896540
transform -1 0 40848 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_156
timestamp 1704896540
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp 1704896540
transform -1 0 40848 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_157
timestamp 1704896540
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp 1704896540
transform -1 0 40848 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Left_158
timestamp 1704896540
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Right_34
timestamp 1704896540
transform -1 0 40848 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Left_159
timestamp 1704896540
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Right_35
timestamp 1704896540
transform -1 0 40848 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Left_160
timestamp 1704896540
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Right_36
timestamp 1704896540
transform -1 0 40848 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Left_161
timestamp 1704896540
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Right_37
timestamp 1704896540
transform -1 0 40848 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Left_162
timestamp 1704896540
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Right_38
timestamp 1704896540
transform -1 0 40848 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Left_163
timestamp 1704896540
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Right_39
timestamp 1704896540
transform -1 0 40848 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Left_164
timestamp 1704896540
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Right_40
timestamp 1704896540
transform -1 0 40848 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Left_165
timestamp 1704896540
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Right_41
timestamp 1704896540
transform -1 0 40848 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Left_166
timestamp 1704896540
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Right_42
timestamp 1704896540
transform -1 0 40848 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Left_167
timestamp 1704896540
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Right_43
timestamp 1704896540
transform -1 0 40848 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Left_168
timestamp 1704896540
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Right_44
timestamp 1704896540
transform -1 0 40848 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Left_169
timestamp 1704896540
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Right_45
timestamp 1704896540
transform -1 0 40848 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Left_170
timestamp 1704896540
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Right_46
timestamp 1704896540
transform -1 0 40848 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Left_171
timestamp 1704896540
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Right_47
timestamp 1704896540
transform -1 0 40848 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Left_172
timestamp 1704896540
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Right_48
timestamp 1704896540
transform -1 0 40848 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_Left_173
timestamp 1704896540
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_Right_49
timestamp 1704896540
transform -1 0 40848 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_Left_174
timestamp 1704896540
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_Right_50
timestamp 1704896540
transform -1 0 40848 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_Left_175
timestamp 1704896540
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_Right_51
timestamp 1704896540
transform -1 0 40848 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_Left_176
timestamp 1704896540
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_Right_52
timestamp 1704896540
transform -1 0 40848 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_Left_177
timestamp 1704896540
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_Right_53
timestamp 1704896540
transform -1 0 40848 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_Left_178
timestamp 1704896540
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_Right_54
timestamp 1704896540
transform -1 0 40848 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_Left_179
timestamp 1704896540
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_Right_55
timestamp 1704896540
transform -1 0 40848 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_Left_180
timestamp 1704896540
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_Right_56
timestamp 1704896540
transform -1 0 40848 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_Left_181
timestamp 1704896540
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_Right_57
timestamp 1704896540
transform -1 0 40848 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_Left_182
timestamp 1704896540
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_Right_58
timestamp 1704896540
transform -1 0 40848 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_Left_183
timestamp 1704896540
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_Right_59
timestamp 1704896540
transform -1 0 40848 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_Left_184
timestamp 1704896540
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_Right_60
timestamp 1704896540
transform -1 0 40848 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_Left_185
timestamp 1704896540
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_Right_61
timestamp 1704896540
transform -1 0 40848 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_Left_186
timestamp 1704896540
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_Right_62
timestamp 1704896540
transform -1 0 40848 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_Left_187
timestamp 1704896540
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_Right_63
timestamp 1704896540
transform -1 0 40848 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_Left_188
timestamp 1704896540
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_Right_64
timestamp 1704896540
transform -1 0 40848 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_Left_189
timestamp 1704896540
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_Right_65
timestamp 1704896540
transform -1 0 40848 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_Left_190
timestamp 1704896540
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_Right_66
timestamp 1704896540
transform -1 0 40848 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_Left_191
timestamp 1704896540
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_Right_67
timestamp 1704896540
transform -1 0 40848 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_Left_192
timestamp 1704896540
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_Right_68
timestamp 1704896540
transform -1 0 40848 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_Left_193
timestamp 1704896540
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_Right_69
timestamp 1704896540
transform -1 0 40848 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_Left_194
timestamp 1704896540
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_Right_70
timestamp 1704896540
transform -1 0 40848 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_Left_195
timestamp 1704896540
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_Right_71
timestamp 1704896540
transform -1 0 40848 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_Left_196
timestamp 1704896540
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_Right_72
timestamp 1704896540
transform -1 0 40848 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_Left_197
timestamp 1704896540
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_Right_73
timestamp 1704896540
transform -1 0 40848 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_74_Left_198
timestamp 1704896540
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_74_Right_74
timestamp 1704896540
transform -1 0 40848 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_75_Left_199
timestamp 1704896540
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_75_Right_75
timestamp 1704896540
transform -1 0 40848 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_76_Left_200
timestamp 1704896540
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_76_Right_76
timestamp 1704896540
transform -1 0 40848 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_77_Left_201
timestamp 1704896540
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_77_Right_77
timestamp 1704896540
transform -1 0 40848 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_78_Left_202
timestamp 1704896540
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_78_Right_78
timestamp 1704896540
transform -1 0 40848 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_79_Left_203
timestamp 1704896540
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_79_Right_79
timestamp 1704896540
transform -1 0 40848 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_80_Left_204
timestamp 1704896540
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_80_Right_80
timestamp 1704896540
transform -1 0 40848 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_81_Left_205
timestamp 1704896540
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_81_Right_81
timestamp 1704896540
transform -1 0 40848 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_82_Left_206
timestamp 1704896540
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_82_Right_82
timestamp 1704896540
transform -1 0 40848 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_83_Left_207
timestamp 1704896540
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_83_Right_83
timestamp 1704896540
transform -1 0 40848 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_84_Left_208
timestamp 1704896540
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_84_Right_84
timestamp 1704896540
transform -1 0 40848 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_85_Left_209
timestamp 1704896540
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_85_Right_85
timestamp 1704896540
transform -1 0 40848 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_86_Left_210
timestamp 1704896540
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_86_Right_86
timestamp 1704896540
transform -1 0 40848 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_87_Left_211
timestamp 1704896540
transform 1 0 1104 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_87_Right_87
timestamp 1704896540
transform -1 0 40848 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_88_Left_212
timestamp 1704896540
transform 1 0 1104 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_88_Right_88
timestamp 1704896540
transform -1 0 40848 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_89_Left_213
timestamp 1704896540
transform 1 0 1104 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_89_Right_89
timestamp 1704896540
transform -1 0 40848 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_90_Left_214
timestamp 1704896540
transform 1 0 1104 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_90_Right_90
timestamp 1704896540
transform -1 0 40848 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_91_Left_215
timestamp 1704896540
transform 1 0 1104 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_91_Right_91
timestamp 1704896540
transform -1 0 40848 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_92_Left_216
timestamp 1704896540
transform 1 0 1104 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_92_Right_92
timestamp 1704896540
transform -1 0 40848 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_93_Left_217
timestamp 1704896540
transform 1 0 1104 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_93_Right_93
timestamp 1704896540
transform -1 0 40848 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_94_Left_218
timestamp 1704896540
transform 1 0 1104 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_94_Right_94
timestamp 1704896540
transform -1 0 40848 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_95_Left_219
timestamp 1704896540
transform 1 0 1104 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_95_Right_95
timestamp 1704896540
transform -1 0 40848 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_96_Left_220
timestamp 1704896540
transform 1 0 1104 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_96_Right_96
timestamp 1704896540
transform -1 0 40848 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_97_Left_221
timestamp 1704896540
transform 1 0 1104 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_97_Right_97
timestamp 1704896540
transform -1 0 40848 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_98_Left_222
timestamp 1704896540
transform 1 0 1104 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_98_Right_98
timestamp 1704896540
transform -1 0 40848 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_99_Left_223
timestamp 1704896540
transform 1 0 1104 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_99_Right_99
timestamp 1704896540
transform -1 0 40848 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_100_Left_224
timestamp 1704896540
transform 1 0 1104 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_100_Right_100
timestamp 1704896540
transform -1 0 40848 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_101_Left_225
timestamp 1704896540
transform 1 0 1104 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_101_Right_101
timestamp 1704896540
transform -1 0 40848 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_102_Left_226
timestamp 1704896540
transform 1 0 1104 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_102_Right_102
timestamp 1704896540
transform -1 0 40848 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_103_Left_227
timestamp 1704896540
transform 1 0 1104 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_103_Right_103
timestamp 1704896540
transform -1 0 40848 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_104_Left_228
timestamp 1704896540
transform 1 0 1104 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_104_Right_104
timestamp 1704896540
transform -1 0 40848 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_105_Left_229
timestamp 1704896540
transform 1 0 1104 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_105_Right_105
timestamp 1704896540
transform -1 0 40848 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_106_Left_230
timestamp 1704896540
transform 1 0 1104 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_106_Right_106
timestamp 1704896540
transform -1 0 40848 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_107_Left_231
timestamp 1704896540
transform 1 0 1104 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_107_Right_107
timestamp 1704896540
transform -1 0 40848 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_108_Left_232
timestamp 1704896540
transform 1 0 1104 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_108_Right_108
timestamp 1704896540
transform -1 0 40848 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_109_Left_233
timestamp 1704896540
transform 1 0 1104 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_109_Right_109
timestamp 1704896540
transform -1 0 40848 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_110_Left_234
timestamp 1704896540
transform 1 0 1104 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_110_Right_110
timestamp 1704896540
transform -1 0 40848 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_111_Left_235
timestamp 1704896540
transform 1 0 1104 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_111_Right_111
timestamp 1704896540
transform -1 0 40848 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_112_Left_236
timestamp 1704896540
transform 1 0 1104 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_112_Right_112
timestamp 1704896540
transform -1 0 40848 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_113_Left_237
timestamp 1704896540
transform 1 0 1104 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_113_Right_113
timestamp 1704896540
transform -1 0 40848 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_114_Left_238
timestamp 1704896540
transform 1 0 1104 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_114_Right_114
timestamp 1704896540
transform -1 0 40848 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_115_Left_239
timestamp 1704896540
transform 1 0 1104 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_115_Right_115
timestamp 1704896540
transform -1 0 40848 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_116_Left_240
timestamp 1704896540
transform 1 0 1104 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_116_Right_116
timestamp 1704896540
transform -1 0 40848 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_117_Left_241
timestamp 1704896540
transform 1 0 1104 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_117_Right_117
timestamp 1704896540
transform -1 0 40848 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_118_Left_242
timestamp 1704896540
transform 1 0 1104 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_118_Right_118
timestamp 1704896540
transform -1 0 40848 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_119_Left_243
timestamp 1704896540
transform 1 0 1104 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_119_Right_119
timestamp 1704896540
transform -1 0 40848 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_120_Left_244
timestamp 1704896540
transform 1 0 1104 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_120_Right_120
timestamp 1704896540
transform -1 0 40848 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_121_Left_245
timestamp 1704896540
transform 1 0 1104 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_121_Right_121
timestamp 1704896540
transform -1 0 40848 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_122_Left_246
timestamp 1704896540
transform 1 0 1104 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_122_Right_122
timestamp 1704896540
transform -1 0 40848 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_123_Left_247
timestamp 1704896540
transform 1 0 1104 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_123_Right_123
timestamp 1704896540
transform -1 0 40848 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  rebuffer1
timestamp 1704896540
transform -1 0 28980 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 32660 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  rebuffer3
timestamp 1704896540
transform 1 0 12420 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  rebuffer4
timestamp 1704896540
transform -1 0 30360 0 1 59840
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  rebuffer5
timestamp 1704896540
transform 1 0 31188 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  rebuffer6
timestamp 1704896540
transform 1 0 20516 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  rebuffer7
timestamp 1704896540
transform -1 0 25300 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  rebuffer8 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 24472 0 1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer9
timestamp 1704896540
transform 1 0 29992 0 1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__buf_6  rebuffer10
timestamp 1704896540
transform 1 0 30636 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer11
timestamp 1704896540
transform 1 0 7728 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  rebuffer12
timestamp 1704896540
transform 1 0 15456 0 1 54400
box -38 -48 958 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer13
timestamp 1704896540
transform 1 0 35144 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer14
timestamp 1704896540
transform 1 0 6716 0 1 58752
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  rebuffer15
timestamp 1704896540
transform -1 0 25944 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer16
timestamp 1704896540
transform -1 0 23920 0 -1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer17
timestamp 1704896540
transform -1 0 17480 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  rebuffer18
timestamp 1704896540
transform 1 0 33212 0 1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer19
timestamp 1704896540
transform 1 0 38732 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer20
timestamp 1704896540
transform -1 0 20976 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s4s_1  rebuffer21 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 11408 0 -1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__buf_12  rebuffer22
timestamp 1704896540
transform 1 0 6992 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer23
timestamp 1704896540
transform -1 0 7636 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  rebuffer24
timestamp 1704896540
transform 1 0 19228 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  rebuffer25
timestamp 1704896540
transform 1 0 15272 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer26
timestamp 1704896540
transform -1 0 33212 0 1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  rebuffer27
timestamp 1704896540
transform 1 0 17020 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s4s_1  rebuffer28
timestamp 1704896540
transform -1 0 39284 0 1 40256
box -38 -48 958 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer29
timestamp 1704896540
transform -1 0 7728 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer30
timestamp 1704896540
transform -1 0 36340 0 -1 52224
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_248 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_249
timestamp 1704896540
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_250
timestamp 1704896540
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_251
timestamp 1704896540
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_252
timestamp 1704896540
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_253
timestamp 1704896540
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_254
timestamp 1704896540
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_255
timestamp 1704896540
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_256
timestamp 1704896540
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_257
timestamp 1704896540
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_258
timestamp 1704896540
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_259
timestamp 1704896540
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_260
timestamp 1704896540
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_261
timestamp 1704896540
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_262
timestamp 1704896540
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_263
timestamp 1704896540
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_264
timestamp 1704896540
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_265
timestamp 1704896540
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_266
timestamp 1704896540
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_267
timestamp 1704896540
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_268
timestamp 1704896540
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_269
timestamp 1704896540
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_270
timestamp 1704896540
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_271
timestamp 1704896540
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_272
timestamp 1704896540
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_273
timestamp 1704896540
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_274
timestamp 1704896540
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_275
timestamp 1704896540
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_276
timestamp 1704896540
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_277
timestamp 1704896540
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_278
timestamp 1704896540
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_279
timestamp 1704896540
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_280
timestamp 1704896540
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_281
timestamp 1704896540
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_282
timestamp 1704896540
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_283
timestamp 1704896540
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_284
timestamp 1704896540
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_285
timestamp 1704896540
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_286
timestamp 1704896540
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_287
timestamp 1704896540
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_288
timestamp 1704896540
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_289
timestamp 1704896540
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_290
timestamp 1704896540
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_291
timestamp 1704896540
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_292
timestamp 1704896540
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_293
timestamp 1704896540
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_294
timestamp 1704896540
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_295
timestamp 1704896540
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_296
timestamp 1704896540
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_297
timestamp 1704896540
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_298
timestamp 1704896540
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_299
timestamp 1704896540
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_300
timestamp 1704896540
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_301
timestamp 1704896540
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_302
timestamp 1704896540
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_303
timestamp 1704896540
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_304
timestamp 1704896540
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_305
timestamp 1704896540
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_306
timestamp 1704896540
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_307
timestamp 1704896540
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_308
timestamp 1704896540
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_309
timestamp 1704896540
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_310
timestamp 1704896540
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_311
timestamp 1704896540
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_312
timestamp 1704896540
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_313
timestamp 1704896540
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_314
timestamp 1704896540
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_315
timestamp 1704896540
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_316
timestamp 1704896540
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_317
timestamp 1704896540
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_318
timestamp 1704896540
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_319
timestamp 1704896540
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_320
timestamp 1704896540
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_321
timestamp 1704896540
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_322
timestamp 1704896540
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_323
timestamp 1704896540
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_324
timestamp 1704896540
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_325
timestamp 1704896540
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_326
timestamp 1704896540
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_327
timestamp 1704896540
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_328
timestamp 1704896540
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_329
timestamp 1704896540
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_330
timestamp 1704896540
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_331
timestamp 1704896540
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_332
timestamp 1704896540
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_333
timestamp 1704896540
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_334
timestamp 1704896540
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_335
timestamp 1704896540
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_336
timestamp 1704896540
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_337
timestamp 1704896540
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_338
timestamp 1704896540
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_339
timestamp 1704896540
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_340
timestamp 1704896540
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_341
timestamp 1704896540
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_342
timestamp 1704896540
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_343
timestamp 1704896540
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_344
timestamp 1704896540
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_345
timestamp 1704896540
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_346
timestamp 1704896540
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_347
timestamp 1704896540
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_348
timestamp 1704896540
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_349
timestamp 1704896540
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_350
timestamp 1704896540
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_351
timestamp 1704896540
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_352
timestamp 1704896540
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_353
timestamp 1704896540
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_354
timestamp 1704896540
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_355
timestamp 1704896540
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_356
timestamp 1704896540
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_357
timestamp 1704896540
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_358
timestamp 1704896540
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_359
timestamp 1704896540
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_360
timestamp 1704896540
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_361
timestamp 1704896540
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_362
timestamp 1704896540
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_363
timestamp 1704896540
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_364
timestamp 1704896540
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_365
timestamp 1704896540
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_366
timestamp 1704896540
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_367
timestamp 1704896540
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_368
timestamp 1704896540
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_369
timestamp 1704896540
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_370
timestamp 1704896540
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_371
timestamp 1704896540
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_372
timestamp 1704896540
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_373
timestamp 1704896540
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_374
timestamp 1704896540
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_375
timestamp 1704896540
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_376
timestamp 1704896540
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_377
timestamp 1704896540
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_378
timestamp 1704896540
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_379
timestamp 1704896540
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_380
timestamp 1704896540
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_381
timestamp 1704896540
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_382
timestamp 1704896540
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_383
timestamp 1704896540
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_384
timestamp 1704896540
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_385
timestamp 1704896540
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_386
timestamp 1704896540
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_387
timestamp 1704896540
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_388
timestamp 1704896540
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_389
timestamp 1704896540
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_390
timestamp 1704896540
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_391
timestamp 1704896540
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_392
timestamp 1704896540
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_393
timestamp 1704896540
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_394
timestamp 1704896540
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_395
timestamp 1704896540
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_396
timestamp 1704896540
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_397
timestamp 1704896540
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_398
timestamp 1704896540
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_399
timestamp 1704896540
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_400
timestamp 1704896540
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_401
timestamp 1704896540
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_402
timestamp 1704896540
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_403
timestamp 1704896540
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_404
timestamp 1704896540
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_405
timestamp 1704896540
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_406
timestamp 1704896540
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_407
timestamp 1704896540
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_408
timestamp 1704896540
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_409
timestamp 1704896540
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_410
timestamp 1704896540
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_411
timestamp 1704896540
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_412
timestamp 1704896540
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_413
timestamp 1704896540
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_414
timestamp 1704896540
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_415
timestamp 1704896540
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_416
timestamp 1704896540
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_417
timestamp 1704896540
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_418
timestamp 1704896540
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_419
timestamp 1704896540
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_420
timestamp 1704896540
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_421
timestamp 1704896540
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_422
timestamp 1704896540
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_423
timestamp 1704896540
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_424
timestamp 1704896540
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_425
timestamp 1704896540
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_426
timestamp 1704896540
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_427
timestamp 1704896540
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_428
timestamp 1704896540
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_429
timestamp 1704896540
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_430
timestamp 1704896540
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_431
timestamp 1704896540
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_432
timestamp 1704896540
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_433
timestamp 1704896540
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_434
timestamp 1704896540
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_435
timestamp 1704896540
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_436
timestamp 1704896540
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_437
timestamp 1704896540
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_438
timestamp 1704896540
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_439
timestamp 1704896540
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_440
timestamp 1704896540
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_441
timestamp 1704896540
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_442
timestamp 1704896540
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_443
timestamp 1704896540
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_444
timestamp 1704896540
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_445
timestamp 1704896540
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_446
timestamp 1704896540
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_447
timestamp 1704896540
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_448
timestamp 1704896540
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_449
timestamp 1704896540
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_450
timestamp 1704896540
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_451
timestamp 1704896540
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_452
timestamp 1704896540
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_453
timestamp 1704896540
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_454
timestamp 1704896540
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_455
timestamp 1704896540
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_456
timestamp 1704896540
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_457
timestamp 1704896540
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_458
timestamp 1704896540
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_459
timestamp 1704896540
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_460
timestamp 1704896540
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_461
timestamp 1704896540
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_462
timestamp 1704896540
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_463
timestamp 1704896540
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_464
timestamp 1704896540
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_465
timestamp 1704896540
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_466
timestamp 1704896540
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_467
timestamp 1704896540
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_468
timestamp 1704896540
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_469
timestamp 1704896540
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_470
timestamp 1704896540
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_471
timestamp 1704896540
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_472
timestamp 1704896540
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_473
timestamp 1704896540
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_474
timestamp 1704896540
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_475
timestamp 1704896540
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_476
timestamp 1704896540
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_477
timestamp 1704896540
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_478
timestamp 1704896540
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_479
timestamp 1704896540
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_480
timestamp 1704896540
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_481
timestamp 1704896540
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_482
timestamp 1704896540
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_483
timestamp 1704896540
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_484
timestamp 1704896540
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_485
timestamp 1704896540
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_486
timestamp 1704896540
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_487
timestamp 1704896540
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_488
timestamp 1704896540
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_489
timestamp 1704896540
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_490
timestamp 1704896540
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_491
timestamp 1704896540
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_492
timestamp 1704896540
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_493
timestamp 1704896540
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_494
timestamp 1704896540
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_495
timestamp 1704896540
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_496
timestamp 1704896540
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_497
timestamp 1704896540
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_498
timestamp 1704896540
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_499
timestamp 1704896540
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_500
timestamp 1704896540
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_501
timestamp 1704896540
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_502
timestamp 1704896540
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_503
timestamp 1704896540
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_504
timestamp 1704896540
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_505
timestamp 1704896540
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_506
timestamp 1704896540
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_507
timestamp 1704896540
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_508
timestamp 1704896540
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_509
timestamp 1704896540
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_510
timestamp 1704896540
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_511
timestamp 1704896540
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_512
timestamp 1704896540
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_513
timestamp 1704896540
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_514
timestamp 1704896540
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_515
timestamp 1704896540
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_516
timestamp 1704896540
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_517
timestamp 1704896540
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_518
timestamp 1704896540
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_519
timestamp 1704896540
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_520
timestamp 1704896540
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_521
timestamp 1704896540
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_522
timestamp 1704896540
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_523
timestamp 1704896540
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_524
timestamp 1704896540
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_525
timestamp 1704896540
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_526
timestamp 1704896540
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_527
timestamp 1704896540
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_528
timestamp 1704896540
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_529
timestamp 1704896540
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_530
timestamp 1704896540
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_531
timestamp 1704896540
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_532
timestamp 1704896540
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_533
timestamp 1704896540
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_534
timestamp 1704896540
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_535
timestamp 1704896540
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_536
timestamp 1704896540
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_537
timestamp 1704896540
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_538
timestamp 1704896540
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_539
timestamp 1704896540
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_540
timestamp 1704896540
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_541
timestamp 1704896540
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_542
timestamp 1704896540
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_543
timestamp 1704896540
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_544
timestamp 1704896540
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_545
timestamp 1704896540
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_546
timestamp 1704896540
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_547
timestamp 1704896540
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_548
timestamp 1704896540
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_549
timestamp 1704896540
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_550
timestamp 1704896540
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_551
timestamp 1704896540
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_552
timestamp 1704896540
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_553
timestamp 1704896540
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_554
timestamp 1704896540
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_555
timestamp 1704896540
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_556
timestamp 1704896540
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_557
timestamp 1704896540
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_558
timestamp 1704896540
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_559
timestamp 1704896540
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_560
timestamp 1704896540
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_561
timestamp 1704896540
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_562
timestamp 1704896540
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_563
timestamp 1704896540
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_564
timestamp 1704896540
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_565
timestamp 1704896540
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_566
timestamp 1704896540
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_567
timestamp 1704896540
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_568
timestamp 1704896540
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_569
timestamp 1704896540
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_570
timestamp 1704896540
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_571
timestamp 1704896540
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_572
timestamp 1704896540
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_573
timestamp 1704896540
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_574
timestamp 1704896540
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_575
timestamp 1704896540
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_576
timestamp 1704896540
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_577
timestamp 1704896540
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_578
timestamp 1704896540
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_579
timestamp 1704896540
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_580
timestamp 1704896540
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_581
timestamp 1704896540
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_582
timestamp 1704896540
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_583
timestamp 1704896540
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_584
timestamp 1704896540
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_585
timestamp 1704896540
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_586
timestamp 1704896540
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_587
timestamp 1704896540
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_588
timestamp 1704896540
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_589
timestamp 1704896540
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_590
timestamp 1704896540
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_591
timestamp 1704896540
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_592
timestamp 1704896540
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_593
timestamp 1704896540
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_594
timestamp 1704896540
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_595
timestamp 1704896540
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_596
timestamp 1704896540
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_597
timestamp 1704896540
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_598
timestamp 1704896540
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_599
timestamp 1704896540
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_600
timestamp 1704896540
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_601
timestamp 1704896540
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_602
timestamp 1704896540
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_603
timestamp 1704896540
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_604
timestamp 1704896540
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_605
timestamp 1704896540
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_606
timestamp 1704896540
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_607
timestamp 1704896540
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_608
timestamp 1704896540
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_609
timestamp 1704896540
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_610
timestamp 1704896540
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_611
timestamp 1704896540
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_612
timestamp 1704896540
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_613
timestamp 1704896540
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_614
timestamp 1704896540
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_615
timestamp 1704896540
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_616
timestamp 1704896540
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_617
timestamp 1704896540
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_618
timestamp 1704896540
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_619
timestamp 1704896540
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_620
timestamp 1704896540
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_621
timestamp 1704896540
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_622
timestamp 1704896540
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_623
timestamp 1704896540
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_624
timestamp 1704896540
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_625
timestamp 1704896540
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_626
timestamp 1704896540
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_627
timestamp 1704896540
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_628
timestamp 1704896540
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_629
timestamp 1704896540
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_630
timestamp 1704896540
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_631
timestamp 1704896540
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_632
timestamp 1704896540
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_633
timestamp 1704896540
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_634
timestamp 1704896540
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_635
timestamp 1704896540
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_636
timestamp 1704896540
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_637
timestamp 1704896540
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_638
timestamp 1704896540
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_639
timestamp 1704896540
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_640
timestamp 1704896540
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_641
timestamp 1704896540
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_642
timestamp 1704896540
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_643
timestamp 1704896540
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_644
timestamp 1704896540
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_645
timestamp 1704896540
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_646
timestamp 1704896540
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_647
timestamp 1704896540
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_648
timestamp 1704896540
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_649
timestamp 1704896540
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_650
timestamp 1704896540
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_651
timestamp 1704896540
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_652
timestamp 1704896540
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_653
timestamp 1704896540
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_654
timestamp 1704896540
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_655
timestamp 1704896540
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_656
timestamp 1704896540
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_657
timestamp 1704896540
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_658
timestamp 1704896540
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_659
timestamp 1704896540
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_660
timestamp 1704896540
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_661
timestamp 1704896540
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_662
timestamp 1704896540
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_663
timestamp 1704896540
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_664
timestamp 1704896540
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_665
timestamp 1704896540
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_666
timestamp 1704896540
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_667
timestamp 1704896540
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_668
timestamp 1704896540
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_669
timestamp 1704896540
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_670
timestamp 1704896540
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_671
timestamp 1704896540
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_672
timestamp 1704896540
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_673
timestamp 1704896540
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_674
timestamp 1704896540
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_675
timestamp 1704896540
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_676
timestamp 1704896540
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_677
timestamp 1704896540
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_678
timestamp 1704896540
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_679
timestamp 1704896540
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_680
timestamp 1704896540
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_681
timestamp 1704896540
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_682
timestamp 1704896540
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_683
timestamp 1704896540
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_684
timestamp 1704896540
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_685
timestamp 1704896540
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_686
timestamp 1704896540
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_687
timestamp 1704896540
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_688
timestamp 1704896540
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_689
timestamp 1704896540
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_690
timestamp 1704896540
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_691
timestamp 1704896540
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_692
timestamp 1704896540
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_693
timestamp 1704896540
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_694
timestamp 1704896540
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_695
timestamp 1704896540
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_696
timestamp 1704896540
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_697
timestamp 1704896540
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_698
timestamp 1704896540
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_699
timestamp 1704896540
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_700
timestamp 1704896540
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_701
timestamp 1704896540
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_702
timestamp 1704896540
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_703
timestamp 1704896540
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_704
timestamp 1704896540
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_705
timestamp 1704896540
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_706
timestamp 1704896540
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_707
timestamp 1704896540
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_708
timestamp 1704896540
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_709
timestamp 1704896540
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_710
timestamp 1704896540
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_711
timestamp 1704896540
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_712
timestamp 1704896540
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_713
timestamp 1704896540
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_714
timestamp 1704896540
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_715
timestamp 1704896540
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_716
timestamp 1704896540
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_717
timestamp 1704896540
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_718
timestamp 1704896540
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_719
timestamp 1704896540
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_720
timestamp 1704896540
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_721
timestamp 1704896540
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_722
timestamp 1704896540
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_723
timestamp 1704896540
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_724
timestamp 1704896540
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_725
timestamp 1704896540
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_726
timestamp 1704896540
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_727
timestamp 1704896540
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_728
timestamp 1704896540
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_729
timestamp 1704896540
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_730
timestamp 1704896540
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_731
timestamp 1704896540
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_732
timestamp 1704896540
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_733
timestamp 1704896540
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_734
timestamp 1704896540
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_735
timestamp 1704896540
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_736
timestamp 1704896540
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_737
timestamp 1704896540
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_738
timestamp 1704896540
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_739
timestamp 1704896540
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_740
timestamp 1704896540
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_741
timestamp 1704896540
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_742
timestamp 1704896540
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_743
timestamp 1704896540
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_744
timestamp 1704896540
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_745
timestamp 1704896540
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_746
timestamp 1704896540
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_747
timestamp 1704896540
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_748
timestamp 1704896540
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_749
timestamp 1704896540
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_750
timestamp 1704896540
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_751
timestamp 1704896540
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_752
timestamp 1704896540
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_753
timestamp 1704896540
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_754
timestamp 1704896540
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_755
timestamp 1704896540
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_756
timestamp 1704896540
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_757
timestamp 1704896540
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_758
timestamp 1704896540
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_759
timestamp 1704896540
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_760
timestamp 1704896540
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_761
timestamp 1704896540
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_762
timestamp 1704896540
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_763
timestamp 1704896540
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_764
timestamp 1704896540
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_765
timestamp 1704896540
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_766
timestamp 1704896540
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_767
timestamp 1704896540
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_768
timestamp 1704896540
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_769
timestamp 1704896540
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_770
timestamp 1704896540
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_771
timestamp 1704896540
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_772
timestamp 1704896540
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_773
timestamp 1704896540
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_774
timestamp 1704896540
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_775
timestamp 1704896540
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_776
timestamp 1704896540
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_777
timestamp 1704896540
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_778
timestamp 1704896540
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_779
timestamp 1704896540
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_780
timestamp 1704896540
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_781
timestamp 1704896540
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_782
timestamp 1704896540
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_783
timestamp 1704896540
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_784
timestamp 1704896540
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_785
timestamp 1704896540
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_786
timestamp 1704896540
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_787
timestamp 1704896540
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_788
timestamp 1704896540
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_789
timestamp 1704896540
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_790
timestamp 1704896540
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_791
timestamp 1704896540
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_792
timestamp 1704896540
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_793
timestamp 1704896540
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_794
timestamp 1704896540
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_795
timestamp 1704896540
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_796
timestamp 1704896540
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_797
timestamp 1704896540
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_798
timestamp 1704896540
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_799
timestamp 1704896540
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_800
timestamp 1704896540
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_801
timestamp 1704896540
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_802
timestamp 1704896540
transform 1 0 39744 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_803
timestamp 1704896540
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_804
timestamp 1704896540
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_805
timestamp 1704896540
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_806
timestamp 1704896540
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_807
timestamp 1704896540
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_808
timestamp 1704896540
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_809
timestamp 1704896540
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_810
timestamp 1704896540
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_811
timestamp 1704896540
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_812
timestamp 1704896540
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_813
timestamp 1704896540
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_814
timestamp 1704896540
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_815
timestamp 1704896540
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_816
timestamp 1704896540
transform 1 0 34592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_817
timestamp 1704896540
transform 1 0 39744 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_818
timestamp 1704896540
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_819
timestamp 1704896540
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_820
timestamp 1704896540
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_821
timestamp 1704896540
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_822
timestamp 1704896540
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_823
timestamp 1704896540
transform 1 0 32016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_824
timestamp 1704896540
transform 1 0 37168 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_825
timestamp 1704896540
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_826
timestamp 1704896540
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_827
timestamp 1704896540
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_828
timestamp 1704896540
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_829
timestamp 1704896540
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_830
timestamp 1704896540
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_831
timestamp 1704896540
transform 1 0 34592 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_832
timestamp 1704896540
transform 1 0 39744 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_833
timestamp 1704896540
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_834
timestamp 1704896540
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_835
timestamp 1704896540
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_836
timestamp 1704896540
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_837
timestamp 1704896540
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_838
timestamp 1704896540
transform 1 0 32016 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_839
timestamp 1704896540
transform 1 0 37168 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_840
timestamp 1704896540
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_841
timestamp 1704896540
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_842
timestamp 1704896540
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_843
timestamp 1704896540
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_844
timestamp 1704896540
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_845
timestamp 1704896540
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_846
timestamp 1704896540
transform 1 0 34592 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_847
timestamp 1704896540
transform 1 0 39744 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_848
timestamp 1704896540
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_849
timestamp 1704896540
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_850
timestamp 1704896540
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_851
timestamp 1704896540
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_852
timestamp 1704896540
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_853
timestamp 1704896540
transform 1 0 32016 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_854
timestamp 1704896540
transform 1 0 37168 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_855
timestamp 1704896540
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_856
timestamp 1704896540
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_857
timestamp 1704896540
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_858
timestamp 1704896540
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_859
timestamp 1704896540
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_860
timestamp 1704896540
transform 1 0 29440 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_861
timestamp 1704896540
transform 1 0 34592 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_862
timestamp 1704896540
transform 1 0 39744 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_863
timestamp 1704896540
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_864
timestamp 1704896540
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_865
timestamp 1704896540
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_866
timestamp 1704896540
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_867
timestamp 1704896540
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_868
timestamp 1704896540
transform 1 0 32016 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_869
timestamp 1704896540
transform 1 0 37168 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_870
timestamp 1704896540
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_871
timestamp 1704896540
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_872
timestamp 1704896540
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_873
timestamp 1704896540
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_874
timestamp 1704896540
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_875
timestamp 1704896540
transform 1 0 29440 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_876
timestamp 1704896540
transform 1 0 34592 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_877
timestamp 1704896540
transform 1 0 39744 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_83_878
timestamp 1704896540
transform 1 0 6256 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_83_879
timestamp 1704896540
transform 1 0 11408 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_83_880
timestamp 1704896540
transform 1 0 16560 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_83_881
timestamp 1704896540
transform 1 0 21712 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_83_882
timestamp 1704896540
transform 1 0 26864 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_83_883
timestamp 1704896540
transform 1 0 32016 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_83_884
timestamp 1704896540
transform 1 0 37168 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_885
timestamp 1704896540
transform 1 0 3680 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_886
timestamp 1704896540
transform 1 0 8832 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_887
timestamp 1704896540
transform 1 0 13984 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_888
timestamp 1704896540
transform 1 0 19136 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_889
timestamp 1704896540
transform 1 0 24288 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_890
timestamp 1704896540
transform 1 0 29440 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_891
timestamp 1704896540
transform 1 0 34592 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_892
timestamp 1704896540
transform 1 0 39744 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_85_893
timestamp 1704896540
transform 1 0 6256 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_85_894
timestamp 1704896540
transform 1 0 11408 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_85_895
timestamp 1704896540
transform 1 0 16560 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_85_896
timestamp 1704896540
transform 1 0 21712 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_85_897
timestamp 1704896540
transform 1 0 26864 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_85_898
timestamp 1704896540
transform 1 0 32016 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_85_899
timestamp 1704896540
transform 1 0 37168 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_900
timestamp 1704896540
transform 1 0 3680 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_901
timestamp 1704896540
transform 1 0 8832 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_902
timestamp 1704896540
transform 1 0 13984 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_903
timestamp 1704896540
transform 1 0 19136 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_904
timestamp 1704896540
transform 1 0 24288 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_905
timestamp 1704896540
transform 1 0 29440 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_906
timestamp 1704896540
transform 1 0 34592 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_907
timestamp 1704896540
transform 1 0 39744 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_87_908
timestamp 1704896540
transform 1 0 6256 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_87_909
timestamp 1704896540
transform 1 0 11408 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_87_910
timestamp 1704896540
transform 1 0 16560 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_87_911
timestamp 1704896540
transform 1 0 21712 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_87_912
timestamp 1704896540
transform 1 0 26864 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_87_913
timestamp 1704896540
transform 1 0 32016 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_87_914
timestamp 1704896540
transform 1 0 37168 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_915
timestamp 1704896540
transform 1 0 3680 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_916
timestamp 1704896540
transform 1 0 8832 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_917
timestamp 1704896540
transform 1 0 13984 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_918
timestamp 1704896540
transform 1 0 19136 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_919
timestamp 1704896540
transform 1 0 24288 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_920
timestamp 1704896540
transform 1 0 29440 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_921
timestamp 1704896540
transform 1 0 34592 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_922
timestamp 1704896540
transform 1 0 39744 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_89_923
timestamp 1704896540
transform 1 0 6256 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_89_924
timestamp 1704896540
transform 1 0 11408 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_89_925
timestamp 1704896540
transform 1 0 16560 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_89_926
timestamp 1704896540
transform 1 0 21712 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_89_927
timestamp 1704896540
transform 1 0 26864 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_89_928
timestamp 1704896540
transform 1 0 32016 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_89_929
timestamp 1704896540
transform 1 0 37168 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_930
timestamp 1704896540
transform 1 0 3680 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_931
timestamp 1704896540
transform 1 0 8832 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_932
timestamp 1704896540
transform 1 0 13984 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_933
timestamp 1704896540
transform 1 0 19136 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_934
timestamp 1704896540
transform 1 0 24288 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_935
timestamp 1704896540
transform 1 0 29440 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_936
timestamp 1704896540
transform 1 0 34592 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_937
timestamp 1704896540
transform 1 0 39744 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_91_938
timestamp 1704896540
transform 1 0 6256 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_91_939
timestamp 1704896540
transform 1 0 11408 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_91_940
timestamp 1704896540
transform 1 0 16560 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_91_941
timestamp 1704896540
transform 1 0 21712 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_91_942
timestamp 1704896540
transform 1 0 26864 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_91_943
timestamp 1704896540
transform 1 0 32016 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_91_944
timestamp 1704896540
transform 1 0 37168 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_945
timestamp 1704896540
transform 1 0 3680 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_946
timestamp 1704896540
transform 1 0 8832 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_947
timestamp 1704896540
transform 1 0 13984 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_948
timestamp 1704896540
transform 1 0 19136 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_949
timestamp 1704896540
transform 1 0 24288 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_950
timestamp 1704896540
transform 1 0 29440 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_951
timestamp 1704896540
transform 1 0 34592 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_952
timestamp 1704896540
transform 1 0 39744 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_93_953
timestamp 1704896540
transform 1 0 6256 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_93_954
timestamp 1704896540
transform 1 0 11408 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_93_955
timestamp 1704896540
transform 1 0 16560 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_93_956
timestamp 1704896540
transform 1 0 21712 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_93_957
timestamp 1704896540
transform 1 0 26864 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_93_958
timestamp 1704896540
transform 1 0 32016 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_93_959
timestamp 1704896540
transform 1 0 37168 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_960
timestamp 1704896540
transform 1 0 3680 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_961
timestamp 1704896540
transform 1 0 8832 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_962
timestamp 1704896540
transform 1 0 13984 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_963
timestamp 1704896540
transform 1 0 19136 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_964
timestamp 1704896540
transform 1 0 24288 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_965
timestamp 1704896540
transform 1 0 29440 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_966
timestamp 1704896540
transform 1 0 34592 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_967
timestamp 1704896540
transform 1 0 39744 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_95_968
timestamp 1704896540
transform 1 0 6256 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_95_969
timestamp 1704896540
transform 1 0 11408 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_95_970
timestamp 1704896540
transform 1 0 16560 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_95_971
timestamp 1704896540
transform 1 0 21712 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_95_972
timestamp 1704896540
transform 1 0 26864 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_95_973
timestamp 1704896540
transform 1 0 32016 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_95_974
timestamp 1704896540
transform 1 0 37168 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_975
timestamp 1704896540
transform 1 0 3680 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_976
timestamp 1704896540
transform 1 0 8832 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_977
timestamp 1704896540
transform 1 0 13984 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_978
timestamp 1704896540
transform 1 0 19136 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_979
timestamp 1704896540
transform 1 0 24288 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_980
timestamp 1704896540
transform 1 0 29440 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_981
timestamp 1704896540
transform 1 0 34592 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_982
timestamp 1704896540
transform 1 0 39744 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_983
timestamp 1704896540
transform 1 0 6256 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_984
timestamp 1704896540
transform 1 0 11408 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_985
timestamp 1704896540
transform 1 0 16560 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_986
timestamp 1704896540
transform 1 0 21712 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_987
timestamp 1704896540
transform 1 0 26864 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_988
timestamp 1704896540
transform 1 0 32016 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_989
timestamp 1704896540
transform 1 0 37168 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_990
timestamp 1704896540
transform 1 0 3680 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_991
timestamp 1704896540
transform 1 0 8832 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_992
timestamp 1704896540
transform 1 0 13984 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_993
timestamp 1704896540
transform 1 0 19136 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_994
timestamp 1704896540
transform 1 0 24288 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_995
timestamp 1704896540
transform 1 0 29440 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_996
timestamp 1704896540
transform 1 0 34592 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_997
timestamp 1704896540
transform 1 0 39744 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_99_998
timestamp 1704896540
transform 1 0 6256 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_99_999
timestamp 1704896540
transform 1 0 11408 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_99_1000
timestamp 1704896540
transform 1 0 16560 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_99_1001
timestamp 1704896540
transform 1 0 21712 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_99_1002
timestamp 1704896540
transform 1 0 26864 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_99_1003
timestamp 1704896540
transform 1 0 32016 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_99_1004
timestamp 1704896540
transform 1 0 37168 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_1005
timestamp 1704896540
transform 1 0 3680 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_1006
timestamp 1704896540
transform 1 0 8832 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_1007
timestamp 1704896540
transform 1 0 13984 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_1008
timestamp 1704896540
transform 1 0 19136 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_1009
timestamp 1704896540
transform 1 0 24288 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_1010
timestamp 1704896540
transform 1 0 29440 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_1011
timestamp 1704896540
transform 1 0 34592 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_1012
timestamp 1704896540
transform 1 0 39744 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1013
timestamp 1704896540
transform 1 0 6256 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1014
timestamp 1704896540
transform 1 0 11408 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1015
timestamp 1704896540
transform 1 0 16560 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1016
timestamp 1704896540
transform 1 0 21712 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1017
timestamp 1704896540
transform 1 0 26864 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1018
timestamp 1704896540
transform 1 0 32016 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1019
timestamp 1704896540
transform 1 0 37168 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_102_1020
timestamp 1704896540
transform 1 0 3680 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_102_1021
timestamp 1704896540
transform 1 0 8832 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_102_1022
timestamp 1704896540
transform 1 0 13984 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_102_1023
timestamp 1704896540
transform 1 0 19136 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_102_1024
timestamp 1704896540
transform 1 0 24288 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_102_1025
timestamp 1704896540
transform 1 0 29440 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_102_1026
timestamp 1704896540
transform 1 0 34592 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_102_1027
timestamp 1704896540
transform 1 0 39744 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_103_1028
timestamp 1704896540
transform 1 0 6256 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_103_1029
timestamp 1704896540
transform 1 0 11408 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_103_1030
timestamp 1704896540
transform 1 0 16560 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_103_1031
timestamp 1704896540
transform 1 0 21712 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_103_1032
timestamp 1704896540
transform 1 0 26864 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_103_1033
timestamp 1704896540
transform 1 0 32016 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_103_1034
timestamp 1704896540
transform 1 0 37168 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_104_1035
timestamp 1704896540
transform 1 0 3680 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_104_1036
timestamp 1704896540
transform 1 0 8832 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_104_1037
timestamp 1704896540
transform 1 0 13984 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_104_1038
timestamp 1704896540
transform 1 0 19136 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_104_1039
timestamp 1704896540
transform 1 0 24288 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_104_1040
timestamp 1704896540
transform 1 0 29440 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_104_1041
timestamp 1704896540
transform 1 0 34592 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_104_1042
timestamp 1704896540
transform 1 0 39744 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_105_1043
timestamp 1704896540
transform 1 0 6256 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_105_1044
timestamp 1704896540
transform 1 0 11408 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_105_1045
timestamp 1704896540
transform 1 0 16560 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_105_1046
timestamp 1704896540
transform 1 0 21712 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_105_1047
timestamp 1704896540
transform 1 0 26864 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_105_1048
timestamp 1704896540
transform 1 0 32016 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_105_1049
timestamp 1704896540
transform 1 0 37168 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_1050
timestamp 1704896540
transform 1 0 3680 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_1051
timestamp 1704896540
transform 1 0 8832 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_1052
timestamp 1704896540
transform 1 0 13984 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_1053
timestamp 1704896540
transform 1 0 19136 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_1054
timestamp 1704896540
transform 1 0 24288 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_1055
timestamp 1704896540
transform 1 0 29440 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_1056
timestamp 1704896540
transform 1 0 34592 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_1057
timestamp 1704896540
transform 1 0 39744 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_107_1058
timestamp 1704896540
transform 1 0 6256 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_107_1059
timestamp 1704896540
transform 1 0 11408 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_107_1060
timestamp 1704896540
transform 1 0 16560 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_107_1061
timestamp 1704896540
transform 1 0 21712 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_107_1062
timestamp 1704896540
transform 1 0 26864 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_107_1063
timestamp 1704896540
transform 1 0 32016 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_107_1064
timestamp 1704896540
transform 1 0 37168 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_108_1065
timestamp 1704896540
transform 1 0 3680 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_108_1066
timestamp 1704896540
transform 1 0 8832 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_108_1067
timestamp 1704896540
transform 1 0 13984 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_108_1068
timestamp 1704896540
transform 1 0 19136 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_108_1069
timestamp 1704896540
transform 1 0 24288 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_108_1070
timestamp 1704896540
transform 1 0 29440 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_108_1071
timestamp 1704896540
transform 1 0 34592 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_108_1072
timestamp 1704896540
transform 1 0 39744 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_109_1073
timestamp 1704896540
transform 1 0 6256 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_109_1074
timestamp 1704896540
transform 1 0 11408 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_109_1075
timestamp 1704896540
transform 1 0 16560 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_109_1076
timestamp 1704896540
transform 1 0 21712 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_109_1077
timestamp 1704896540
transform 1 0 26864 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_109_1078
timestamp 1704896540
transform 1 0 32016 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_109_1079
timestamp 1704896540
transform 1 0 37168 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_110_1080
timestamp 1704896540
transform 1 0 3680 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_110_1081
timestamp 1704896540
transform 1 0 8832 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_110_1082
timestamp 1704896540
transform 1 0 13984 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_110_1083
timestamp 1704896540
transform 1 0 19136 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_110_1084
timestamp 1704896540
transform 1 0 24288 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_110_1085
timestamp 1704896540
transform 1 0 29440 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_110_1086
timestamp 1704896540
transform 1 0 34592 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_110_1087
timestamp 1704896540
transform 1 0 39744 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_111_1088
timestamp 1704896540
transform 1 0 6256 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_111_1089
timestamp 1704896540
transform 1 0 11408 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_111_1090
timestamp 1704896540
transform 1 0 16560 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_111_1091
timestamp 1704896540
transform 1 0 21712 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_111_1092
timestamp 1704896540
transform 1 0 26864 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_111_1093
timestamp 1704896540
transform 1 0 32016 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_111_1094
timestamp 1704896540
transform 1 0 37168 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_112_1095
timestamp 1704896540
transform 1 0 3680 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_112_1096
timestamp 1704896540
transform 1 0 8832 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_112_1097
timestamp 1704896540
transform 1 0 13984 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_112_1098
timestamp 1704896540
transform 1 0 19136 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_112_1099
timestamp 1704896540
transform 1 0 24288 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_112_1100
timestamp 1704896540
transform 1 0 29440 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_112_1101
timestamp 1704896540
transform 1 0 34592 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_112_1102
timestamp 1704896540
transform 1 0 39744 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_113_1103
timestamp 1704896540
transform 1 0 6256 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_113_1104
timestamp 1704896540
transform 1 0 11408 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_113_1105
timestamp 1704896540
transform 1 0 16560 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_113_1106
timestamp 1704896540
transform 1 0 21712 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_113_1107
timestamp 1704896540
transform 1 0 26864 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_113_1108
timestamp 1704896540
transform 1 0 32016 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_113_1109
timestamp 1704896540
transform 1 0 37168 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_114_1110
timestamp 1704896540
transform 1 0 3680 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_114_1111
timestamp 1704896540
transform 1 0 8832 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_114_1112
timestamp 1704896540
transform 1 0 13984 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_114_1113
timestamp 1704896540
transform 1 0 19136 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_114_1114
timestamp 1704896540
transform 1 0 24288 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_114_1115
timestamp 1704896540
transform 1 0 29440 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_114_1116
timestamp 1704896540
transform 1 0 34592 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_114_1117
timestamp 1704896540
transform 1 0 39744 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_115_1118
timestamp 1704896540
transform 1 0 6256 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_115_1119
timestamp 1704896540
transform 1 0 11408 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_115_1120
timestamp 1704896540
transform 1 0 16560 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_115_1121
timestamp 1704896540
transform 1 0 21712 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_115_1122
timestamp 1704896540
transform 1 0 26864 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_115_1123
timestamp 1704896540
transform 1 0 32016 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_115_1124
timestamp 1704896540
transform 1 0 37168 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_116_1125
timestamp 1704896540
transform 1 0 3680 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_116_1126
timestamp 1704896540
transform 1 0 8832 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_116_1127
timestamp 1704896540
transform 1 0 13984 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_116_1128
timestamp 1704896540
transform 1 0 19136 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_116_1129
timestamp 1704896540
transform 1 0 24288 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_116_1130
timestamp 1704896540
transform 1 0 29440 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_116_1131
timestamp 1704896540
transform 1 0 34592 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_116_1132
timestamp 1704896540
transform 1 0 39744 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1133
timestamp 1704896540
transform 1 0 6256 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1134
timestamp 1704896540
transform 1 0 11408 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1135
timestamp 1704896540
transform 1 0 16560 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1136
timestamp 1704896540
transform 1 0 21712 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1137
timestamp 1704896540
transform 1 0 26864 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1138
timestamp 1704896540
transform 1 0 32016 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1139
timestamp 1704896540
transform 1 0 37168 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_1140
timestamp 1704896540
transform 1 0 3680 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_1141
timestamp 1704896540
transform 1 0 8832 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_1142
timestamp 1704896540
transform 1 0 13984 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_1143
timestamp 1704896540
transform 1 0 19136 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_1144
timestamp 1704896540
transform 1 0 24288 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_1145
timestamp 1704896540
transform 1 0 29440 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_1146
timestamp 1704896540
transform 1 0 34592 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_1147
timestamp 1704896540
transform 1 0 39744 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_1148
timestamp 1704896540
transform 1 0 6256 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_1149
timestamp 1704896540
transform 1 0 11408 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_1150
timestamp 1704896540
transform 1 0 16560 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_1151
timestamp 1704896540
transform 1 0 21712 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_1152
timestamp 1704896540
transform 1 0 26864 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_1153
timestamp 1704896540
transform 1 0 32016 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_1154
timestamp 1704896540
transform 1 0 37168 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1155
timestamp 1704896540
transform 1 0 3680 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1156
timestamp 1704896540
transform 1 0 8832 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1157
timestamp 1704896540
transform 1 0 13984 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1158
timestamp 1704896540
transform 1 0 19136 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1159
timestamp 1704896540
transform 1 0 24288 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1160
timestamp 1704896540
transform 1 0 29440 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1161
timestamp 1704896540
transform 1 0 34592 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1162
timestamp 1704896540
transform 1 0 39744 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_1163
timestamp 1704896540
transform 1 0 6256 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_1164
timestamp 1704896540
transform 1 0 11408 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_1165
timestamp 1704896540
transform 1 0 16560 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_1166
timestamp 1704896540
transform 1 0 21712 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_1167
timestamp 1704896540
transform 1 0 26864 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_1168
timestamp 1704896540
transform 1 0 32016 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_1169
timestamp 1704896540
transform 1 0 37168 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_1170
timestamp 1704896540
transform 1 0 3680 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_1171
timestamp 1704896540
transform 1 0 8832 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_1172
timestamp 1704896540
transform 1 0 13984 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_1173
timestamp 1704896540
transform 1 0 19136 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_1174
timestamp 1704896540
transform 1 0 24288 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_1175
timestamp 1704896540
transform 1 0 29440 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_1176
timestamp 1704896540
transform 1 0 34592 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_1177
timestamp 1704896540
transform 1 0 39744 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_1178
timestamp 1704896540
transform 1 0 3680 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_1179
timestamp 1704896540
transform 1 0 6256 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_1180
timestamp 1704896540
transform 1 0 8832 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_1181
timestamp 1704896540
transform 1 0 11408 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_1182
timestamp 1704896540
transform 1 0 13984 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_1183
timestamp 1704896540
transform 1 0 16560 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_1184
timestamp 1704896540
transform 1 0 19136 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_1185
timestamp 1704896540
transform 1 0 21712 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_1186
timestamp 1704896540
transform 1 0 24288 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_1187
timestamp 1704896540
transform 1 0 26864 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_1188
timestamp 1704896540
transform 1 0 29440 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_1189
timestamp 1704896540
transform 1 0 32016 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_1190
timestamp 1704896540
transform 1 0 34592 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_1191
timestamp 1704896540
transform 1 0 37168 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_1192
timestamp 1704896540
transform 1 0 39744 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  wire28
timestamp 1704896540
transform -1 0 10580 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  wire29
timestamp 1704896540
transform -1 0 24748 0 1 57664
box -38 -48 406 592
<< labels >>
flabel metal3 s 0 67192 800 67312 0 FreeSans 480 0 0 0 A[0]
port 0 nsew signal input
flabel metal3 s 0 58216 800 58336 0 FreeSans 480 0 0 0 A[1]
port 1 nsew signal input
flabel metal3 s 0 49240 800 49360 0 FreeSans 480 0 0 0 A[2]
port 2 nsew signal input
flabel metal3 s 0 40264 800 40384 0 FreeSans 480 0 0 0 A[3]
port 3 nsew signal input
flabel metal3 s 0 31288 800 31408 0 FreeSans 480 0 0 0 A[4]
port 4 nsew signal input
flabel metal3 s 0 22312 800 22432 0 FreeSans 480 0 0 0 A[5]
port 5 nsew signal input
flabel metal3 s 0 13336 800 13456 0 FreeSans 480 0 0 0 A[6]
port 6 nsew signal input
flabel metal3 s 0 4360 800 4480 0 FreeSans 480 0 0 0 A[7]
port 7 nsew signal input
flabel metal3 s 41200 67192 42000 67312 0 FreeSans 480 0 0 0 B[0]
port 8 nsew signal input
flabel metal3 s 41200 58216 42000 58336 0 FreeSans 480 0 0 0 B[1]
port 9 nsew signal input
flabel metal3 s 41200 49240 42000 49360 0 FreeSans 480 0 0 0 B[2]
port 10 nsew signal input
flabel metal3 s 41200 40264 42000 40384 0 FreeSans 480 0 0 0 B[3]
port 11 nsew signal input
flabel metal3 s 41200 31288 42000 31408 0 FreeSans 480 0 0 0 B[4]
port 12 nsew signal input
flabel metal3 s 41200 22312 42000 22432 0 FreeSans 480 0 0 0 B[5]
port 13 nsew signal input
flabel metal3 s 41200 13336 42000 13456 0 FreeSans 480 0 0 0 B[6]
port 14 nsew signal input
flabel metal3 s 41200 4360 42000 4480 0 FreeSans 480 0 0 0 B[7]
port 15 nsew signal input
flabel metal4 s 2604 2128 2924 69680 0 FreeSans 1920 90 0 0 VGND
port 16 nsew ground bidirectional
flabel metal4 s 7604 2128 7924 69680 0 FreeSans 1920 90 0 0 VGND
port 16 nsew ground bidirectional
flabel metal4 s 12604 2128 12924 69680 0 FreeSans 1920 90 0 0 VGND
port 16 nsew ground bidirectional
flabel metal4 s 17604 2128 17924 69680 0 FreeSans 1920 90 0 0 VGND
port 16 nsew ground bidirectional
flabel metal4 s 22604 2128 22924 69680 0 FreeSans 1920 90 0 0 VGND
port 16 nsew ground bidirectional
flabel metal4 s 27604 2128 27924 69680 0 FreeSans 1920 90 0 0 VGND
port 16 nsew ground bidirectional
flabel metal4 s 32604 2128 32924 69680 0 FreeSans 1920 90 0 0 VGND
port 16 nsew ground bidirectional
flabel metal4 s 37604 2128 37924 69680 0 FreeSans 1920 90 0 0 VGND
port 16 nsew ground bidirectional
flabel metal5 s 1056 3676 40896 3996 0 FreeSans 2560 0 0 0 VGND
port 16 nsew ground bidirectional
flabel metal5 s 1056 8676 40896 8996 0 FreeSans 2560 0 0 0 VGND
port 16 nsew ground bidirectional
flabel metal5 s 1056 13676 40896 13996 0 FreeSans 2560 0 0 0 VGND
port 16 nsew ground bidirectional
flabel metal5 s 1056 18676 40896 18996 0 FreeSans 2560 0 0 0 VGND
port 16 nsew ground bidirectional
flabel metal5 s 1056 23676 40896 23996 0 FreeSans 2560 0 0 0 VGND
port 16 nsew ground bidirectional
flabel metal5 s 1056 28676 40896 28996 0 FreeSans 2560 0 0 0 VGND
port 16 nsew ground bidirectional
flabel metal5 s 1056 33676 40896 33996 0 FreeSans 2560 0 0 0 VGND
port 16 nsew ground bidirectional
flabel metal5 s 1056 38676 40896 38996 0 FreeSans 2560 0 0 0 VGND
port 16 nsew ground bidirectional
flabel metal5 s 1056 43676 40896 43996 0 FreeSans 2560 0 0 0 VGND
port 16 nsew ground bidirectional
flabel metal5 s 1056 48676 40896 48996 0 FreeSans 2560 0 0 0 VGND
port 16 nsew ground bidirectional
flabel metal5 s 1056 53676 40896 53996 0 FreeSans 2560 0 0 0 VGND
port 16 nsew ground bidirectional
flabel metal5 s 1056 58676 40896 58996 0 FreeSans 2560 0 0 0 VGND
port 16 nsew ground bidirectional
flabel metal5 s 1056 63676 40896 63996 0 FreeSans 2560 0 0 0 VGND
port 16 nsew ground bidirectional
flabel metal5 s 1056 68676 40896 68996 0 FreeSans 2560 0 0 0 VGND
port 16 nsew ground bidirectional
flabel metal4 s 1944 2128 2264 69680 0 FreeSans 1920 90 0 0 VPWR
port 17 nsew power bidirectional
flabel metal4 s 6944 2128 7264 69680 0 FreeSans 1920 90 0 0 VPWR
port 17 nsew power bidirectional
flabel metal4 s 11944 2128 12264 69680 0 FreeSans 1920 90 0 0 VPWR
port 17 nsew power bidirectional
flabel metal4 s 16944 2128 17264 69680 0 FreeSans 1920 90 0 0 VPWR
port 17 nsew power bidirectional
flabel metal4 s 21944 2128 22264 69680 0 FreeSans 1920 90 0 0 VPWR
port 17 nsew power bidirectional
flabel metal4 s 26944 2128 27264 69680 0 FreeSans 1920 90 0 0 VPWR
port 17 nsew power bidirectional
flabel metal4 s 31944 2128 32264 69680 0 FreeSans 1920 90 0 0 VPWR
port 17 nsew power bidirectional
flabel metal4 s 36944 2128 37264 69680 0 FreeSans 1920 90 0 0 VPWR
port 17 nsew power bidirectional
flabel metal5 s 1056 3016 40896 3336 0 FreeSans 2560 0 0 0 VPWR
port 17 nsew power bidirectional
flabel metal5 s 1056 8016 40896 8336 0 FreeSans 2560 0 0 0 VPWR
port 17 nsew power bidirectional
flabel metal5 s 1056 13016 40896 13336 0 FreeSans 2560 0 0 0 VPWR
port 17 nsew power bidirectional
flabel metal5 s 1056 18016 40896 18336 0 FreeSans 2560 0 0 0 VPWR
port 17 nsew power bidirectional
flabel metal5 s 1056 23016 40896 23336 0 FreeSans 2560 0 0 0 VPWR
port 17 nsew power bidirectional
flabel metal5 s 1056 28016 40896 28336 0 FreeSans 2560 0 0 0 VPWR
port 17 nsew power bidirectional
flabel metal5 s 1056 33016 40896 33336 0 FreeSans 2560 0 0 0 VPWR
port 17 nsew power bidirectional
flabel metal5 s 1056 38016 40896 38336 0 FreeSans 2560 0 0 0 VPWR
port 17 nsew power bidirectional
flabel metal5 s 1056 43016 40896 43336 0 FreeSans 2560 0 0 0 VPWR
port 17 nsew power bidirectional
flabel metal5 s 1056 48016 40896 48336 0 FreeSans 2560 0 0 0 VPWR
port 17 nsew power bidirectional
flabel metal5 s 1056 53016 40896 53336 0 FreeSans 2560 0 0 0 VPWR
port 17 nsew power bidirectional
flabel metal5 s 1056 58016 40896 58336 0 FreeSans 2560 0 0 0 VPWR
port 17 nsew power bidirectional
flabel metal5 s 1056 63016 40896 63336 0 FreeSans 2560 0 0 0 VPWR
port 17 nsew power bidirectional
flabel metal5 s 1056 68016 40896 68336 0 FreeSans 2560 0 0 0 VPWR
port 17 nsew power bidirectional
flabel metal2 s 34886 71200 34942 72000 0 FreeSans 224 90 0 0 opcode[0]
port 18 nsew signal input
flabel metal2 s 20902 71200 20958 72000 0 FreeSans 224 90 0 0 opcode[1]
port 19 nsew signal input
flabel metal2 s 6918 71200 6974 72000 0 FreeSans 224 90 0 0 opcode[2]
port 20 nsew signal input
flabel metal2 s 39302 0 39358 800 0 FreeSans 224 90 0 0 out[0]
port 21 nsew signal output
flabel metal2 s 34058 0 34114 800 0 FreeSans 224 90 0 0 out[1]
port 22 nsew signal output
flabel metal2 s 28814 0 28870 800 0 FreeSans 224 90 0 0 out[2]
port 23 nsew signal output
flabel metal2 s 23570 0 23626 800 0 FreeSans 224 90 0 0 out[3]
port 24 nsew signal output
flabel metal2 s 18326 0 18382 800 0 FreeSans 224 90 0 0 out[4]
port 25 nsew signal output
flabel metal2 s 13082 0 13138 800 0 FreeSans 224 90 0 0 out[5]
port 26 nsew signal output
flabel metal2 s 7838 0 7894 800 0 FreeSans 224 90 0 0 out[6]
port 27 nsew signal output
flabel metal2 s 2594 0 2650 800 0 FreeSans 224 90 0 0 out[7]
port 28 nsew signal output
rlabel metal1 20976 69632 20976 69632 0 VGND
rlabel metal1 20976 69088 20976 69088 0 VPWR
rlabel metal3 1050 67252 1050 67252 0 A[0]
rlabel metal3 751 58276 751 58276 0 A[1]
rlabel metal3 1050 49300 1050 49300 0 A[2]
rlabel metal3 751 40324 751 40324 0 A[3]
rlabel metal3 1050 31348 1050 31348 0 A[4]
rlabel metal3 751 22372 751 22372 0 A[5]
rlabel metal3 1050 13396 1050 13396 0 A[6]
rlabel metal3 751 4420 751 4420 0 A[7]
rlabel via2 40526 67235 40526 67235 0 B[0]
rlabel metal1 40158 59602 40158 59602 0 B[1]
rlabel metal2 40526 49555 40526 49555 0 B[2]
rlabel metal1 40572 40018 40572 40018 0 B[3]
rlabel via2 40526 31331 40526 31331 0 B[4]
rlabel metal2 40526 22491 40526 22491 0 B[5]
rlabel metal1 40158 13906 40158 13906 0 B[6]
rlabel metal2 40526 4301 40526 4301 0 B[7]
rlabel metal1 2162 16082 2162 16082 0 _000_
rlabel metal2 31786 43588 31786 43588 0 _001_
rlabel metal2 24702 26214 24702 26214 0 _002_
rlabel metal2 22448 29988 22448 29988 0 _003_
rlabel metal1 35236 57290 35236 57290 0 _004_
rlabel metal2 32338 39372 32338 39372 0 _005_
rlabel metal1 32476 38998 32476 38998 0 _006_
rlabel metal1 21160 42602 21160 42602 0 _007_
rlabel metal1 21574 41106 21574 41106 0 _008_
rlabel metal1 38548 52462 38548 52462 0 _009_
rlabel metal1 34316 52598 34316 52598 0 _010_
rlabel metal2 36846 52020 36846 52020 0 _011_
rlabel metal2 6854 57086 6854 57086 0 _012_
rlabel metal1 9890 43282 9890 43282 0 _013_
rlabel metal1 9062 62662 9062 62662 0 _014_
rlabel metal2 6670 33796 6670 33796 0 _015_
rlabel metal1 8372 32538 8372 32538 0 _016_
rlabel metal1 10212 43214 10212 43214 0 _017_
rlabel metal1 5750 16014 5750 16014 0 _018_
rlabel metal1 6394 4590 6394 4590 0 _019_
rlabel metal2 25024 20468 25024 20468 0 _020_
rlabel metal1 5474 4658 5474 4658 0 _021_
rlabel metal1 10304 41446 10304 41446 0 _022_
rlabel metal2 7130 54400 7130 54400 0 _023_
rlabel metal2 7866 21114 7866 21114 0 _024_
rlabel metal1 4922 55284 4922 55284 0 _025_
rlabel metal1 2530 33932 2530 33932 0 _026_
rlabel metal1 31418 28084 31418 28084 0 _027_
rlabel metal2 22310 58140 22310 58140 0 _028_
rlabel metal1 16698 12240 16698 12240 0 _029_
rlabel metal1 23322 58990 23322 58990 0 _030_
rlabel metal2 23690 58106 23690 58106 0 _031_
rlabel metal1 35420 21454 35420 21454 0 _032_
rlabel metal1 5750 55250 5750 55250 0 _033_
rlabel metal1 6072 55046 6072 55046 0 _034_
rlabel metal1 36386 49776 36386 49776 0 _035_
rlabel metal1 25300 25942 25300 25942 0 _036_
rlabel metal1 16790 9350 16790 9350 0 _037_
rlabel metal2 24794 31076 24794 31076 0 _038_
rlabel metal1 17572 9554 17572 9554 0 _039_
rlabel metal1 15617 7990 15617 7990 0 _040_
rlabel metal1 12880 67694 12880 67694 0 _041_
rlabel metal1 16054 7820 16054 7820 0 _042_
rlabel metal1 15962 32946 15962 32946 0 _043_
rlabel metal1 14122 9554 14122 9554 0 _044_
rlabel metal1 16146 7922 16146 7922 0 _045_
rlabel metal1 31648 25738 31648 25738 0 _046_
rlabel metal1 28888 17646 28888 17646 0 _047_
rlabel metal1 7222 4658 7222 4658 0 _048_
rlabel metal1 7314 4794 7314 4794 0 _049_
rlabel metal1 23782 27574 23782 27574 0 _050_
rlabel metal1 37720 17850 37720 17850 0 _051_
rlabel metal2 22402 18802 22402 18802 0 _052_
rlabel metal3 23529 59500 23529 59500 0 _053_
rlabel metal1 5750 66130 5750 66130 0 _054_
rlabel metal1 7222 16558 7222 16558 0 _055_
rlabel metal1 6302 52666 6302 52666 0 _056_
rlabel metal1 4416 53550 4416 53550 0 _057_
rlabel metal1 22678 60078 22678 60078 0 _058_
rlabel metal1 34224 20434 34224 20434 0 _059_
rlabel metal1 20654 23052 20654 23052 0 _060_
rlabel metal1 31326 30124 31326 30124 0 _061_
rlabel metal2 16560 31892 16560 31892 0 _062_
rlabel metal1 37950 4556 37950 4556 0 _063_
rlabel metal1 38042 4522 38042 4522 0 _064_
rlabel metal1 38410 4692 38410 4692 0 _065_
rlabel metal1 19918 4624 19918 4624 0 _066_
rlabel metal2 38594 4862 38594 4862 0 _067_
rlabel metal2 38410 14535 38410 14535 0 _068_
rlabel metal2 26082 24888 26082 24888 0 _069_
rlabel metal2 26174 24055 26174 24055 0 _070_
rlabel metal1 23736 2822 23736 2822 0 _071_
rlabel metal1 15502 22474 15502 22474 0 _072_
rlabel metal1 19182 62390 19182 62390 0 _073_
rlabel metal1 20240 62186 20240 62186 0 _074_
rlabel metal1 19366 62322 19366 62322 0 _075_
rlabel metal2 30958 29444 30958 29444 0 _076_
rlabel metal1 10948 48246 10948 48246 0 _077_
rlabel metal1 8694 20842 8694 20842 0 _078_
rlabel metal1 35788 29682 35788 29682 0 _079_
rlabel metal1 31648 6290 31648 6290 0 _080_
rlabel metal1 2898 65586 2898 65586 0 _081_
rlabel metal1 39238 14416 39238 14416 0 _082_
rlabel metal2 4186 36159 4186 36159 0 _083_
rlabel metal2 21850 49266 21850 49266 0 _084_
rlabel metal2 39514 30430 39514 30430 0 _085_
rlabel metal1 37490 14280 37490 14280 0 _086_
rlabel metal2 24702 19924 24702 19924 0 _087_
rlabel metal1 28612 41446 28612 41446 0 _088_
rlabel metal1 29118 14450 29118 14450 0 _089_
rlabel metal1 10212 52462 10212 52462 0 _090_
rlabel metal2 33074 40970 33074 40970 0 _091_
rlabel metal1 2530 50252 2530 50252 0 _092_
rlabel metal1 5014 44336 5014 44336 0 _093_
rlabel metal1 4738 44302 4738 44302 0 _094_
rlabel metal2 23598 29546 23598 29546 0 _095_
rlabel metal1 4738 51918 4738 51918 0 _096_
rlabel metal2 5106 43758 5106 43758 0 _097_
rlabel metal1 12098 43248 12098 43248 0 _098_
rlabel metal2 3082 13974 3082 13974 0 _099_
rlabel metal1 12328 43146 12328 43146 0 _100_
rlabel metal1 33580 19822 33580 19822 0 _101_
rlabel metal1 37628 15062 37628 15062 0 _102_
rlabel metal1 2484 61166 2484 61166 0 _103_
rlabel metal2 2346 59160 2346 59160 0 _104_
rlabel metal1 2714 10676 2714 10676 0 _105_
rlabel metal1 7176 19346 7176 19346 0 _106_
rlabel metal1 7498 19380 7498 19380 0 _107_
rlabel metal1 8694 19346 8694 19346 0 _108_
rlabel metal1 9246 3434 9246 3434 0 _109_
rlabel metal1 2714 50354 2714 50354 0 _110_
rlabel metal1 10028 61098 10028 61098 0 _111_
rlabel metal2 10994 7174 10994 7174 0 _112_
rlabel metal2 24610 38879 24610 38879 0 _113_
rlabel metal1 31832 60078 31832 60078 0 _114_
rlabel metal1 29578 60078 29578 60078 0 _115_
rlabel metal1 2530 65654 2530 65654 0 _116_
rlabel metal1 1794 20502 1794 20502 0 _117_
rlabel metal2 1702 22440 1702 22440 0 _118_
rlabel metal1 23230 12784 23230 12784 0 _119_
rlabel metal1 18906 44506 18906 44506 0 _120_
rlabel metal2 29118 58344 29118 58344 0 _121_
rlabel viali 19642 44847 19642 44847 0 _122_
rlabel metal1 23913 68374 23913 68374 0 _123_
rlabel metal1 24334 20230 24334 20230 0 _124_
rlabel metal1 33258 20298 33258 20298 0 _125_
rlabel metal1 37306 34510 37306 34510 0 _126_
rlabel metal1 37444 34714 37444 34714 0 _127_
rlabel metal1 23736 20502 23736 20502 0 _128_
rlabel metal1 24932 20570 24932 20570 0 _129_
rlabel metal2 34730 57936 34730 57936 0 _130_
rlabel metal1 30682 66538 30682 66538 0 _131_
rlabel metal1 18262 67082 18262 67082 0 _132_
rlabel metal2 33626 63563 33626 63563 0 _133_
rlabel metal2 36754 49606 36754 49606 0 _134_
rlabel metal1 17296 25738 17296 25738 0 _135_
rlabel metal1 26542 66572 26542 66572 0 _136_
rlabel metal2 26450 66300 26450 66300 0 _137_
rlabel metal1 17572 33558 17572 33558 0 _138_
rlabel metal2 26358 66164 26358 66164 0 _139_
rlabel metal2 20654 65552 20654 65552 0 _140_
rlabel metal1 6210 6256 6210 6256 0 _141_
rlabel metal1 23552 20978 23552 20978 0 _142_
rlabel metal1 30130 65926 30130 65926 0 _143_
rlabel metal1 26174 40970 26174 40970 0 _144_
rlabel metal2 3910 55488 3910 55488 0 _145_
rlabel metal1 15548 59466 15548 59466 0 _146_
rlabel metal2 13386 62492 13386 62492 0 _147_
rlabel metal1 14950 11152 14950 11152 0 _148_
rlabel metal2 20746 64226 20746 64226 0 _149_
rlabel metal2 24150 61438 24150 61438 0 _150_
rlabel metal1 38088 59058 38088 59058 0 _151_
rlabel metal3 21689 63580 21689 63580 0 _152_
rlabel metal1 34914 36176 34914 36176 0 _153_
rlabel metal2 24886 56134 24886 56134 0 _154_
rlabel metal2 3818 8143 3818 8143 0 _155_
rlabel metal2 10902 51476 10902 51476 0 _156_
rlabel metal1 19044 44370 19044 44370 0 _157_
rlabel metal1 38180 36822 38180 36822 0 _158_
rlabel metal2 39330 57256 39330 57256 0 _159_
rlabel metal1 5566 52530 5566 52530 0 _160_
rlabel metal2 35282 43282 35282 43282 0 _161_
rlabel metal1 30958 14382 30958 14382 0 _162_
rlabel metal1 30452 14314 30452 14314 0 _163_
rlabel metal2 20654 48450 20654 48450 0 _164_
rlabel metal1 29808 18258 29808 18258 0 _165_
rlabel metal1 28014 18190 28014 18190 0 _166_
rlabel metal1 3036 50422 3036 50422 0 _167_
rlabel metal1 17848 6154 17848 6154 0 _168_
rlabel metal1 5934 6324 5934 6324 0 _169_
rlabel metal1 12098 50218 12098 50218 0 _170_
rlabel metal1 32522 62322 32522 62322 0 _171_
rlabel metal1 13294 50728 13294 50728 0 _172_
rlabel metal1 29532 66470 29532 66470 0 _173_
rlabel metal2 13570 37706 13570 37706 0 _174_
rlabel metal1 14214 3502 14214 3502 0 _175_
rlabel metal1 4968 45458 4968 45458 0 _176_
rlabel metal1 24656 38522 24656 38522 0 _177_
rlabel metal2 13754 41820 13754 41820 0 _178_
rlabel metal1 13662 33082 13662 33082 0 _179_
rlabel metal1 5566 59058 5566 59058 0 _180_
rlabel metal1 13202 35088 13202 35088 0 _181_
rlabel metal1 4600 61098 4600 61098 0 _182_
rlabel metal1 16698 43214 16698 43214 0 _183_
rlabel metal2 27462 23919 27462 23919 0 _184_
rlabel metal1 38134 48722 38134 48722 0 _185_
rlabel metal1 19642 44948 19642 44948 0 _186_
rlabel metal1 8234 3604 8234 3604 0 _187_
rlabel metal1 38042 67694 38042 67694 0 _188_
rlabel metal2 19642 43520 19642 43520 0 _189_
rlabel metal1 3772 9010 3772 9010 0 _190_
rlabel metal2 1886 10047 1886 10047 0 _191_
rlabel via2 38042 67813 38042 67813 0 _192_
rlabel metal1 19167 62866 19167 62866 0 _193_
rlabel metal1 21896 50830 21896 50830 0 _194_
rlabel metal1 2990 16218 2990 16218 0 _195_
rlabel metal2 5566 60894 5566 60894 0 _196_
rlabel metal1 37996 37978 37996 37978 0 _197_
rlabel metal2 6808 5780 6808 5780 0 _198_
rlabel metal1 27876 63206 27876 63206 0 _199_
rlabel metal1 37030 7922 37030 7922 0 _200_
rlabel metal1 17250 48654 17250 48654 0 _201_
rlabel metal1 17204 62798 17204 62798 0 _202_
rlabel metal1 3266 21012 3266 21012 0 _203_
rlabel metal1 37490 19822 37490 19822 0 _204_
rlabel metal1 33488 42194 33488 42194 0 _205_
rlabel metal1 16422 28492 16422 28492 0 _206_
rlabel metal1 16146 28526 16146 28526 0 _207_
rlabel metal1 37950 19890 37950 19890 0 _208_
rlabel metal1 24794 20536 24794 20536 0 _209_
rlabel metal1 14858 38182 14858 38182 0 _210_
rlabel metal1 4094 20842 4094 20842 0 _211_
rlabel metal1 32292 40494 32292 40494 0 _212_
rlabel metal1 38916 14042 38916 14042 0 _213_
rlabel metal1 21160 59942 21160 59942 0 _214_
rlabel metal1 21298 42568 21298 42568 0 _215_
rlabel metal1 3910 20774 3910 20774 0 _216_
rlabel metal1 1426 61234 1426 61234 0 _217_
rlabel metal1 20746 42704 20746 42704 0 _218_
rlabel metal1 6440 44846 6440 44846 0 _219_
rlabel metal1 15456 50830 15456 50830 0 _220_
rlabel metal1 16698 42670 16698 42670 0 _221_
rlabel metal2 6762 47532 6762 47532 0 _222_
rlabel metal1 32522 44812 32522 44812 0 _223_
rlabel metal1 9614 62866 9614 62866 0 _224_
rlabel metal2 32338 43112 32338 43112 0 _225_
rlabel metal1 13800 55726 13800 55726 0 _226_
rlabel metal1 36110 33048 36110 33048 0 _227_
rlabel metal1 26910 8942 26910 8942 0 _228_
rlabel metal1 18423 64294 18423 64294 0 _229_
rlabel metal1 37766 4624 37766 4624 0 _230_
rlabel metal1 3634 6358 3634 6358 0 _231_
rlabel metal1 1978 30702 1978 30702 0 _232_
rlabel metal1 2024 40494 2024 40494 0 _233_
rlabel metal3 20447 63580 20447 63580 0 _234_
rlabel metal1 22540 64294 22540 64294 0 _235_
rlabel metal1 2438 30770 2438 30770 0 _236_
rlabel metal1 14582 54026 14582 54026 0 _237_
rlabel metal1 19366 6698 19366 6698 0 _238_
rlabel metal2 7866 64634 7866 64634 0 _239_
rlabel metal1 38962 60622 38962 60622 0 _240_
rlabel metal1 37030 32878 37030 32878 0 _241_
rlabel metal1 37306 32980 37306 32980 0 _242_
rlabel metal2 16698 7310 16698 7310 0 _243_
rlabel metal2 38778 56814 38778 56814 0 _244_
rlabel metal1 17480 6358 17480 6358 0 _245_
rlabel metal2 10994 56882 10994 56882 0 _246_
rlabel metal2 39146 60384 39146 60384 0 _247_
rlabel metal1 20654 42636 20654 42636 0 net1
rlabel metal1 19044 4590 19044 4590 0 net10
rlabel metal2 22310 20060 22310 20060 0 net11
rlabel metal1 37766 40562 37766 40562 0 net12
rlabel metal2 27554 24157 27554 24157 0 net13
rlabel metal2 26174 22916 26174 22916 0 net14
rlabel metal1 37950 36720 37950 36720 0 net15
rlabel metal1 18906 44404 18906 44404 0 net16
rlabel metal1 4370 59058 4370 59058 0 net17
rlabel metal1 4094 19890 4094 19890 0 net18
rlabel metal2 32890 42228 32890 42228 0 net19
rlabel metal2 6762 58786 6762 58786 0 net2
rlabel metal1 39238 2414 39238 2414 0 net20
rlabel metal1 18354 61574 18354 61574 0 net21
rlabel via2 28658 2363 28658 2363 0 net22
rlabel metal1 23506 2414 23506 2414 0 net23
rlabel metal2 34638 5406 34638 5406 0 net24
rlabel metal2 24610 11458 24610 11458 0 net25
rlabel metal1 9154 2414 9154 2414 0 net26
rlabel metal1 2990 2448 2990 2448 0 net27
rlabel metal1 3450 20434 3450 20434 0 net28
rlabel metal1 11454 44438 11454 44438 0 net29
rlabel metal2 7314 51646 7314 51646 0 net3
rlabel metal1 16284 33014 16284 33014 0 net30
rlabel metal1 37076 63954 37076 63954 0 net31
rlabel metal1 4370 66096 4370 66096 0 net32
rlabel metal1 21298 38964 21298 38964 0 net33
rlabel metal2 31924 29036 31924 29036 0 net34
rlabel metal2 30130 66130 30130 66130 0 net35
rlabel metal2 29670 63376 29670 63376 0 net36
rlabel metal1 32200 29546 32200 29546 0 net37
rlabel metal2 30406 28764 30406 28764 0 net38
rlabel metal1 24472 28594 24472 28594 0 net39
rlabel metal2 4370 4794 4370 4794 0 net4
rlabel metal2 20746 26622 20746 26622 0 net40
rlabel metal1 32798 62254 32798 62254 0 net41
rlabel metal1 33166 39508 33166 39508 0 net42
rlabel metal2 8510 4182 8510 4182 0 net43
rlabel metal1 35052 37230 35052 37230 0 net44
rlabel metal2 38042 36924 38042 36924 0 net45
rlabel metal1 7360 59126 7360 59126 0 net46
rlabel metal1 19964 7378 19964 7378 0 net47
rlabel metal2 23414 10948 23414 10948 0 net48
rlabel metal1 17158 31926 17158 31926 0 net49
rlabel metal1 2070 25942 2070 25942 0 net5
rlabel metal1 38502 32878 38502 32878 0 net50
rlabel metal1 38686 32980 38686 32980 0 net51
rlabel metal1 7130 21012 7130 21012 0 net52
rlabel metal1 7498 20944 7498 20944 0 net53
rlabel metal1 7820 19890 7820 19890 0 net54
rlabel metal1 5428 4522 5428 4522 0 net55
rlabel metal1 19504 18598 19504 18598 0 net56
rlabel metal1 40250 57392 40250 57392 0 net57
rlabel metal1 32292 39270 32292 39270 0 net58
rlabel metal2 28014 37468 28014 37468 0 net59
rlabel metal1 21022 7446 21022 7446 0 net6
rlabel metal1 38548 15062 38548 15062 0 net60
rlabel metal1 4462 4488 4462 4488 0 net61
rlabel metal2 35834 52292 35834 52292 0 net62
rlabel metal1 39008 57426 39008 57426 0 net63
rlabel metal2 23138 40698 23138 40698 0 net64
rlabel metal1 6762 45492 6762 45492 0 net65
rlabel metal1 4445 16082 4445 16082 0 net66
rlabel metal2 4830 60894 4830 60894 0 net7
rlabel metal1 2990 4658 2990 4658 0 net8
rlabel metal1 5566 60520 5566 60520 0 net9
rlabel metal2 35006 70397 35006 70397 0 opcode[0]
rlabel metal1 21436 69394 21436 69394 0 opcode[1]
rlabel metal2 7130 70363 7130 70363 0 opcode[2]
rlabel metal2 39330 1520 39330 1520 0 out[0]
rlabel metal2 34086 1520 34086 1520 0 out[1]
rlabel metal2 28842 1520 28842 1520 0 out[2]
rlabel metal2 23598 1520 23598 1520 0 out[3]
rlabel metal2 18354 1520 18354 1520 0 out[4]
rlabel metal2 13110 1520 13110 1520 0 out[5]
rlabel metal2 7866 959 7866 959 0 out[6]
rlabel metal2 2622 959 2622 959 0 out[7]
<< properties >>
string FIXED_BBOX 0 0 42000 72000
<< end >>

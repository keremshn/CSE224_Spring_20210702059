magic
tech sky130A
magscale 1 2
timestamp 1746359155
<< nwell >>
rect 1066 2159 40886 69649
<< obsli1 >>
rect 1104 2159 40848 69649
<< obsm1 >>
rect 842 2128 40926 69680
<< metal2 >>
rect 6918 71200 6974 72000
rect 20902 71200 20958 72000
rect 34886 71200 34942 72000
rect 2594 0 2650 800
rect 7838 0 7894 800
rect 13082 0 13138 800
rect 18326 0 18382 800
rect 23570 0 23626 800
rect 28814 0 28870 800
rect 34058 0 34114 800
rect 39302 0 39358 800
<< obsm2 >>
rect 846 71144 6862 71346
rect 7030 71144 20846 71346
rect 21014 71144 34830 71346
rect 34998 71144 40922 71346
rect 846 856 40922 71144
rect 846 800 2538 856
rect 2706 800 7782 856
rect 7950 800 13026 856
rect 13194 800 18270 856
rect 18438 800 23514 856
rect 23682 800 28758 856
rect 28926 800 34002 856
rect 34170 800 39246 856
rect 39414 800 40922 856
<< metal3 >>
rect 0 67192 800 67312
rect 41200 67192 42000 67312
rect 0 58216 800 58336
rect 41200 58216 42000 58336
rect 0 49240 800 49360
rect 41200 49240 42000 49360
rect 0 40264 800 40384
rect 41200 40264 42000 40384
rect 0 31288 800 31408
rect 41200 31288 42000 31408
rect 0 22312 800 22432
rect 41200 22312 42000 22432
rect 0 13336 800 13456
rect 41200 13336 42000 13456
rect 0 4360 800 4480
rect 41200 4360 42000 4480
<< obsm3 >>
rect 798 67392 41200 69665
rect 880 67112 41120 67392
rect 798 58416 41200 67112
rect 880 58136 41120 58416
rect 798 49440 41200 58136
rect 880 49160 41120 49440
rect 798 40464 41200 49160
rect 880 40184 41120 40464
rect 798 31488 41200 40184
rect 880 31208 41120 31488
rect 798 22512 41200 31208
rect 880 22232 41120 22512
rect 798 13536 41200 22232
rect 880 13256 41120 13536
rect 798 4560 41200 13256
rect 880 4280 41120 4560
rect 798 2143 41200 4280
<< metal4 >>
rect 1944 2128 2264 69680
rect 2604 2128 2924 69680
rect 6944 2128 7264 69680
rect 7604 2128 7924 69680
rect 11944 2128 12264 69680
rect 12604 2128 12924 69680
rect 16944 2128 17264 69680
rect 17604 2128 17924 69680
rect 21944 2128 22264 69680
rect 22604 2128 22924 69680
rect 26944 2128 27264 69680
rect 27604 2128 27924 69680
rect 31944 2128 32264 69680
rect 32604 2128 32924 69680
rect 36944 2128 37264 69680
rect 37604 2128 37924 69680
<< obsm4 >>
rect 3371 2347 6864 67829
rect 7344 2347 7524 67829
rect 8004 2347 11864 67829
rect 12344 2347 12524 67829
rect 13004 2347 16864 67829
rect 17344 2347 17524 67829
rect 18004 2347 21864 67829
rect 22344 2347 22524 67829
rect 23004 2347 26864 67829
rect 27344 2347 27524 67829
rect 28004 2347 31864 67829
rect 32344 2347 32524 67829
rect 33004 2347 34901 67829
<< metal5 >>
rect 1056 68676 40896 68996
rect 1056 68016 40896 68336
rect 1056 63676 40896 63996
rect 1056 63016 40896 63336
rect 1056 58676 40896 58996
rect 1056 58016 40896 58336
rect 1056 53676 40896 53996
rect 1056 53016 40896 53336
rect 1056 48676 40896 48996
rect 1056 48016 40896 48336
rect 1056 43676 40896 43996
rect 1056 43016 40896 43336
rect 1056 38676 40896 38996
rect 1056 38016 40896 38336
rect 1056 33676 40896 33996
rect 1056 33016 40896 33336
rect 1056 28676 40896 28996
rect 1056 28016 40896 28336
rect 1056 23676 40896 23996
rect 1056 23016 40896 23336
rect 1056 18676 40896 18996
rect 1056 18016 40896 18336
rect 1056 13676 40896 13996
rect 1056 13016 40896 13336
rect 1056 8676 40896 8996
rect 1056 8016 40896 8336
rect 1056 3676 40896 3996
rect 1056 3016 40896 3336
<< labels >>
rlabel metal3 s 0 67192 800 67312 6 A[0]
port 1 nsew signal input
rlabel metal3 s 0 58216 800 58336 6 A[1]
port 2 nsew signal input
rlabel metal3 s 0 49240 800 49360 6 A[2]
port 3 nsew signal input
rlabel metal3 s 0 40264 800 40384 6 A[3]
port 4 nsew signal input
rlabel metal3 s 0 31288 800 31408 6 A[4]
port 5 nsew signal input
rlabel metal3 s 0 22312 800 22432 6 A[5]
port 6 nsew signal input
rlabel metal3 s 0 13336 800 13456 6 A[6]
port 7 nsew signal input
rlabel metal3 s 0 4360 800 4480 6 A[7]
port 8 nsew signal input
rlabel metal3 s 41200 67192 42000 67312 6 B[0]
port 9 nsew signal input
rlabel metal3 s 41200 58216 42000 58336 6 B[1]
port 10 nsew signal input
rlabel metal3 s 41200 49240 42000 49360 6 B[2]
port 11 nsew signal input
rlabel metal3 s 41200 40264 42000 40384 6 B[3]
port 12 nsew signal input
rlabel metal3 s 41200 31288 42000 31408 6 B[4]
port 13 nsew signal input
rlabel metal3 s 41200 22312 42000 22432 6 B[5]
port 14 nsew signal input
rlabel metal3 s 41200 13336 42000 13456 6 B[6]
port 15 nsew signal input
rlabel metal3 s 41200 4360 42000 4480 6 B[7]
port 16 nsew signal input
rlabel metal4 s 2604 2128 2924 69680 6 VGND
port 17 nsew ground bidirectional
rlabel metal4 s 7604 2128 7924 69680 6 VGND
port 17 nsew ground bidirectional
rlabel metal4 s 12604 2128 12924 69680 6 VGND
port 17 nsew ground bidirectional
rlabel metal4 s 17604 2128 17924 69680 6 VGND
port 17 nsew ground bidirectional
rlabel metal4 s 22604 2128 22924 69680 6 VGND
port 17 nsew ground bidirectional
rlabel metal4 s 27604 2128 27924 69680 6 VGND
port 17 nsew ground bidirectional
rlabel metal4 s 32604 2128 32924 69680 6 VGND
port 17 nsew ground bidirectional
rlabel metal4 s 37604 2128 37924 69680 6 VGND
port 17 nsew ground bidirectional
rlabel metal5 s 1056 3676 40896 3996 6 VGND
port 17 nsew ground bidirectional
rlabel metal5 s 1056 8676 40896 8996 6 VGND
port 17 nsew ground bidirectional
rlabel metal5 s 1056 13676 40896 13996 6 VGND
port 17 nsew ground bidirectional
rlabel metal5 s 1056 18676 40896 18996 6 VGND
port 17 nsew ground bidirectional
rlabel metal5 s 1056 23676 40896 23996 6 VGND
port 17 nsew ground bidirectional
rlabel metal5 s 1056 28676 40896 28996 6 VGND
port 17 nsew ground bidirectional
rlabel metal5 s 1056 33676 40896 33996 6 VGND
port 17 nsew ground bidirectional
rlabel metal5 s 1056 38676 40896 38996 6 VGND
port 17 nsew ground bidirectional
rlabel metal5 s 1056 43676 40896 43996 6 VGND
port 17 nsew ground bidirectional
rlabel metal5 s 1056 48676 40896 48996 6 VGND
port 17 nsew ground bidirectional
rlabel metal5 s 1056 53676 40896 53996 6 VGND
port 17 nsew ground bidirectional
rlabel metal5 s 1056 58676 40896 58996 6 VGND
port 17 nsew ground bidirectional
rlabel metal5 s 1056 63676 40896 63996 6 VGND
port 17 nsew ground bidirectional
rlabel metal5 s 1056 68676 40896 68996 6 VGND
port 17 nsew ground bidirectional
rlabel metal4 s 1944 2128 2264 69680 6 VPWR
port 18 nsew power bidirectional
rlabel metal4 s 6944 2128 7264 69680 6 VPWR
port 18 nsew power bidirectional
rlabel metal4 s 11944 2128 12264 69680 6 VPWR
port 18 nsew power bidirectional
rlabel metal4 s 16944 2128 17264 69680 6 VPWR
port 18 nsew power bidirectional
rlabel metal4 s 21944 2128 22264 69680 6 VPWR
port 18 nsew power bidirectional
rlabel metal4 s 26944 2128 27264 69680 6 VPWR
port 18 nsew power bidirectional
rlabel metal4 s 31944 2128 32264 69680 6 VPWR
port 18 nsew power bidirectional
rlabel metal4 s 36944 2128 37264 69680 6 VPWR
port 18 nsew power bidirectional
rlabel metal5 s 1056 3016 40896 3336 6 VPWR
port 18 nsew power bidirectional
rlabel metal5 s 1056 8016 40896 8336 6 VPWR
port 18 nsew power bidirectional
rlabel metal5 s 1056 13016 40896 13336 6 VPWR
port 18 nsew power bidirectional
rlabel metal5 s 1056 18016 40896 18336 6 VPWR
port 18 nsew power bidirectional
rlabel metal5 s 1056 23016 40896 23336 6 VPWR
port 18 nsew power bidirectional
rlabel metal5 s 1056 28016 40896 28336 6 VPWR
port 18 nsew power bidirectional
rlabel metal5 s 1056 33016 40896 33336 6 VPWR
port 18 nsew power bidirectional
rlabel metal5 s 1056 38016 40896 38336 6 VPWR
port 18 nsew power bidirectional
rlabel metal5 s 1056 43016 40896 43336 6 VPWR
port 18 nsew power bidirectional
rlabel metal5 s 1056 48016 40896 48336 6 VPWR
port 18 nsew power bidirectional
rlabel metal5 s 1056 53016 40896 53336 6 VPWR
port 18 nsew power bidirectional
rlabel metal5 s 1056 58016 40896 58336 6 VPWR
port 18 nsew power bidirectional
rlabel metal5 s 1056 63016 40896 63336 6 VPWR
port 18 nsew power bidirectional
rlabel metal5 s 1056 68016 40896 68336 6 VPWR
port 18 nsew power bidirectional
rlabel metal2 s 34886 71200 34942 72000 6 opcode[0]
port 19 nsew signal input
rlabel metal2 s 20902 71200 20958 72000 6 opcode[1]
port 20 nsew signal input
rlabel metal2 s 6918 71200 6974 72000 6 opcode[2]
port 21 nsew signal input
rlabel metal2 s 39302 0 39358 800 6 out[0]
port 22 nsew signal output
rlabel metal2 s 34058 0 34114 800 6 out[1]
port 23 nsew signal output
rlabel metal2 s 28814 0 28870 800 6 out[2]
port 24 nsew signal output
rlabel metal2 s 23570 0 23626 800 6 out[3]
port 25 nsew signal output
rlabel metal2 s 18326 0 18382 800 6 out[4]
port 26 nsew signal output
rlabel metal2 s 13082 0 13138 800 6 out[5]
port 27 nsew signal output
rlabel metal2 s 7838 0 7894 800 6 out[6]
port 28 nsew signal output
rlabel metal2 s 2594 0 2650 800 6 out[7]
port 29 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 42000 72000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 3235834
string GDS_FILE /openlane/designs/ALU/runs/RUN_2025.05.04_11.45.11/results/signoff/ALU.magic.gds
string GDS_START 729516
<< end >>


// This is the unpowered netlist.
module ALU (A,
    B,
    opcode,
    out);
 input [7:0] A;
 input [7:0] B;
 input [2:0] opcode;
 output [7:0] out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire net1;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net7;
 wire net8;
 wire net9;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_006_));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(_191_));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(_213_));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(_213_));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(_213_));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(_213_));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(_240_));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(_244_));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(_245_));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(_247_));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_021_));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(_041_));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_082_));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(_141_));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(_240_));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_36 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_094_));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(_095_));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(_103_));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(_116_));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(_183_));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(_189_));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_10 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_34 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_16 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_224 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_225 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_102_Left_226 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_102_Right_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_103_Left_227 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_103_Right_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_104_Left_228 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_104_Right_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_105_Left_229 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_105_Right_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_106_Left_230 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_106_Right_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_107_Left_231 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_107_Right_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_108_Left_232 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_108_Right_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_109_Left_233 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_109_Right_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_110_Left_234 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_110_Right_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_111_Left_235 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_111_Right_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_112_Left_236 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_112_Right_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_113_Left_237 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_113_Right_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_114_Left_238 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_114_Right_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_115_Left_239 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_115_Right_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_116_Left_240 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_116_Right_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_117_Left_241 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_117_Right_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_118_Left_242 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_118_Right_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_119_Left_243 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_119_Right_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_120_Left_244 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_120_Right_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_121_Left_245 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_121_Right_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_122_Left_246 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_122_Right_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_123_Left_247 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_123_Right_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_203 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_204 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_205 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_206 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_207 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_208 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_209 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_210 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_211 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_212 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_213 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_214 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_215 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_216 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_217 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_218 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_219 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_220 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_221 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_222 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_223 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_329 ();
 sky130_fd_sc_hd__buf_8 _248_ (.A(net1),
    .X(_176_));
 sky130_fd_sc_hd__or2_4 _249_ (.A(net17),
    .B(net18),
    .X(_180_));
 sky130_fd_sc_hd__or2_2 _250_ (.A(net19),
    .B(_180_),
    .X(_181_));
 sky130_fd_sc_hd__clkbuf_16 _251_ (.A(net9),
    .X(_182_));
 sky130_fd_sc_hd__buf_12 _252_ (.A(_182_),
    .X(_183_));
 sky130_fd_sc_hd__or2_1 _253_ (.A(_176_),
    .B(_183_),
    .X(_184_));
 sky130_fd_sc_hd__nand2_4 _254_ (.A(net17),
    .B(net18),
    .Y(_185_));
 sky130_fd_sc_hd__inv_4 _255_ (.A(net19),
    .Y(_186_));
 sky130_fd_sc_hd__nand2_8 _256_ (.A(net17),
    .B(_186_),
    .Y(_187_));
 sky130_fd_sc_hd__nand3_4 _257_ (.A(_176_),
    .B(_183_),
    .C(_187_),
    .Y(_188_));
 sky130_fd_sc_hd__nor2_8 _258_ (.A(_186_),
    .B(_180_),
    .Y(_189_));
 sky130_fd_sc_hd__nor2_4 _259_ (.A(net19),
    .B(_185_),
    .Y(_190_));
 sky130_fd_sc_hd__o211a_4 _260_ (.A1(_189_),
    .A2(_190_),
    .B1(_176_),
    .C1(_183_),
    .X(_191_));
 sky130_fd_sc_hd__a31o_2 _261_ (.A1(_180_),
    .A2(_185_),
    .A3(_188_),
    .B1(_191_),
    .X(_192_));
 sky130_fd_sc_hd__a2bb2o_2 _262_ (.A1_N(_176_),
    .A2_N(_181_),
    .B1(_184_),
    .B2(_192_),
    .X(net20));
 sky130_fd_sc_hd__buf_8 _263_ (.A(net44),
    .X(_193_));
 sky130_fd_sc_hd__nor2_2 _264_ (.A(net19),
    .B(_180_),
    .Y(_194_));
 sky130_fd_sc_hd__clkbuf_8 _265_ (.A(_194_),
    .X(_195_));
 sky130_fd_sc_hd__buf_12 _266_ (.A(net10),
    .X(_196_));
 sky130_fd_sc_hd__clkbuf_8 _267_ (.A(_196_),
    .X(_197_));
 sky130_fd_sc_hd__nor2_8 _268_ (.A(net18),
    .B(_187_),
    .Y(_198_));
 sky130_fd_sc_hd__or3b_2 _269_ (.A(net17),
    .B(net19),
    .C_N(net18),
    .X(_199_));
 sky130_fd_sc_hd__clkbuf_8 _270_ (.A(_199_),
    .X(_200_));
 sky130_fd_sc_hd__a21oi_2 _271_ (.A1(_193_),
    .A2(_197_),
    .B1(_200_),
    .Y(_201_));
 sky130_fd_sc_hd__o22a_1 _272_ (.A1(_193_),
    .A2(_197_),
    .B1(_198_),
    .B2(_201_),
    .X(_202_));
 sky130_fd_sc_hd__and3_4 _273_ (.A(net19),
    .B(_180_),
    .C(_185_),
    .X(_203_));
 sky130_fd_sc_hd__or2b_2 _274_ (.A(net1),
    .B_N(_183_),
    .X(_204_));
 sky130_fd_sc_hd__nand3b_4 _275_ (.A_N(net17),
    .B(net18),
    .C(net19),
    .Y(_205_));
 sky130_fd_sc_hd__a21oi_2 _276_ (.A1(_183_),
    .A2(net32),
    .B1(_197_),
    .Y(_206_));
 sky130_fd_sc_hd__and3_1 _277_ (.A(net63),
    .B(_197_),
    .C(_205_),
    .X(_207_));
 sky130_fd_sc_hd__o21a_2 _278_ (.A1(_206_),
    .A2(_207_),
    .B1(_193_),
    .X(_208_));
 sky130_fd_sc_hd__or3_4 _279_ (.A(_193_),
    .B(_206_),
    .C(_207_),
    .X(_209_));
 sky130_fd_sc_hd__or2b_1 _280_ (.A(_208_),
    .B_N(_209_),
    .X(_210_));
 sky130_fd_sc_hd__xnor2_1 _281_ (.A(_204_),
    .B(_210_),
    .Y(_211_));
 sky130_fd_sc_hd__and4_2 _282_ (.A(_176_),
    .B(_183_),
    .C(_193_),
    .D(_197_),
    .X(_212_));
 sky130_fd_sc_hd__a22o_2 _283_ (.A1(_183_),
    .A2(_193_),
    .B1(_197_),
    .B2(_176_),
    .X(_213_));
 sky130_fd_sc_hd__and3b_1 _284_ (.A_N(_212_),
    .B(_189_),
    .C(_213_),
    .X(_214_));
 sky130_fd_sc_hd__a31o_2 _285_ (.A1(_193_),
    .A2(_197_),
    .A3(_190_),
    .B1(_214_),
    .X(_215_));
 sky130_fd_sc_hd__a211o_2 _286_ (.A1(_203_),
    .A2(_211_),
    .B1(_215_),
    .C1(_195_),
    .X(_216_));
 sky130_fd_sc_hd__o2bb2a_2 _287_ (.A1_N(_193_),
    .A2_N(_195_),
    .B1(_202_),
    .B2(_216_),
    .X(net21));
 sky130_fd_sc_hd__buf_8 _288_ (.A(net54),
    .X(_217_));
 sky130_fd_sc_hd__buf_12 _289_ (.A(net11),
    .X(_218_));
 sky130_fd_sc_hd__nand2_2 _290_ (.A(_176_),
    .B(net65),
    .Y(_219_));
 sky130_fd_sc_hd__and3_1 _291_ (.A(_193_),
    .B(_197_),
    .C(_217_),
    .X(_220_));
 sky130_fd_sc_hd__a22o_1 _292_ (.A1(net2),
    .A2(net47),
    .B1(_217_),
    .B2(net63),
    .X(_221_));
 sky130_fd_sc_hd__a21bo_2 _293_ (.A1(_183_),
    .A2(_220_),
    .B1_N(_221_),
    .X(_222_));
 sky130_fd_sc_hd__xor2_4 _294_ (.A(_219_),
    .B(_222_),
    .X(_223_));
 sky130_fd_sc_hd__and2_4 _295_ (.A(_212_),
    .B(_223_),
    .X(_224_));
 sky130_fd_sc_hd__o21ai_2 _296_ (.A1(_212_),
    .A2(_223_),
    .B1(_189_),
    .Y(_225_));
 sky130_fd_sc_hd__nor2_1 _297_ (.A(_224_),
    .B(_225_),
    .Y(_226_));
 sky130_fd_sc_hd__o21a_4 _298_ (.A1(_183_),
    .A2(_197_),
    .B1(net50),
    .X(_227_));
 sky130_fd_sc_hd__xnor2_4 _299_ (.A(_218_),
    .B(_227_),
    .Y(_228_));
 sky130_fd_sc_hd__xor2_4 _300_ (.A(_217_),
    .B(_228_),
    .X(_229_));
 sky130_fd_sc_hd__a21o_4 _301_ (.A1(_204_),
    .A2(_209_),
    .B1(_208_),
    .X(_230_));
 sky130_fd_sc_hd__nand2_2 _302_ (.A(_229_),
    .B(_230_),
    .Y(_231_));
 sky130_fd_sc_hd__o21a_2 _303_ (.A1(_229_),
    .A2(_230_),
    .B1(_203_),
    .X(_232_));
 sky130_fd_sc_hd__nand2_8 _304_ (.A(net54),
    .B(net11),
    .Y(_233_));
 sky130_fd_sc_hd__and2b_2 _305_ (.A_N(_200_),
    .B(_233_),
    .X(_234_));
 sky130_fd_sc_hd__o22a_1 _306_ (.A1(_217_),
    .A2(net65),
    .B1(_198_),
    .B2(_234_),
    .X(_235_));
 sky130_fd_sc_hd__a31o_2 _307_ (.A1(_217_),
    .A2(net65),
    .A3(_190_),
    .B1(_235_),
    .X(_236_));
 sky130_fd_sc_hd__a211o_1 _308_ (.A1(_231_),
    .A2(_232_),
    .B1(_236_),
    .C1(_195_),
    .X(_237_));
 sky130_fd_sc_hd__o2bb2a_2 _309_ (.A1_N(_217_),
    .A2_N(_195_),
    .B1(_226_),
    .B2(_237_),
    .X(net22));
 sky130_fd_sc_hd__buf_12 _310_ (.A(net4),
    .X(_238_));
 sky130_fd_sc_hd__and2_1 _311_ (.A(_217_),
    .B(_228_),
    .X(_239_));
 sky130_fd_sc_hd__a21o_4 _312_ (.A1(_229_),
    .A2(_230_),
    .B1(_239_),
    .X(_240_));
 sky130_fd_sc_hd__buf_8 _313_ (.A(net62),
    .X(_241_));
 sky130_fd_sc_hd__a211oi_4 _314_ (.A1(net65),
    .A2(net51),
    .B1(_227_),
    .C1(_241_),
    .Y(_242_));
 sky130_fd_sc_hd__o311a_4 _315_ (.A1(_183_),
    .A2(_197_),
    .A3(net65),
    .B1(_241_),
    .C1(net32),
    .X(_243_));
 sky130_fd_sc_hd__o21ai_4 _316_ (.A1(net30),
    .A2(_243_),
    .B1(net66),
    .Y(_244_));
 sky130_fd_sc_hd__or3_4 _317_ (.A(_238_),
    .B(_242_),
    .C(_243_),
    .X(_245_));
 sky130_fd_sc_hd__and3_2 _318_ (.A(_240_),
    .B(_244_),
    .C(_245_),
    .X(_246_));
 sky130_fd_sc_hd__a21o_1 _319_ (.A1(_244_),
    .A2(_245_),
    .B1(_240_),
    .X(_247_));
 sky130_fd_sc_hd__and3b_2 _320_ (.A_N(_246_),
    .B(_247_),
    .C(_203_),
    .X(_000_));
 sky130_fd_sc_hd__nand2_4 _321_ (.A(_176_),
    .B(_241_),
    .Y(_001_));
 sky130_fd_sc_hd__nand2_4 _322_ (.A(net46),
    .B(_218_),
    .Y(_002_));
 sky130_fd_sc_hd__and4_4 _323_ (.A(net9),
    .B(net10),
    .C(net56),
    .D(net4),
    .X(_003_));
 sky130_fd_sc_hd__a22oi_4 _324_ (.A1(_196_),
    .A2(net57),
    .B1(_238_),
    .B2(net63),
    .Y(_004_));
 sky130_fd_sc_hd__or3_4 _325_ (.A(_002_),
    .B(_003_),
    .C(net39),
    .X(_005_));
 sky130_fd_sc_hd__o21ai_4 _326_ (.A1(net40),
    .A2(_003_),
    .B1(_002_),
    .Y(_006_));
 sky130_fd_sc_hd__and4_4 _327_ (.A(net63),
    .B(net43),
    .C(net47),
    .D(_217_),
    .X(_007_));
 sky130_fd_sc_hd__a31o_4 _328_ (.A1(net1),
    .A2(_218_),
    .A3(_221_),
    .B1(_007_),
    .X(_008_));
 sky130_fd_sc_hd__and3_1 _329_ (.A(_006_),
    .B(_005_),
    .C(_008_),
    .X(_009_));
 sky130_fd_sc_hd__a21o_4 _330_ (.A1(_005_),
    .A2(_006_),
    .B1(_008_),
    .X(_010_));
 sky130_fd_sc_hd__and2b_2 _331_ (.A_N(_009_),
    .B(_010_),
    .X(_011_));
 sky130_fd_sc_hd__xnor2_4 _332_ (.A(_001_),
    .B(_011_),
    .Y(_012_));
 sky130_fd_sc_hd__nand2_4 _333_ (.A(_012_),
    .B(_224_),
    .Y(_013_));
 sky130_fd_sc_hd__or2_1 _334_ (.A(_224_),
    .B(_012_),
    .X(_014_));
 sky130_fd_sc_hd__a21oi_1 _335_ (.A1(net66),
    .A2(_241_),
    .B1(_200_),
    .Y(_015_));
 sky130_fd_sc_hd__o22a_1 _336_ (.A1(net66),
    .A2(_241_),
    .B1(_198_),
    .B2(_015_),
    .X(_016_));
 sky130_fd_sc_hd__a311o_1 _337_ (.A1(net66),
    .A2(_241_),
    .A3(_190_),
    .B1(_195_),
    .C1(_016_),
    .X(_017_));
 sky130_fd_sc_hd__a31o_1 _338_ (.A1(_189_),
    .A2(_013_),
    .A3(_014_),
    .B1(_017_),
    .X(_018_));
 sky130_fd_sc_hd__o2bb2a_1 _339_ (.A1_N(net66),
    .A2_N(_195_),
    .B1(_000_),
    .B2(_018_),
    .X(net23));
 sky130_fd_sc_hd__buf_12 _340_ (.A(net5),
    .X(_019_));
 sky130_fd_sc_hd__a31o_4 _341_ (.A1(_176_),
    .A2(_241_),
    .A3(_010_),
    .B1(net58),
    .X(_020_));
 sky130_fd_sc_hd__buf_8 _342_ (.A(net13),
    .X(_021_));
 sky130_fd_sc_hd__a22o_2 _343_ (.A1(net43),
    .A2(net61),
    .B1(_021_),
    .B2(net1),
    .X(_022_));
 sky130_fd_sc_hd__and4_2 _344_ (.A(net1),
    .B(net2),
    .C(net12),
    .D(net13),
    .X(_023_));
 sky130_fd_sc_hd__clkinv_4 _345_ (.A(_023_),
    .Y(_024_));
 sky130_fd_sc_hd__and2_4 _346_ (.A(_022_),
    .B(_024_),
    .X(_025_));
 sky130_fd_sc_hd__and4_4 _347_ (.A(net9),
    .B(net10),
    .C(net4),
    .D(net5),
    .X(_026_));
 sky130_fd_sc_hd__a22oi_4 _348_ (.A1(net4),
    .A2(net10),
    .B1(net5),
    .B2(net9),
    .Y(_027_));
 sky130_fd_sc_hd__or3_4 _349_ (.A(_233_),
    .B(_027_),
    .C(_026_),
    .X(_028_));
 sky130_fd_sc_hd__o21ai_4 _350_ (.A1(_026_),
    .A2(_027_),
    .B1(_233_),
    .Y(_029_));
 sky130_fd_sc_hd__o21bai_4 _351_ (.A1(_002_),
    .A2(net64),
    .B1_N(_003_),
    .Y(_030_));
 sky130_fd_sc_hd__and3_4 _352_ (.A(_028_),
    .B(_029_),
    .C(_030_),
    .X(_031_));
 sky130_fd_sc_hd__a21o_4 _353_ (.A1(_028_),
    .A2(_029_),
    .B1(_030_),
    .X(_032_));
 sky130_fd_sc_hd__or2b_4 _354_ (.A(_031_),
    .B_N(_032_),
    .X(_033_));
 sky130_fd_sc_hd__xnor2_4 _355_ (.A(_025_),
    .B(_033_),
    .Y(_034_));
 sky130_fd_sc_hd__nand2_8 _356_ (.A(_020_),
    .B(_034_),
    .Y(_035_));
 sky130_fd_sc_hd__or2_4 _357_ (.A(_020_),
    .B(_034_),
    .X(_036_));
 sky130_fd_sc_hd__a21bo_1 _358_ (.A1(_035_),
    .A2(_036_),
    .B1_N(_013_),
    .X(_037_));
 sky130_fd_sc_hd__nand3b_4 _359_ (.A_N(_013_),
    .B(_035_),
    .C(_036_),
    .Y(_038_));
 sky130_fd_sc_hd__and3_2 _360_ (.A(_189_),
    .B(_037_),
    .C(_038_),
    .X(_039_));
 sky130_fd_sc_hd__o31a_4 _361_ (.A1(_218_),
    .A2(_241_),
    .A3(_227_),
    .B1(net49),
    .X(_040_));
 sky130_fd_sc_hd__xnor2_4 _362_ (.A(_021_),
    .B(_040_),
    .Y(_041_));
 sky130_fd_sc_hd__and2_2 _363_ (.A(_019_),
    .B(_041_),
    .X(_042_));
 sky130_fd_sc_hd__nor2_2 _364_ (.A(_019_),
    .B(_041_),
    .Y(_043_));
 sky130_fd_sc_hd__nor2_2 _365_ (.A(_042_),
    .B(_043_),
    .Y(_044_));
 sky130_fd_sc_hd__a21bo_2 _366_ (.A1(_240_),
    .A2(_245_),
    .B1_N(_244_),
    .X(_045_));
 sky130_fd_sc_hd__nand2_2 _367_ (.A(_044_),
    .B(_045_),
    .Y(_046_));
 sky130_fd_sc_hd__or2_2 _368_ (.A(_044_),
    .B(_045_),
    .X(_047_));
 sky130_fd_sc_hd__a21oi_4 _369_ (.A1(_019_),
    .A2(_021_),
    .B1(_200_),
    .Y(_048_));
 sky130_fd_sc_hd__o22a_2 _370_ (.A1(_019_),
    .A2(_021_),
    .B1(_198_),
    .B2(_048_),
    .X(_049_));
 sky130_fd_sc_hd__a311o_1 _371_ (.A1(_019_),
    .A2(_021_),
    .A3(_190_),
    .B1(_194_),
    .C1(_049_),
    .X(_050_));
 sky130_fd_sc_hd__a31o_1 _372_ (.A1(_203_),
    .A2(_046_),
    .A3(_047_),
    .B1(_050_),
    .X(_051_));
 sky130_fd_sc_hd__o2bb2a_2 _373_ (.A1_N(_019_),
    .A2_N(_195_),
    .B1(_039_),
    .B2(_051_),
    .X(net24));
 sky130_fd_sc_hd__buf_12 _374_ (.A(net6),
    .X(_052_));
 sky130_fd_sc_hd__a21o_4 _375_ (.A1(_044_),
    .A2(_045_),
    .B1(_042_),
    .X(_053_));
 sky130_fd_sc_hd__a21o_4 _376_ (.A1(_021_),
    .A2(net32),
    .B1(_040_),
    .X(_054_));
 sky130_fd_sc_hd__xnor2_4 _377_ (.A(net14),
    .B(_054_),
    .Y(_055_));
 sky130_fd_sc_hd__and2_4 _378_ (.A(_052_),
    .B(_055_),
    .X(_056_));
 sky130_fd_sc_hd__nor2_1 _379_ (.A(_052_),
    .B(_055_),
    .Y(_057_));
 sky130_fd_sc_hd__nor2_4 _380_ (.A(_056_),
    .B(_057_),
    .Y(_058_));
 sky130_fd_sc_hd__xor2_1 _381_ (.A(_053_),
    .B(_058_),
    .X(_059_));
 sky130_fd_sc_hd__nand4_4 _382_ (.A(net47),
    .B(_182_),
    .C(_019_),
    .D(net6),
    .Y(_060_));
 sky130_fd_sc_hd__a22o_4 _383_ (.A1(net5),
    .A2(_196_),
    .B1(net6),
    .B2(net9),
    .X(_061_));
 sky130_fd_sc_hd__and2_4 _384_ (.A(net11),
    .B(net4),
    .X(_062_));
 sky130_fd_sc_hd__a21o_4 _385_ (.A1(_061_),
    .A2(_060_),
    .B1(_062_),
    .X(_063_));
 sky130_fd_sc_hd__nand3_4 _386_ (.A(_062_),
    .B(net38),
    .C(net37),
    .Y(_064_));
 sky130_fd_sc_hd__o21bai_4 _387_ (.A1(_233_),
    .A2(_027_),
    .B1_N(_026_),
    .Y(_065_));
 sky130_fd_sc_hd__nand3_4 _388_ (.A(_063_),
    .B(_064_),
    .C(_065_),
    .Y(_066_));
 sky130_fd_sc_hd__a21o_4 _389_ (.A1(_064_),
    .A2(_063_),
    .B1(_065_),
    .X(_067_));
 sky130_fd_sc_hd__nand2_4 _390_ (.A(net1),
    .B(net14),
    .Y(_068_));
 sky130_fd_sc_hd__and4_4 _391_ (.A(net13),
    .B(net3),
    .C(net12),
    .D(net2),
    .X(_069_));
 sky130_fd_sc_hd__a22o_2 _392_ (.A1(net3),
    .A2(net12),
    .B1(net13),
    .B2(net2),
    .X(_070_));
 sky130_fd_sc_hd__and2b_2 _393_ (.A_N(_069_),
    .B(_070_),
    .X(_071_));
 sky130_fd_sc_hd__xnor2_4 _394_ (.A(_071_),
    .B(_068_),
    .Y(_072_));
 sky130_fd_sc_hd__a21o_4 _395_ (.A1(_067_),
    .A2(_066_),
    .B1(net31),
    .X(_073_));
 sky130_fd_sc_hd__nand3_4 _396_ (.A(_072_),
    .B(_066_),
    .C(_067_),
    .Y(_074_));
 sky130_fd_sc_hd__a21o_4 _397_ (.A1(_025_),
    .A2(_032_),
    .B1(_031_),
    .X(_075_));
 sky130_fd_sc_hd__and3_4 _398_ (.A(_073_),
    .B(_074_),
    .C(_075_),
    .X(_076_));
 sky130_fd_sc_hd__a21oi_4 _399_ (.A1(_074_),
    .A2(_073_),
    .B1(_075_),
    .Y(_077_));
 sky130_fd_sc_hd__o21ai_4 _400_ (.A1(net52),
    .A2(net53),
    .B1(_024_),
    .Y(_078_));
 sky130_fd_sc_hd__or3_4 _401_ (.A(_024_),
    .B(_077_),
    .C(_076_),
    .X(_079_));
 sky130_fd_sc_hd__nand2_4 _402_ (.A(_078_),
    .B(net34),
    .Y(_080_));
 sky130_fd_sc_hd__a21o_4 _403_ (.A1(_035_),
    .A2(_038_),
    .B1(_080_),
    .X(_081_));
 sky130_fd_sc_hd__nand3_2 _404_ (.A(_035_),
    .B(_038_),
    .C(_080_),
    .Y(_082_));
 sky130_fd_sc_hd__a21oi_2 _405_ (.A1(_052_),
    .A2(net14),
    .B1(_200_),
    .Y(_083_));
 sky130_fd_sc_hd__o22a_1 _406_ (.A1(_052_),
    .A2(net14),
    .B1(_198_),
    .B2(_083_),
    .X(_084_));
 sky130_fd_sc_hd__a311o_2 _407_ (.A1(_052_),
    .A2(net14),
    .A3(_190_),
    .B1(_194_),
    .C1(_084_),
    .X(_085_));
 sky130_fd_sc_hd__a31o_1 _408_ (.A1(_189_),
    .A2(_081_),
    .A3(_082_),
    .B1(_085_),
    .X(_086_));
 sky130_fd_sc_hd__a21oi_1 _409_ (.A1(_203_),
    .A2(_059_),
    .B1(_086_),
    .Y(_087_));
 sky130_fd_sc_hd__a21oi_2 _410_ (.A1(_052_),
    .A2(_195_),
    .B1(_087_),
    .Y(net25));
 sky130_fd_sc_hd__nand3_4 _411_ (.A(_073_),
    .B(_074_),
    .C(_075_),
    .Y(_088_));
 sky130_fd_sc_hd__a31o_2 _412_ (.A1(net1),
    .A2(net14),
    .A3(_070_),
    .B1(_069_),
    .X(_089_));
 sky130_fd_sc_hd__and3_4 _413_ (.A(net1),
    .B(net15),
    .C(_089_),
    .X(_090_));
 sky130_fd_sc_hd__a21oi_4 _414_ (.A1(_176_),
    .A2(net15),
    .B1(_089_),
    .Y(_091_));
 sky130_fd_sc_hd__nor2_4 _415_ (.A(_090_),
    .B(_091_),
    .Y(_092_));
 sky130_fd_sc_hd__nand4_4 _416_ (.A(_182_),
    .B(net47),
    .C(_052_),
    .D(net7),
    .Y(_093_));
 sky130_fd_sc_hd__a22o_4 _417_ (.A1(_196_),
    .A2(_052_),
    .B1(net7),
    .B2(net63),
    .X(_094_));
 sky130_fd_sc_hd__and2_4 _418_ (.A(net11),
    .B(_019_),
    .X(_095_));
 sky130_fd_sc_hd__a21o_2 _419_ (.A1(_093_),
    .A2(_094_),
    .B1(_095_),
    .X(_096_));
 sky130_fd_sc_hd__nand3_2 _420_ (.A(_095_),
    .B(_093_),
    .C(_094_),
    .Y(_097_));
 sky130_fd_sc_hd__a21bo_4 _421_ (.A1(_062_),
    .A2(_061_),
    .B1_N(net38),
    .X(_098_));
 sky130_fd_sc_hd__nand3_4 _422_ (.A(_096_),
    .B(_097_),
    .C(_098_),
    .Y(_099_));
 sky130_fd_sc_hd__a21o_4 _423_ (.A1(_096_),
    .A2(_097_),
    .B1(_098_),
    .X(_100_));
 sky130_fd_sc_hd__nand2_4 _424_ (.A(_193_),
    .B(net14),
    .Y(_101_));
 sky130_fd_sc_hd__and3_4 _425_ (.A(_238_),
    .B(net60),
    .C(net13),
    .X(_102_));
 sky130_fd_sc_hd__a22o_2 _426_ (.A1(net4),
    .A2(net12),
    .B1(_021_),
    .B2(net57),
    .X(_103_));
 sky130_fd_sc_hd__a21bo_4 _427_ (.A1(_217_),
    .A2(_102_),
    .B1_N(_103_),
    .X(_104_));
 sky130_fd_sc_hd__xor2_4 _428_ (.A(_101_),
    .B(_104_),
    .X(_105_));
 sky130_fd_sc_hd__a21o_4 _429_ (.A1(_099_),
    .A2(_100_),
    .B1(_105_),
    .X(_106_));
 sky130_fd_sc_hd__nand3_4 _430_ (.A(_105_),
    .B(_099_),
    .C(_100_),
    .Y(_107_));
 sky130_fd_sc_hd__a21bo_4 _431_ (.A1(net31),
    .A2(_067_),
    .B1_N(_066_),
    .X(_108_));
 sky130_fd_sc_hd__nand3_4 _432_ (.A(_106_),
    .B(_107_),
    .C(_108_),
    .Y(_109_));
 sky130_fd_sc_hd__a21o_4 _433_ (.A1(_106_),
    .A2(_107_),
    .B1(_108_),
    .X(_110_));
 sky130_fd_sc_hd__and3_4 _434_ (.A(_092_),
    .B(_109_),
    .C(_110_),
    .X(_111_));
 sky130_fd_sc_hd__a21oi_4 _435_ (.A1(_109_),
    .A2(_110_),
    .B1(_092_),
    .Y(_112_));
 sky130_fd_sc_hd__a211oi_4 _436_ (.A1(net33),
    .A2(_088_),
    .B1(_111_),
    .C1(_112_),
    .Y(_113_));
 sky130_fd_sc_hd__o211a_2 _437_ (.A1(_111_),
    .A2(_112_),
    .B1(_088_),
    .C1(_079_),
    .X(_114_));
 sky130_fd_sc_hd__a2111oi_4 _438_ (.A1(_035_),
    .A2(_038_),
    .B1(_080_),
    .C1(net42),
    .D1(_114_),
    .Y(_115_));
 sky130_fd_sc_hd__or2_4 _439_ (.A(_113_),
    .B(_114_),
    .X(_116_));
 sky130_fd_sc_hd__a21bo_2 _440_ (.A1(_081_),
    .A2(_116_),
    .B1_N(_189_),
    .X(_117_));
 sky130_fd_sc_hd__or2_4 _441_ (.A(net28),
    .B(_117_),
    .X(_118_));
 sky130_fd_sc_hd__a21o_4 _442_ (.A1(_053_),
    .A2(_058_),
    .B1(_056_),
    .X(_119_));
 sky130_fd_sc_hd__or2_4 _443_ (.A(net14),
    .B(_054_),
    .X(_120_));
 sky130_fd_sc_hd__nand2_4 _444_ (.A(net32),
    .B(_120_),
    .Y(_121_));
 sky130_fd_sc_hd__xor2_4 _445_ (.A(net15),
    .B(_121_),
    .X(_122_));
 sky130_fd_sc_hd__xor2_4 _446_ (.A(net7),
    .B(_122_),
    .X(_123_));
 sky130_fd_sc_hd__nand2_1 _447_ (.A(_119_),
    .B(net48),
    .Y(_124_));
 sky130_fd_sc_hd__o21a_1 _448_ (.A1(_119_),
    .A2(net48),
    .B1(_203_),
    .X(_125_));
 sky130_fd_sc_hd__a21oi_1 _449_ (.A1(net7),
    .A2(net15),
    .B1(_200_),
    .Y(_126_));
 sky130_fd_sc_hd__o22a_1 _450_ (.A1(net7),
    .A2(net15),
    .B1(_198_),
    .B2(_126_),
    .X(_127_));
 sky130_fd_sc_hd__a311o_2 _451_ (.A1(net7),
    .A2(net15),
    .A3(_190_),
    .B1(_195_),
    .C1(_127_),
    .X(_128_));
 sky130_fd_sc_hd__a21oi_4 _452_ (.A1(_124_),
    .A2(_125_),
    .B1(_128_),
    .Y(_129_));
 sky130_fd_sc_hd__a22oi_4 _453_ (.A1(net7),
    .A2(_195_),
    .B1(_129_),
    .B2(_118_),
    .Y(net26));
 sky130_fd_sc_hd__and2_2 _454_ (.A(net7),
    .B(_122_),
    .X(_130_));
 sky130_fd_sc_hd__a21oi_1 _455_ (.A1(_119_),
    .A2(_123_),
    .B1(_130_),
    .Y(_131_));
 sky130_fd_sc_hd__o21ai_4 _456_ (.A1(net15),
    .A2(_120_),
    .B1(net32),
    .Y(_132_));
 sky130_fd_sc_hd__nand2_2 _457_ (.A(net8),
    .B(net16),
    .Y(_133_));
 sky130_fd_sc_hd__or2_2 _458_ (.A(net8),
    .B(net16),
    .X(_134_));
 sky130_fd_sc_hd__nand2_1 _459_ (.A(_133_),
    .B(_134_),
    .Y(_135_));
 sky130_fd_sc_hd__and2b_2 _460_ (.A_N(_132_),
    .B(_135_),
    .X(_136_));
 sky130_fd_sc_hd__and2b_2 _461_ (.A_N(_135_),
    .B(_132_),
    .X(_137_));
 sky130_fd_sc_hd__nor2_1 _462_ (.A(_136_),
    .B(_137_),
    .Y(_138_));
 sky130_fd_sc_hd__a211o_2 _463_ (.A1(_119_),
    .A2(_123_),
    .B1(_138_),
    .C1(_130_),
    .X(_139_));
 sky130_fd_sc_hd__o311a_2 _464_ (.A1(_131_),
    .A2(_136_),
    .A3(_137_),
    .B1(_139_),
    .C1(_203_),
    .X(_140_));
 sky130_fd_sc_hd__a211o_4 _465_ (.A1(_079_),
    .A2(_088_),
    .B1(_111_),
    .C1(_112_),
    .X(_141_));
 sky130_fd_sc_hd__a22o_4 _466_ (.A1(_238_),
    .A2(_021_),
    .B1(_052_),
    .B2(net11),
    .X(_142_));
 sky130_fd_sc_hd__nand4_4 _467_ (.A(_218_),
    .B(_238_),
    .C(_021_),
    .D(_052_),
    .Y(_143_));
 sky130_fd_sc_hd__a22oi_4 _468_ (.A1(net47),
    .A2(net7),
    .B1(net8),
    .B2(net59),
    .Y(_144_));
 sky130_fd_sc_hd__and4_2 _469_ (.A(_182_),
    .B(_196_),
    .C(net7),
    .D(net8),
    .X(_145_));
 sky130_fd_sc_hd__a211o_4 _470_ (.A1(_143_),
    .A2(_142_),
    .B1(_144_),
    .C1(_145_),
    .X(_146_));
 sky130_fd_sc_hd__o211ai_4 _471_ (.A1(_144_),
    .A2(_145_),
    .B1(_142_),
    .C1(_143_),
    .Y(_147_));
 sky130_fd_sc_hd__a22o_4 _472_ (.A1(_241_),
    .A2(_019_),
    .B1(_146_),
    .B2(_147_),
    .X(_148_));
 sky130_fd_sc_hd__nand4_4 _473_ (.A(_147_),
    .B(_019_),
    .C(_146_),
    .D(_241_),
    .Y(_149_));
 sky130_fd_sc_hd__a21bo_2 _474_ (.A1(_095_),
    .A2(_094_),
    .B1_N(_093_),
    .X(_150_));
 sky130_fd_sc_hd__nand2_2 _475_ (.A(_217_),
    .B(net14),
    .Y(_151_));
 sky130_fd_sc_hd__xor2_4 _476_ (.A(_151_),
    .B(_150_),
    .X(_152_));
 sky130_fd_sc_hd__a21o_4 _477_ (.A1(_148_),
    .A2(_149_),
    .B1(_152_),
    .X(_153_));
 sky130_fd_sc_hd__nand3_4 _478_ (.A(_152_),
    .B(_148_),
    .C(_149_),
    .Y(_154_));
 sky130_fd_sc_hd__and4_4 _479_ (.A(net55),
    .B(net4),
    .C(net61),
    .D(_021_),
    .X(_155_));
 sky130_fd_sc_hd__a31o_2 _480_ (.A1(net44),
    .A2(net14),
    .A3(_103_),
    .B1(_155_),
    .X(_156_));
 sky130_fd_sc_hd__nand2_4 _481_ (.A(net1),
    .B(net16),
    .Y(_157_));
 sky130_fd_sc_hd__nand2_2 _482_ (.A(net45),
    .B(net15),
    .Y(_158_));
 sky130_fd_sc_hd__xor2_4 _483_ (.A(_157_),
    .B(_158_),
    .X(_159_));
 sky130_fd_sc_hd__xnor2_2 _484_ (.A(_156_),
    .B(_159_),
    .Y(_160_));
 sky130_fd_sc_hd__xnor2_4 _485_ (.A(_090_),
    .B(_160_),
    .Y(_161_));
 sky130_fd_sc_hd__a21o_4 _486_ (.A1(_153_),
    .A2(_154_),
    .B1(_161_),
    .X(_162_));
 sky130_fd_sc_hd__nand3_4 _487_ (.A(_153_),
    .B(_154_),
    .C(_161_),
    .Y(_163_));
 sky130_fd_sc_hd__nand2_4 _488_ (.A(_099_),
    .B(_107_),
    .Y(_164_));
 sky130_fd_sc_hd__a21o_2 _489_ (.A1(_162_),
    .A2(_163_),
    .B1(_164_),
    .X(_165_));
 sky130_fd_sc_hd__nand3_4 _490_ (.A(_164_),
    .B(_162_),
    .C(_163_),
    .Y(_166_));
 sky130_fd_sc_hd__a21boi_4 _491_ (.A1(_092_),
    .A2(_110_),
    .B1_N(_109_),
    .Y(_167_));
 sky130_fd_sc_hd__a21oi_4 _492_ (.A1(_165_),
    .A2(_166_),
    .B1(_167_),
    .Y(_168_));
 sky130_fd_sc_hd__and3_4 _493_ (.A(_165_),
    .B(_167_),
    .C(_166_),
    .X(_169_));
 sky130_fd_sc_hd__or3_4 _494_ (.A(_169_),
    .B(_168_),
    .C(_141_),
    .X(_170_));
 sky130_fd_sc_hd__o21ai_4 _495_ (.A1(_168_),
    .A2(_169_),
    .B1(net41),
    .Y(_171_));
 sky130_fd_sc_hd__and3_1 _496_ (.A(_170_),
    .B(net29),
    .C(_171_),
    .X(_172_));
 sky130_fd_sc_hd__a21oi_4 _497_ (.A1(net35),
    .A2(_171_),
    .B1(net36),
    .Y(_173_));
 sky130_fd_sc_hd__o21a_1 _498_ (.A1(_173_),
    .A2(_172_),
    .B1(_189_),
    .X(_174_));
 sky130_fd_sc_hd__o21ai_4 _499_ (.A1(net8),
    .A2(net16),
    .B1(_198_),
    .Y(_175_));
 sky130_fd_sc_hd__o221a_1 _500_ (.A1(_187_),
    .A2(_133_),
    .B1(_135_),
    .B2(_200_),
    .C1(_181_),
    .X(_177_));
 sky130_fd_sc_hd__nand2_1 _501_ (.A(_175_),
    .B(_177_),
    .Y(_178_));
 sky130_fd_sc_hd__inv_2 _502_ (.A(net8),
    .Y(_179_));
 sky130_fd_sc_hd__o32a_4 _503_ (.A1(_140_),
    .A2(_178_),
    .A3(_174_),
    .B1(_181_),
    .B2(_179_),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_16 clone15 (.A(net10),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_16 clone16 (.A(net11),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_16 clone17 (.A(net4),
    .X(net66));
 sky130_fd_sc_hd__buf_12 clone31 (.A(net9),
    .X(net63));
 sky130_fd_sc_hd__buf_8 input1 (.A(A[0]),
    .X(net1));
 sky130_fd_sc_hd__buf_8 input10 (.A(B[1]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_8 input11 (.A(B[2]),
    .X(net11));
 sky130_fd_sc_hd__buf_12 input12 (.A(B[3]),
    .X(net12));
 sky130_fd_sc_hd__buf_8 input13 (.A(B[4]),
    .X(net13));
 sky130_fd_sc_hd__buf_8 input14 (.A(B[5]),
    .X(net14));
 sky130_fd_sc_hd__buf_8 input15 (.A(B[6]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_8 input16 (.A(B[7]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_8 input17 (.A(opcode[0]),
    .X(net17));
 sky130_fd_sc_hd__buf_6 input18 (.A(opcode[1]),
    .X(net18));
 sky130_fd_sc_hd__buf_6 input19 (.A(opcode[2]),
    .X(net19));
 sky130_fd_sc_hd__buf_12 input2 (.A(A[1]),
    .X(net2));
 sky130_fd_sc_hd__buf_12 input3 (.A(A[2]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_8 input4 (.A(A[3]),
    .X(net4));
 sky130_fd_sc_hd__buf_4 input5 (.A(A[4]),
    .X(net5));
 sky130_fd_sc_hd__buf_4 input6 (.A(A[5]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_16 input7 (.A(A[6]),
    .X(net7));
 sky130_fd_sc_hd__buf_8 input8 (.A(A[7]),
    .X(net8));
 sky130_fd_sc_hd__buf_8 input9 (.A(B[0]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_2 max_cap30 (.A(_242_),
    .X(net30));
 sky130_fd_sc_hd__buf_6 max_cap31 (.A(_072_),
    .X(net31));
 sky130_fd_sc_hd__buf_6 max_cap32 (.A(_205_),
    .X(net32));
 sky130_fd_sc_hd__buf_2 output20 (.A(net20),
    .X(out[0]));
 sky130_fd_sc_hd__buf_2 output21 (.A(net21),
    .X(out[1]));
 sky130_fd_sc_hd__buf_2 output22 (.A(net22),
    .X(out[2]));
 sky130_fd_sc_hd__buf_2 output23 (.A(net23),
    .X(out[3]));
 sky130_fd_sc_hd__buf_2 output24 (.A(net24),
    .X(out[4]));
 sky130_fd_sc_hd__buf_2 output25 (.A(net25),
    .X(out[5]));
 sky130_fd_sc_hd__buf_6 output26 (.A(net26),
    .X(out[6]));
 sky130_fd_sc_hd__buf_8 output27 (.A(net27),
    .X(out[7]));
 sky130_fd_sc_hd__clkbuf_2 rebuffer1 (.A(_079_),
    .X(net33));
 sky130_fd_sc_hd__buf_6 rebuffer10 (.A(_113_),
    .X(net42));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer11 (.A(net2),
    .X(net43));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer12 (.A(net2),
    .X(net44));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer13 (.A(net44),
    .X(net45));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer14 (.A(net2),
    .X(net46));
 sky130_fd_sc_hd__buf_2 rebuffer15 (.A(_004_),
    .X(net64));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer16 (.A(_123_),
    .X(net48));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer17 (.A(_205_),
    .X(net49));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer18 (.A(_205_),
    .X(net50));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer19 (.A(net50),
    .X(net51));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer2 (.A(_079_),
    .X(net34));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer20 (.A(_076_),
    .X(net52));
 sky130_fd_sc_hd__dlymetal6s4s_1 rebuffer21 (.A(_077_),
    .X(net53));
 sky130_fd_sc_hd__buf_12 rebuffer22 (.A(net3),
    .X(net54));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer23 (.A(net54),
    .X(net55));
 sky130_fd_sc_hd__buf_2 rebuffer24 (.A(net54),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_2 rebuffer25 (.A(net3),
    .X(net57));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer26 (.A(_009_),
    .X(net58));
 sky130_fd_sc_hd__buf_2 rebuffer27 (.A(_182_),
    .X(net59));
 sky130_fd_sc_hd__dlymetal6s4s_1 rebuffer28 (.A(net12),
    .X(net60));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer29 (.A(net12),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_2 rebuffer3 (.A(_170_),
    .X(net35));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer30 (.A(net12),
    .X(net62));
 sky130_fd_sc_hd__buf_6 rebuffer4 (.A(_115_),
    .X(net36));
 sky130_fd_sc_hd__buf_6 rebuffer5 (.A(_061_),
    .X(net37));
 sky130_fd_sc_hd__buf_6 rebuffer6 (.A(_060_),
    .X(net38));
 sky130_fd_sc_hd__buf_6 rebuffer7 (.A(_004_),
    .X(net39));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer8 (.A(net39),
    .X(net40));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer9 (.A(_141_),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_2 wire28 (.A(net29),
    .X(net28));
 sky130_fd_sc_hd__buf_2 wire29 (.A(_115_),
    .X(net29));
endmodule

